// IWLS benchmark module "pm1" printed on Wed May 29 17:28:07 2002
module pm1(a, b, c, d, e, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, \xx , y, z, a0, b0, c0, d0);
input
  a,
  b,
  c,
  d,
  e,
  g,
  h,
  i,
  j,
  k,
  l,
  m,
  n,
  o,
  p,
  q;
output
  r,
  s,
  t,
  u,
  v,
  w,
  \xx ,
  y,
  z,
  a0,
  b0,
  c0,
  d0;
wire
  k1,
  l1,
  m1,
  n1,
  o1,
  r1,
  s0,
  s1,
  \[0] ,
  a1,
  t0,
  t1,
  \[1] ,
  u1,
  \[2] ,
  v1,
  \[3] ,
  d1,
  \[4] ,
  e1,
  \[5] ,
  y0,
  \[6] ,
  z0,
  \[7] ,
  \[8] ,
  \[10] ,
  i1,
  \[9] ,
  \[11] ,
  \[12] ;
assign
  k1 = ~b & (~m & ~n),
  l1 = ~m & n,
  m1 = ~o1 | (~g | ~h),
  n1 = ~m1 & (m & n),
  o1 = i & (j & k),
  r = \[0] ,
  s = \[1] ,
  r1 = (n & ~s1) | ((n & ~g) | (n & ~h)),
  t = \[2] ,
  u = \[3] ,
  v = \[4] ,
  w = \[5] ,
  \xx  = \[6] ,
  y = \[7] ,
  z = \[8] ,
  s0 = (m & ~t0) | ((m & ~c) | (m & ~d)),
  s1 = i & j,
  \[0]  = ~k1,
  a0 = \[9] ,
  a1 = (a & (k & ~e)) | ((a & (k & ~d)) | (a & (k & ~c))),
  t0 = e & (k & n),
  t1 = d & e,
  \[1]  = ~l1,
  b0 = \[10] ,
  u1 = m | ~n,
  \[2]  = ~n1,
  c0 = \[11] ,
  v1 = ~b | ~k,
  \[3]  = ~r1 | (~k | ~m),
  d0 = \[12] ,
  d1 = (e & (d & c)) | (~n | ~k),
  \[4]  = ~p,
  e1 = (n & ~b) | (~a | l),
  \[5]  = ~o,
  y0 = (n & ~m) | (~a | l),
  \[6]  = (~v1 & ~u1) | ((~v1 & ~t1) | (~v1 & ~c)),
  z0 = ~a1 | l,
  \[7]  = ~q,
  \[8]  = ~s0 | (l | ~a),
  \[10]  = ~z0 & (m & n),
  i1 = ~a | (k | l),
  \[9]  = (~y0 & ~m) | (~y0 & n),
  \[11]  = (~e1 & (m & ~d1)) | (~e1 & (m & ~b)),
  \[12]  = ~i1 & (m & n);
endmodule

