module s1488 (
  CK,
  CLR,
  v0,
  v1,
  v2,
  v3,
  v4,
  v5,
  v6,
  v13_D_9,
  v13_D_24,
  v13_D_15,
  v13_D_21,
  v13_D_10,
  v13_D_13,
  v13_D_17,
  v13_D_22,
  v13_D_20,
  v13_D_16,
  v13_D_19,
  v13_D_6,
  v13_D_8,
  v13_D_18,
  v13_D_14,
  v13_D_12,
  v13_D_23,
  v13_D_11,
  v13_D_7
);
  input CK;
  wire CK;
  input CLR;
  wire CLR;
  input v0;
  wire v0;
  input v1;
  wire v1;
  input v2;
  wire v2;
  input v3;
  wire v3;
  input v4;
  wire v4;
  input v5;
  wire v5;
  input v6;
  wire v6;
  output v13_D_9;
  wire v13_D_9;
  output v13_D_24;
  wire v13_D_24;
  output v13_D_15;
  wire v13_D_15;
  output v13_D_21;
  wire v13_D_21;
  output v13_D_10;
  wire v13_D_10;
  output v13_D_13;
  wire v13_D_13;
  output v13_D_17;
  wire v13_D_17;
  output v13_D_22;
  wire v13_D_22;
  output v13_D_20;
  wire v13_D_20;
  output v13_D_16;
  wire v13_D_16;
  output v13_D_19;
  wire v13_D_19;
  output v13_D_6;
  wire v13_D_6;
  output v13_D_8;
  wire v13_D_8;
  output v13_D_18;
  wire v13_D_18;
  output v13_D_14;
  wire v13_D_14;
  output v13_D_12;
  wire v13_D_12;
  output v13_D_23;
  wire v13_D_23;
  output v13_D_11;
  wire v13_D_11;
  output v13_D_7;
  wire v13_D_7;
  wire __0__;
  wire __1__;
  wire __2__;
  wire __3__;
  wire __4__;
  wire __5__;
  wire __6__;
  wire __7__;
  wire __8__;
  wire __9__;
  wire __10__;
  wire __11__;
  wire __12__;
  wire __13__;
  wire __14__;
  wire __15__;
  wire __16__;
  wire __17__;
  wire __18__;
  wire __19__;
  wire __20__;
  wire __21__;
  wire __22__;
  wire __23__;
  wire __24__;
  wire __25__;
  wire __26__;
  wire __27__;
  wire __28__;
  wire __29__;
  wire __30__;
  wire __31__;
  wire __33__;
  wire __34__;
  wire __35__;
  wire __36__;
  wire __37__;
  wire __38__;
  wire __39__;
  wire __40__;
  wire __41__;
  wire __42__;
  wire __43__;
  wire __44__;
  wire __45__;
  wire __46__;
  wire __47__;
  wire __48__;
  wire __49__;
  wire __50__;
  wire __51__;
  wire __52__;
  wire __53__;
  wire __54__;
  wire __55__;
  wire __56__;
  wire __57__;
  wire __58__;
  wire __59__;
  wire __60__;
  wire __61__;
  wire __62__;
  wire __63__;
  wire __64__;
  wire __65__;
  wire __66__;
  wire __67__;
  wire __68__;
  wire __69__;
  wire __70__;
  wire __71__;
  wire __72__;
  wire __73__;
  wire __74__;
  wire __75__;
  wire __76__;
  wire __77__;
  wire __78__;
  wire __79__;
  wire __80__;
  wire __81__;
  wire __82__;
  wire __83__;
  wire __84__;
  wire __85__;
  wire __86__;
  wire __87__;
  wire __88__;
  wire __89__;
  wire __90__;
  wire __91__;
  wire __92__;
  wire __93__;
  wire __94__;
  wire __95__;
  wire __96__;
  wire __97__;
  wire __98__;
  wire __99__;
  wire __100__;
  wire __101__;
  wire __102__;
  wire __103__;
  wire __104__;
  wire __105__;
  wire __106__;
  wire __107__;
  wire __108__;
  wire __109__;
  wire __110__;
  wire __111__;
  wire __112__;
  wire __113__;
  wire __114__;
  wire __115__;
  wire __116__;
  wire __117__;
  wire __118__;
  wire __119__;
  wire __121__;
  wire __122__;
  wire __123__;
  wire __124__;
  wire __125__;
  wire __126__;
  wire __127__;
  wire __128__;
  wire __129__;
  wire __130__;
  wire __131__;
  wire __132__;
  wire __133__;
  wire __134__;
  wire __135__;
  wire __136__;
  wire __137__;
  wire __138__;
  wire __139__;
  wire __140__;
  wire __141__;
  wire __142__;
  wire __143__;
  wire __144__;
  wire __145__;
  wire __146__;
  wire __147__;
  wire __148__;
  wire __149__;
  wire __150__;
  wire __151__;
  wire __152__;
  wire __153__;
  wire __154__;
  wire __155__;
  wire __156__;
  wire __157__;
  wire __158__;
  wire __159__;
  wire __160__;
  wire __161__;
  wire __162__;
  wire __163__;
  wire __164__;
  FDRE #(
    .INIT(1'bx)
  ) __165__ (
    .D(__115__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__0__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __166__ (
    .D(__106__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __167__ (
    .D(__70__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__2__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __168__ (
    .D(__85__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__3__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __169__ (
    .D(__46__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__4__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __170__ (
    .D(__60__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__5__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __171__ (
    .I1(__4__),
    .I0(__1__),
    .O(__6__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __172__ (
    .I1(__2__),
    .I0(__3__),
    .O(__7__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __173__ (
    .I1(v6),
    .I0(v3),
    .O(__8__)
  );
  LUT6 #(
    .INIT(64'h33330f0fff005555)
  ) __174__ (
    .I5(__2__),
    .I4(__4__),
    .I3(__8__),
    .I2(v0),
    .I1(v2),
    .I0(__1__),
    .O(__9__)
  );
  LUT6 #(
    .INIT(64'h000000007707ff07)
  ) __175__ (
    .I5(__3__),
    .I4(__2__),
    .I3(__4__),
    .I2(__5__),
    .I1(v5),
    .I0(v4),
    .O(__10__)
  );
  LUT4 #(
    .INIT(16'h1f00)
  ) __176__ (
    .I3(__4__),
    .I2(__5__),
    .I1(__2__),
    .I0(__1__),
    .O(__11__)
  );
  LUT6 #(
    .INIT(64'hffff8888ffff8fff)
  ) __177__ (
    .I5(__0__),
    .I4(__11__),
    .I3(__10__),
    .I2(__9__),
    .I1(__7__),
    .I0(__6__),
    .O(__12__)
  );
  LUT3 #(
    .INIT(8'h04)
  ) __178__ (
    .I2(__3__),
    .I1(__1__),
    .I0(__2__),
    .O(__13__)
  );
  LUT5 #(
    .INIT(32'hffee0fff)
  ) __179__ (
    .I4(__4__),
    .I3(__3__),
    .I2(__5__),
    .I1(__2__),
    .I0(v2),
    .O(__14__)
  );
  LUT6 #(
    .INIT(64'h80808080000000ff)
  ) __180__ (
    .I5(__0__),
    .I4(__1__),
    .I3(__14__),
    .I2(__4__),
    .I1(__5__),
    .I0(__13__),
    .O(__15__)
  );
  LUT5 #(
    .INIT(32'heeee0fff)
  ) __181__ (
    .I4(__4__),
    .I3(__2__),
    .I2(v0),
    .I1(__5__),
    .I0(v2),
    .O(__16__)
  );
  LUT6 #(
    .INIT(64'h0a323ffffafaffff)
  ) __182__ (
    .I5(__5__),
    .I4(__1__),
    .I3(__4__),
    .I2(__0__),
    .I1(__2__),
    .I0(__16__),
    .O(__17__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __183__ (
    .I1(__3__),
    .I0(__17__),
    .O(__18__)
  );
  LUT6 #(
    .INIT(64'h00000000fffcf0fa)
  ) __184__ (
    .I5(__4__),
    .I4(__2__),
    .I3(__3__),
    .I2(__5__),
    .I1(v0),
    .I0(__1__),
    .O(__19__)
  );
  LUT5 #(
    .INIT(32'h0000cacc)
  ) __185__ (
    .I4(__2__),
    .I3(__1__),
    .I2(__3__),
    .I1(__4__),
    .I0(v2),
    .O(__20__)
  );
  LUT6 #(
    .INIT(64'h4044f0ff40444044)
  ) __186__ (
    .I5(__2__),
    .I4(__4__),
    .I3(v5),
    .I2(v4),
    .I1(__5__),
    .I0(v2),
    .O(__21__)
  );
  LUT4 #(
    .INIT(16'h30ab)
  ) __187__ (
    .I3(__5__),
    .I2(__2__),
    .I1(__3__),
    .I0(__1__),
    .O(__22__)
  );
  LUT5 #(
    .INIT(32'he8ffffcf)
  ) __188__ (
    .I4(__4__),
    .I3(__1__),
    .I2(__2__),
    .I1(__3__),
    .I0(__5__),
    .O(__23__)
  );
  LUT6 #(
    .INIT(64'h0000fffffefffeff)
  ) __189__ (
    .I5(__0__),
    .I4(__23__),
    .I3(__22__),
    .I2(__21__),
    .I1(__20__),
    .I0(__19__),
    .O(__24__)
  );
  LUT6 #(
    .INIT(64'hf0f3f0faf0f0f0f0)
  ) __190__ (
    .I5(__4__),
    .I4(__5__),
    .I3(__1__),
    .I2(__24__),
    .I1(__2__),
    .I0(__3__),
    .O(__25__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __191__ (
    .I1(__0__),
    .I0(__3__),
    .O(__26__)
  );
  LUT5 #(
    .INIT(32'h0000fdf0)
  ) __192__ (
    .I4(__4__),
    .I3(__2__),
    .I2(__5__),
    .I1(v0),
    .I0(__1__),
    .O(__27__)
  );
  LUT3 #(
    .INIT(8'hf8)
  ) __193__ (
    .I2(__3__),
    .I1(__4__),
    .I0(v2),
    .O(__28__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __194__ (
    .I1(__1__),
    .I0(__2__),
    .O(__29__)
  );
  LUT6 #(
    .INIT(64'h5555555455545555)
  ) __195__ (
    .I5(v5),
    .I4(v4),
    .I3(__29__),
    .I2(__28__),
    .I1(__27__),
    .I0(__0__),
    .O(__30__)
  );
  LUT6 #(
    .INIT(64'hfffffffff1a0ff20)
  ) __196__ (
    .I5(__30__),
    .I4(__5__),
    .I3(__4__),
    .I2(__26__),
    .I1(__1__),
    .I0(__2__),
    .O(__31__)
  );
  LUT3 #(
    .INIT(8'h08)
  ) __198__ (
    .I2(v3),
    .I1(__3__),
    .I0(__1__),
    .O(__33__)
  );
  LUT3 #(
    .INIT(8'h08)
  ) __199__ (
    .I2(__1__),
    .I1(__3__),
    .I0(__2__),
    .O(__34__)
  );
  LUT6 #(
    .INIT(64'h00f0eefe00000000)
  ) __200__ (
    .I5(v2),
    .I4(__4__),
    .I3(v1),
    .I2(__34__),
    .I1(__5__),
    .I0(__33__),
    .O(__35__)
  );
  LUT6 #(
    .INIT(64'h00ff0f0f000f00ef)
  ) __201__ (
    .I5(__1__),
    .I4(__2__),
    .I3(__5__),
    .I2(__3__),
    .I1(v6),
    .I0(v3),
    .O(__36__)
  );
  LUT3 #(
    .INIT(8'h25)
  ) __202__ (
    .I2(__2__),
    .I1(v0),
    .I0(__1__),
    .O(__37__)
  );
  LUT6 #(
    .INIT(64'h000055550000d555)
  ) __203__ (
    .I5(__3__),
    .I4(__4__),
    .I3(v5),
    .I2(v4),
    .I1(__37__),
    .I0(__36__),
    .O(__38__)
  );
  LUT5 #(
    .INIT(32'h0fffffbb)
  ) __204__ (
    .I4(__3__),
    .I3(__5__),
    .I2(__2__),
    .I1(__4__),
    .I0(__1__),
    .O(__39__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __205__ (
    .I1(__2__),
    .I0(__0__),
    .O(__40__)
  );
  LUT6 #(
    .INIT(64'hffff00ff7f7f7f7f)
  ) __206__ (
    .I5(__3__),
    .I4(__1__),
    .I3(v1),
    .I2(__4__),
    .I1(v5),
    .I0(v4),
    .O(__41__)
  );
  LUT6 #(
    .INIT(64'hf0ff7777ffffffff)
  ) __207__ (
    .I5(__4__),
    .I4(__3__),
    .I3(__0__),
    .I2(__5__),
    .I1(__2__),
    .I0(__1__),
    .O(__42__)
  );
  LUT6 #(
    .INIT(64'h000f004400000000)
  ) __208__ (
    .I5(__4__),
    .I4(__3__),
    .I3(__2__),
    .I2(__5__),
    .I1(v3),
    .I0(__1__),
    .O(__43__)
  );
  LUT6 #(
    .INIT(64'h0e0043cc00000000)
  ) __209__ (
    .I5(__0__),
    .I4(__1__),
    .I3(__2__),
    .I2(__3__),
    .I1(__4__),
    .I0(__5__),
    .O(__44__)
  );
  LUT6 #(
    .INIT(64'h000000000000fdf0)
  ) __210__ (
    .I5(__44__),
    .I4(__43__),
    .I3(__42__),
    .I2(v2),
    .I1(__41__),
    .I0(__40__),
    .O(__45__)
  );
  LUT6 #(
    .INIT(64'h00ef0000ffff0000)
  ) __211__ (
    .I5(__45__),
    .I4(CLR),
    .I3(__0__),
    .I2(__39__),
    .I1(__38__),
    .I0(__35__),
    .O(__46__)
  );
  LUT6 #(
    .INIT(64'hfffffffaff0f30ff)
  ) __212__ (
    .I5(__5__),
    .I4(__3__),
    .I3(__1__),
    .I2(__2__),
    .I1(v0),
    .I0(v6),
    .O(__47__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __213__ (
    .I1(__4__),
    .I0(__47__),
    .O(__48__)
  );
  LUT6 #(
    .INIT(64'hffff337ffff0fcff)
  ) __214__ (
    .I5(__2__),
    .I4(__1__),
    .I3(__5__),
    .I2(__3__),
    .I1(__4__),
    .I0(v1),
    .O(__49__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __215__ (
    .I1(v2),
    .I0(__49__),
    .O(__50__)
  );
  LUT3 #(
    .INIT(8'h01)
  ) __216__ (
    .I2(__3__),
    .I1(__2__),
    .I0(__5__),
    .O(__51__)
  );
  LUT6 #(
    .INIT(64'h030000000000000a)
  ) __217__ (
    .I5(__3__),
    .I4(__2__),
    .I3(__4__),
    .I2(v1),
    .I1(v2),
    .I0(__5__),
    .O(__52__)
  );
  LUT5 #(
    .INIT(32'hfffa3fff)
  ) __218__ (
    .I4(__1__),
    .I3(__4__),
    .I2(__5__),
    .I1(__2__),
    .I0(__3__),
    .O(__53__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __219__ (
    .I1(v5),
    .I0(v4),
    .O(__54__)
  );
  LUT6 #(
    .INIT(64'hf3f333fffffff5ff)
  ) __220__ (
    .I5(__3__),
    .I4(__1__),
    .I3(__4__),
    .I2(__2__),
    .I1(__5__),
    .I0(v3),
    .O(__55__)
  );
  LUT6 #(
    .INIT(64'hcdcdcf0000000000)
  ) __221__ (
    .I5(__55__),
    .I4(__54__),
    .I3(__53__),
    .I2(__52__),
    .I1(__1__),
    .I0(__51__),
    .O(__56__)
  );
  LUT6 #(
    .INIT(64'hef03cf0fcf00ffff)
  ) __222__ (
    .I5(__1__),
    .I4(__2__),
    .I3(__3__),
    .I2(__4__),
    .I1(__5__),
    .I0(v2),
    .O(__57__)
  );
  LUT5 #(
    .INIT(32'hfffe30ff)
  ) __223__ (
    .I4(__3__),
    .I3(__4__),
    .I2(v3),
    .I1(__0__),
    .I0(v6),
    .O(__58__)
  );
  LUT5 #(
    .INIT(32'haaa8fffc)
  ) __224__ (
    .I4(__0__),
    .I3(__5__),
    .I2(__1__),
    .I1(__58__),
    .I0(__57__),
    .O(__59__)
  );
  LUT6 #(
    .INIT(64'h00ef0000ffff0000)
  ) __225__ (
    .I5(__59__),
    .I4(CLR),
    .I3(__0__),
    .I2(__56__),
    .I1(__50__),
    .I0(__48__),
    .O(__60__)
  );
  LUT6 #(
    .INIT(64'hff00fcffffffefef)
  ) __226__ (
    .I5(__1__),
    .I4(__3__),
    .I3(__2__),
    .I2(__5__),
    .I1(__4__),
    .I0(v1),
    .O(__61__)
  );
  LUT6 #(
    .INIT(64'ha0aa0a88aaaa08aa)
  ) __227__ (
    .I5(__3__),
    .I4(__2__),
    .I3(__5__),
    .I2(__1__),
    .I1(v6),
    .I0(__61__),
    .O(__62__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __228__ (
    .I1(__3__),
    .I0(v2),
    .O(__63__)
  );
  LUT6 #(
    .INIT(64'hffffffaa00f000c0)
  ) __229__ (
    .I5(__1__),
    .I4(__5__),
    .I3(__3__),
    .I2(__2__),
    .I1(v3),
    .I0(v2),
    .O(__64__)
  );
  LUT6 #(
    .INIT(64'h40fffffffffff0f0)
  ) __230__ (
    .I5(__3__),
    .I4(__2__),
    .I3(v3),
    .I2(v6),
    .I1(v0),
    .I0(v1),
    .O(__65__)
  );
  LUT6 #(
    .INIT(64'h8f0f0000ff0f0000)
  ) __231__ (
    .I5(__65__),
    .I4(__4__),
    .I3(__5__),
    .I2(__64__),
    .I1(__54__),
    .I0(__63__),
    .O(__66__)
  );
  LUT6 #(
    .INIT(64'hf7ffffffffffff0f)
  ) __232__ (
    .I5(__0__),
    .I4(__3__),
    .I3(__1__),
    .I2(__5__),
    .I1(__2__),
    .I0(__4__),
    .O(__67__)
  );
  LUT6 #(
    .INIT(64'hfffbff0ffffff1ff)
  ) __233__ (
    .I5(__4__),
    .I4(__1__),
    .I3(__2__),
    .I2(__3__),
    .I1(__0__),
    .I0(__5__),
    .O(__68__)
  );
  LUT3 #(
    .INIT(8'hb0)
  ) __234__ (
    .I2(__68__),
    .I1(v2),
    .I0(__67__),
    .O(__69__)
  );
  LUT5 #(
    .INIT(32'h0fdf0000)
  ) __235__ (
    .I4(CLR),
    .I3(__0__),
    .I2(__69__),
    .I1(__66__),
    .I0(__62__),
    .O(__70__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __236__ (
    .I1(__3__),
    .I0(v3),
    .O(__71__)
  );
  LUT5 #(
    .INIT(32'h07000000)
  ) __237__ (
    .I4(__5__),
    .I3(__1__),
    .I2(v2),
    .I1(v5),
    .I0(v4),
    .O(__72__)
  );
  LUT5 #(
    .INIT(32'h44f00000)
  ) __238__ (
    .I4(__4__),
    .I3(__5__),
    .I2(__1__),
    .I1(__2__),
    .I0(__3__),
    .O(__73__)
  );
  LUT6 #(
    .INIT(64'hd000000000000000)
  ) __239__ (
    .I5(__2__),
    .I4(__4__),
    .I3(__1__),
    .I2(v0),
    .I1(v1),
    .I0(v6),
    .O(__74__)
  );
  LUT4 #(
    .INIT(16'h0001)
  ) __240__ (
    .I3(__2__),
    .I2(__4__),
    .I1(__5__),
    .I0(__1__),
    .O(__75__)
  );
  LUT6 #(
    .INIT(64'h0f00000000000008)
  ) __241__ (
    .I5(__2__),
    .I4(__5__),
    .I3(__1__),
    .I2(__4__),
    .I1(__3__),
    .I0(v6),
    .O(__76__)
  );
  LUT6 #(
    .INIT(64'h00000000454545cf)
  ) __242__ (
    .I5(__76__),
    .I4(__75__),
    .I3(__74__),
    .I2(__73__),
    .I1(__72__),
    .I0(__71__),
    .O(__77__)
  );
  LUT6 #(
    .INIT(64'h4000000000000000)
  ) __243__ (
    .I5(__3__),
    .I4(__2__),
    .I3(__4__),
    .I2(v6),
    .I1(v3),
    .I0(v1),
    .O(__78__)
  );
  LUT4 #(
    .INIT(16'h0008)
  ) __244__ (
    .I3(__3__),
    .I2(__5__),
    .I1(v5),
    .I0(v4),
    .O(__79__)
  );
  LUT5 #(
    .INIT(32'hf0fe0000)
  ) __245__ (
    .I4(__1__),
    .I3(v0),
    .I2(__51__),
    .I1(__79__),
    .I0(__78__),
    .O(__80__)
  );
  LUT6 #(
    .INIT(64'h0000000000000004)
  ) __246__ (
    .I5(__0__),
    .I4(__3__),
    .I3(__2__),
    .I2(__4__),
    .I1(__5__),
    .I0(__1__),
    .O(__81__)
  );
  LUT4 #(
    .INIT(16'h4000)
  ) __247__ (
    .I3(__2__),
    .I2(__4__),
    .I1(__1__),
    .I0(__5__),
    .O(__82__)
  );
  LUT6 #(
    .INIT(64'hf1fbfbfbfc37ffff)
  ) __248__ (
    .I5(__1__),
    .I4(__0__),
    .I3(__2__),
    .I2(__3__),
    .I1(__4__),
    .I0(__5__),
    .O(__83__)
  );
  LUT6 #(
    .INIT(64'hffff0000007f0000)
  ) __249__ (
    .I5(v2),
    .I4(__83__),
    .I3(__82__),
    .I2(v1),
    .I1(v6),
    .I0(__81__),
    .O(__84__)
  );
  LUT5 #(
    .INIT(32'h0fdf0000)
  ) __250__ (
    .I4(CLR),
    .I3(__0__),
    .I2(__84__),
    .I1(__80__),
    .I0(__77__),
    .O(__85__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __251__ (
    .I1(__5__),
    .I0(__1__),
    .O(__86__)
  );
  LUT6 #(
    .INIT(64'hfffff0ff0fff5f13)
  ) __252__ (
    .I5(__3__),
    .I4(__5__),
    .I3(__1__),
    .I2(__2__),
    .I1(__54__),
    .I0(v0),
    .O(__87__)
  );
  LUT6 #(
    .INIT(64'hf0ffffff11155555)
  ) __253__ (
    .I5(__3__),
    .I4(__2__),
    .I3(__1__),
    .I2(__5__),
    .I1(v2),
    .I0(__0__),
    .O(__88__)
  );
  LUT6 #(
    .INIT(64'h0000ffff888f888f)
  ) __254__ (
    .I5(__4__),
    .I4(__88__),
    .I3(__0__),
    .I2(__87__),
    .I1(__7__),
    .I0(__86__),
    .O(__89__)
  );
  LUT3 #(
    .INIT(8'he8)
  ) __255__ (
    .I2(__3__),
    .I1(__5__),
    .I0(__1__),
    .O(__90__)
  );
  LUT5 #(
    .INIT(32'hff0f111f)
  ) __256__ (
    .I4(__3__),
    .I3(__5__),
    .I2(__1__),
    .I1(__0__),
    .I0(v2),
    .O(__91__)
  );
  LUT5 #(
    .INIT(32'hf3f350ff)
  ) __257__ (
    .I4(__2__),
    .I3(__1__),
    .I2(__4__),
    .I1(v0),
    .I0(v2),
    .O(__92__)
  );
  LUT6 #(
    .INIT(64'ha003000000000000)
  ) __258__ (
    .I5(v5),
    .I4(v4),
    .I3(__4__),
    .I2(__5__),
    .I1(__0__),
    .I0(__2__),
    .O(__93__)
  );
  LUT4 #(
    .INIT(16'h4100)
  ) __259__ (
    .I3(__2__),
    .I2(__5__),
    .I1(__1__),
    .I0(__4__),
    .O(__94__)
  );
  LUT6 #(
    .INIT(64'h00000000ffffff01)
  ) __260__ (
    .I5(__3__),
    .I4(__94__),
    .I3(__93__),
    .I2(__0__),
    .I1(__5__),
    .I0(__92__),
    .O(__95__)
  );
  LUT6 #(
    .INIT(64'hff0fff44ff00ff00)
  ) __261__ (
    .I5(__4__),
    .I4(__2__),
    .I3(__95__),
    .I2(__91__),
    .I1(__0__),
    .I0(__90__),
    .O(__96__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __262__ (
    .I1(__3__),
    .I0(__2__),
    .O(__97__)
  );
  LUT4 #(
    .INIT(16'h0037)
  ) __263__ (
    .I3(__5__),
    .I2(__2__),
    .I1(__1__),
    .I0(v2),
    .O(__98__)
  );
  LUT6 #(
    .INIT(64'h000000008acf8a8a)
  ) __264__ (
    .I5(__98__),
    .I4(__54__),
    .I3(__97__),
    .I2(__5__),
    .I1(__65__),
    .I0(__1__),
    .O(__99__)
  );
  LUT5 #(
    .INIT(32'h000f0088)
  ) __265__ (
    .I4(__3__),
    .I3(v3),
    .I2(__1__),
    .I1(__4__),
    .I0(__5__),
    .O(__100__)
  );
  LUT5 #(
    .INIT(32'h00000008)
  ) __266__ (
    .I4(__3__),
    .I3(__5__),
    .I2(__1__),
    .I1(v5),
    .I0(v4),
    .O(__101__)
  );
  LUT5 #(
    .INIT(32'h02300000)
  ) __267__ (
    .I4(v2),
    .I3(__1__),
    .I2(__4__),
    .I1(__3__),
    .I0(__5__),
    .O(__102__)
  );
  LUT6 #(
    .INIT(64'h003000ce00000000)
  ) __268__ (
    .I5(__3__),
    .I4(__1__),
    .I3(__4__),
    .I2(__2__),
    .I1(__5__),
    .I0(v6),
    .O(__103__)
  );
  LUT5 #(
    .INIT(32'h000000f1)
  ) __269__ (
    .I4(__103__),
    .I3(__102__),
    .I2(__2__),
    .I1(__101__),
    .I0(__100__),
    .O(__104__)
  );
  LUT6 #(
    .INIT(64'hf7f7f7f7cf30ffff)
  ) __270__ (
    .I5(__2__),
    .I4(__4__),
    .I3(__1__),
    .I2(__3__),
    .I1(__5__),
    .I0(__0__),
    .O(__105__)
  );
  LUT6 #(
    .INIT(64'h00ff4fff00000000)
  ) __271__ (
    .I5(CLR),
    .I4(__0__),
    .I3(__105__),
    .I2(__104__),
    .I1(__4__),
    .I0(__99__),
    .O(__106__)
  );
  LUT6 #(
    .INIT(64'h00ff0000ffbfffff)
  ) __272__ (
    .I5(__5__),
    .I4(__1__),
    .I3(__3__),
    .I2(v5),
    .I1(v4),
    .I0(v0),
    .O(__107__)
  );
  LUT6 #(
    .INIT(64'h005500a0005500b0)
  ) __273__ (
    .I5(__3__),
    .I4(__2__),
    .I3(__4__),
    .I2(__5__),
    .I1(v6),
    .I0(__107__),
    .O(__108__)
  );
  LUT6 #(
    .INIT(64'hf000fffff0f0ff88)
  ) __274__ (
    .I5(__4__),
    .I4(__3__),
    .I3(__2__),
    .I2(__1__),
    .I1(v1),
    .I0(v3),
    .O(__109__)
  );
  LUT6 #(
    .INIT(64'h4fff00ff00000000)
  ) __275__ (
    .I5(__5__),
    .I4(__97__),
    .I3(__109__),
    .I2(v3),
    .I1(v6),
    .I0(v1),
    .O(__110__)
  );
  LUT4 #(
    .INIT(16'h4000)
  ) __276__ (
    .I3(__0__),
    .I2(__3__),
    .I1(__4__),
    .I0(__5__),
    .O(__111__)
  );
  LUT3 #(
    .INIT(8'h04)
  ) __277__ (
    .I2(__0__),
    .I1(__5__),
    .I0(__3__),
    .O(__112__)
  );
  LUT6 #(
    .INIT(64'h00000000eccfcccc)
  ) __278__ (
    .I5(v2),
    .I4(__112__),
    .I3(__2__),
    .I2(__4__),
    .I1(__111__),
    .I0(__54__),
    .O(__113__)
  );
  LUT6 #(
    .INIT(64'h1170000000000000)
  ) __279__ (
    .I5(__0__),
    .I4(__4__),
    .I3(__5__),
    .I2(__3__),
    .I1(__2__),
    .I0(__1__),
    .O(__114__)
  );
  LUT6 #(
    .INIT(64'hff00ff00ff000e00)
  ) __280__ (
    .I5(__114__),
    .I4(__113__),
    .I3(CLR),
    .I2(__0__),
    .I1(__110__),
    .I0(__108__),
    .O(__115__)
  );
  LUT4 #(
    .INIT(16'h0004)
  ) __281__ (
    .I3(__0__),
    .I2(__3__),
    .I1(v4),
    .I0(v5),
    .O(__116__)
  );
  LUT6 #(
    .INIT(64'h440000f000000000)
  ) __282__ (
    .I5(__116__),
    .I4(__4__),
    .I3(__5__),
    .I2(__37__),
    .I1(__2__),
    .I0(v2),
    .O(__117__)
  );
  LUT3 #(
    .INIT(8'h01)
  ) __283__ (
    .I2(__0__),
    .I1(__3__),
    .I0(__1__),
    .O(__118__)
  );
  LUT6 #(
    .INIT(64'hf000004400000000)
  ) __284__ (
    .I5(__118__),
    .I4(__4__),
    .I3(__5__),
    .I2(v2),
    .I1(__54__),
    .I0(__2__),
    .O(__119__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __286__ (
    .I1(__1__),
    .I0(__0__),
    .O(__121__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __287__ (
    .I1(__4__),
    .I0(__5__),
    .O(__122__)
  );
  LUT6 #(
    .INIT(64'hd000000000000000)
  ) __288__ (
    .I5(__122__),
    .I4(v3),
    .I3(__97__),
    .I2(__121__),
    .I1(v1),
    .I0(v6),
    .O(__123__)
  );
  LUT5 #(
    .INIT(32'hfffe7fff)
  ) __289__ (
    .I4(__3__),
    .I3(__4__),
    .I2(__5__),
    .I1(__1__),
    .I0(v6),
    .O(__124__)
  );
  LUT6 #(
    .INIT(64'h4000000000000000)
  ) __290__ (
    .I5(__0__),
    .I4(__3__),
    .I3(__2__),
    .I2(__4__),
    .I1(__1__),
    .I0(__5__),
    .O(__125__)
  );
  LUT6 #(
    .INIT(64'hffff010001000100)
  ) __291__ (
    .I5(v2),
    .I4(__125__),
    .I3(v3),
    .I2(__0__),
    .I1(__2__),
    .I0(__124__),
    .O(__126__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __292__ (
    .I1(__5__),
    .I0(v2),
    .O(__127__)
  );
  LUT3 #(
    .INIT(8'h0d)
  ) __293__ (
    .I2(__1__),
    .I1(v4),
    .I0(v5),
    .O(__128__)
  );
  LUT6 #(
    .INIT(64'h5500fdfc5500fcfc)
  ) __294__ (
    .I5(__98__),
    .I4(__2__),
    .I3(__4__),
    .I2(__3__),
    .I1(__128__),
    .I0(__127__),
    .O(__129__)
  );
  LUT5 #(
    .INIT(32'hcc04cccc)
  ) __295__ (
    .I4(__2__),
    .I3(__3__),
    .I2(__4__),
    .I1(__5__),
    .I0(__1__),
    .O(__130__)
  );
  LUT5 #(
    .INIT(32'h1e030000)
  ) __296__ (
    .I4(__4__),
    .I3(__3__),
    .I2(__5__),
    .I1(__1__),
    .I0(__2__),
    .O(__131__)
  );
  LUT6 #(
    .INIT(64'hffffffff0f0f0f08)
  ) __297__ (
    .I5(__131__),
    .I4(__130__),
    .I3(__129__),
    .I2(__0__),
    .I1(__3__),
    .I0(__1__),
    .O(__132__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __298__ (
    .I1(__2__),
    .I0(__1__),
    .O(__133__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __299__ (
    .I1(__0__),
    .I0(__4__),
    .O(__134__)
  );
  LUT6 #(
    .INIT(64'h2000750000000000)
  ) __300__ (
    .I5(__0__),
    .I4(__3__),
    .I3(__2__),
    .I2(__4__),
    .I1(__5__),
    .I0(__1__),
    .O(__135__)
  );
  LUT6 #(
    .INIT(64'h000f33ff0303fbf3)
  ) __301__ (
    .I5(__5__),
    .I4(__4__),
    .I3(__2__),
    .I2(__0__),
    .I1(__1__),
    .I0(v0),
    .O(__136__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __302__ (
    .I1(__3__),
    .I0(__136__),
    .O(__137__)
  );
  LUT6 #(
    .INIT(64'hffffff8080808080)
  ) __303__ (
    .I5(v2),
    .I4(__137__),
    .I3(__135__),
    .I2(__134__),
    .I1(__79__),
    .I0(__133__),
    .O(__138__)
  );
  LUT6 #(
    .INIT(64'hf5ffffffffffff3f)
  ) __304__ (
    .I5(__0__),
    .I4(__3__),
    .I3(__2__),
    .I2(__5__),
    .I1(__8__),
    .I0(v2),
    .O(__139__)
  );
  LUT3 #(
    .INIT(8'h08)
  ) __305__ (
    .I2(__139__),
    .I1(__4__),
    .I0(__1__),
    .O(__140__)
  );
  LUT6 #(
    .INIT(64'hfffff0ffffbbffff)
  ) __306__ (
    .I5(__0__),
    .I4(__1__),
    .I3(__4__),
    .I2(v2),
    .I1(__2__),
    .I0(v5),
    .O(__141__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __307__ (
    .I1(__3__),
    .I0(__5__),
    .O(__142__)
  );
  LUT5 #(
    .INIT(32'hff3faeff)
  ) __308__ (
    .I4(__3__),
    .I3(__5__),
    .I2(__1__),
    .I1(__0__),
    .I0(v5),
    .O(__143__)
  );
  LUT6 #(
    .INIT(64'h0ee0eeeeff00ffff)
  ) __309__ (
    .I5(__4__),
    .I4(__26__),
    .I3(__1__),
    .I2(__5__),
    .I1(v2),
    .I0(__143__),
    .O(__144__)
  );
  LUT6 #(
    .INIT(64'h0003030000000001)
  ) __310__ (
    .I5(__3__),
    .I4(__2__),
    .I3(__1__),
    .I2(__4__),
    .I1(__5__),
    .I0(v5),
    .O(__145__)
  );
  LUT6 #(
    .INIT(64'h00000000ff80ff00)
  ) __311__ (
    .I5(__0__),
    .I4(__4__),
    .I3(__145__),
    .I2(__5__),
    .I1(__13__),
    .I0(__8__),
    .O(__146__)
  );
  LUT6 #(
    .INIT(64'hffffffff10ff1010)
  ) __312__ (
    .I5(__146__),
    .I4(__2__),
    .I3(__144__),
    .I2(__142__),
    .I1(v0),
    .I0(__141__),
    .O(__147__)
  );
  LUT6 #(
    .INIT(64'h0ffffff5f3ffffff)
  ) __313__ (
    .I5(__3__),
    .I4(__2__),
    .I3(__1__),
    .I2(__5__),
    .I1(v0),
    .I0(v6),
    .O(__148__)
  );
  LUT3 #(
    .INIT(8'h01)
  ) __314__ (
    .I2(__0__),
    .I1(__4__),
    .I0(__148__),
    .O(__149__)
  );
  LUT6 #(
    .INIT(64'hff0fffff33f2fffa)
  ) __315__ (
    .I5(__5__),
    .I4(__2__),
    .I3(__3__),
    .I2(v1),
    .I1(__4__),
    .I0(__0__),
    .O(__150__)
  );
  LUT5 #(
    .INIT(32'h0fffffd0)
  ) __316__ (
    .I4(__4__),
    .I3(__5__),
    .I2(__2__),
    .I1(v0),
    .I0(__1__),
    .O(__151__)
  );
  LUT5 #(
    .INIT(32'he0000000)
  ) __317__ (
    .I4(__2__),
    .I3(__4__),
    .I2(v2),
    .I1(__5__),
    .I0(__1__),
    .O(__152__)
  );
  LUT5 #(
    .INIT(32'hfffbf8ff)
  ) __318__ (
    .I4(__2__),
    .I3(__1__),
    .I2(__5__),
    .I1(__3__),
    .I0(__4__),
    .O(__153__)
  );
  LUT6 #(
    .INIT(64'h0000000000fff4ff)
  ) __319__ (
    .I5(__0__),
    .I4(__3__),
    .I3(__153__),
    .I2(__152__),
    .I1(__54__),
    .I0(__151__),
    .O(__154__)
  );
  LUT6 #(
    .INIT(64'h0040150c00000000)
  ) __320__ (
    .I5(__0__),
    .I4(__1__),
    .I3(__2__),
    .I2(__5__),
    .I1(__4__),
    .I0(__3__),
    .O(__155__)
  );
  LUT4 #(
    .INIT(16'hfff2)
  ) __321__ (
    .I3(__155__),
    .I2(__154__),
    .I1(__150__),
    .I0(__1__),
    .O(__156__)
  );
  LUT5 #(
    .INIT(32'hf0ffffbb)
  ) __322__ (
    .I4(__4__),
    .I3(__5__),
    .I2(v2),
    .I1(__1__),
    .I0(v0),
    .O(__157__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __323__ (
    .I1(__0__),
    .I0(__3__),
    .O(__158__)
  );
  LUT6 #(
    .INIT(64'h8f0c880000000000)
  ) __324__ (
    .I5(__158__),
    .I4(__2__),
    .I3(v5),
    .I2(__157__),
    .I1(v4),
    .I0(__75__),
    .O(__159__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __325__ (
    .I1(v5),
    .I0(v4),
    .O(__160__)
  );
  LUT6 #(
    .INIT(64'hbbbbfffffffff0ff)
  ) __326__ (
    .I5(__4__),
    .I4(__5__),
    .I3(__1__),
    .I2(v0),
    .I1(__2__),
    .I0(v2),
    .O(__161__)
  );
  LUT6 #(
    .INIT(64'h0003000000000b00)
  ) __327__ (
    .I5(__3__),
    .I4(__2__),
    .I3(__1__),
    .I2(__5__),
    .I1(__4__),
    .I0(v2),
    .O(__162__)
  );
  LUT5 #(
    .INIT(32'hffef731f)
  ) __328__ (
    .I4(__3__),
    .I3(__2__),
    .I2(__4__),
    .I1(__5__),
    .I0(__1__),
    .O(__163__)
  );
  LUT6 #(
    .INIT(64'h0000ffffff01ff01)
  ) __329__ (
    .I5(__0__),
    .I4(__163__),
    .I3(__162__),
    .I2(__3__),
    .I1(__161__),
    .I0(__160__),
    .O(__164__)
  );
  assign v13_D_9 = __18__;
  assign v13_D_24 = __147__;
  assign v13_D_15 = __117__;
  assign v13_D_21 = __119__;
  assign v13_D_10 = __96__;
  assign v13_D_13 = __156__;
  assign v13_D_17 = __138__;
  assign v13_D_22 = __15__;
  assign v13_D_20 = __123__;
  assign v13_D_16 = __140__;
  assign v13_D_19 = __126__;
  assign v13_D_6 = __132__;
  assign v13_D_8 = __25__;
  assign v13_D_18 = __159__;
  assign v13_D_14 = __31__;
  assign v13_D_12 = __89__;
  assign v13_D_23 = __149__;
  assign v13_D_11 = __12__;
  assign v13_D_7 = __164__;
endmodule
