// IWLS benchmark module "s953.bench" printed on Wed May 29 21:45:20 2002
module s953 (Rdy1RtHS1, Rdy2RtHS1, Rdy1BmHS1, Rdy2BmHS1, IInDoneHS1, RtTSHS1, TpArrayHS1, OutputHS1, WantBmHS1, WantRtHS1, OutAvHS1, FullOHS1, FullIIHS1, Prog_2, Prog_1, Prog_0, ReWhBufHS1, TgWhBufHS1, SeOutAvHS1, LdProgHS1, Mode2HS1, ReRtTSHS1, ShftIIRHS1, NewTrHS1, Mode1HS1, ShftORHS1, ActRtHS1, Mode0HS1, TxHIInHS1, LxHIInHS1, NewLineHS1, ActBmHS1, GoBmHS1, LoadOHHS1, DumpIIHS1, SeFullOHS1, GoRtHS1, LoadIIHHS1, SeFullIIHS1);
input
  WantBmHS1,
  IInDoneHS1,
  WantRtHS1,
  Prog_0,
  Prog_1,
  Prog_2,
  Rdy2BmHS1,
  FullIIHS1,
  OutAvHS1,
  Rdy2RtHS1,
  TpArrayHS1,
  RtTSHS1,
  FullOHS1,
  Rdy1BmHS1,
  Rdy1RtHS1,
  OutputHS1;
output
  LoadOHHS1,
  GoBmHS1,
  GoRtHS1,
  SeFullIIHS1,
  LxHIInHS1,
  ReWhBufHS1,
  NewTrHS1,
  SeFullOHS1,
  Mode0HS1,
  ShftIIRHS1,
  Mode1HS1,
  Mode2HS1,
  LoadIIHHS1,
  ActBmHS1,
  ActRtHS1,
  TxHIInHS1,
  TgWhBufHS1,
  SeOutAvHS1,
  DumpIIHS1,
  LdProgHS1,
  ReRtTSHS1,
  NewLineHS1,
  ShftORHS1;
reg
  \[8373] ,
  \[8374] ,
  \[8375] ,
  \[8376] ,
  \[8377] ,
  \[8378] ,
  \[8379] ,
  \[8380] ,
  \[8381] ,
  \[8382] ,
  \[8383] ,
  \[8384] ,
  \[8385] ,
  \[8386] ,
  \[8387] ,
  \[8388] ,
  \[8389] ,
  \[8390] ,
  \[8391] ,
  \[8392] ,
  \[8393] ,
  \[8394] ,
  \[8395] ,
  State_0,
  State_1,
  State_2,
  State_3,
  State_4,
  State_5;
wire
  II829_1,
  \[77] ,
  \[78] ,
  II857_1,
  \[79] ,
  \[80] ,
  II1037_1,
  II2,
  II3,
  II4,
  II5,
  II6,
  II7,
  II8,
  II9,
  II1028_1,
  II1188_1,
  II1188_2,
  II910_1,
  II1143_1,
  II1143_2,
  II1047_1,
  II1047_2,
  II896_1,
  II1125_1,
  II1163_1,
  II1199_1,
  II1199_2,
  II1100_1,
  II263,
  II264,
  II265,
  II266,
  II267,
  II269,
  II271,
  II272,
  II274,
  II275,
  II276,
  II277,
  II278,
  II279,
  II280,
  II281,
  II282,
  II283,
  II284,
  II1154_1,
  II287,
  II294,
  II295,
  II297,
  II1173_1,
  II300,
  II303,
  II1110_1,
  II1077_1,
  II311,
  II315,
  II317,
  II318,
  II1136_1,
  II320,
  II322,
  II323,
  II325,
  II326,
  II327,
  II328,
  II329,
  II330,
  II331,
  II333,
  II335,
  II336,
  II338,
  II339,
  II340,
  II341,
  II342,
  II343,
  II344,
  II345,
  II347,
  II348,
  II350,
  II351,
  II353,
  II354,
  II355,
  II357,
  II358,
  II359,
  II360,
  II362,
  II363,
  II364,
  II366,
  II367,
  II370,
  II371,
  II372,
  II374,
  II376,
  II377,
  II378,
  II379,
  II380,
  II381,
  II382,
  II384,
  II386,
  II388,
  II390,
  II391,
  II393,
  II394,
  II396,
  II397,
  II398,
  II399,
  II1087_1,
  II403,
  II10,
  II404,
  II11,
  II405,
  II12,
  II13,
  II407,
  II14,
  II408,
  II15,
  II16,
  II17,
  II18,
  II19,
  II410,
  II411,
  II412,
  II20,
  II414,
  II21,
  II415,
  II22,
  II416,
  II23,
  II24,
  II418,
  II25,
  II26,
  II27,
  II28,
  II29,
  II421,
  II422,
  II423,
  II30,
  II424,
  II425,
  II428,
  II429,
  II430,
  II431,
  II432,
  II434,
  II435,
  II436,
  II437,
  II439,
  II440,
  II441,
  II442,
  II444,
  II445,
  II446,
  II447,
  II449,
  II450,
  II451,
  II1193_1,
  II452,
  II453,
  II455,
  II457,
  II458,
  II459,
  II461,
  II463,
  II465,
  II466,
  II467,
  II468,
  II469,
  II1097_1,
  II470,
  II473,
  II474,
  II475,
  II476,
  II477,
  II479,
  II481,
  II482,
  II485,
  II486,
  II487,
  II489,
  II491,
  II493,
  II494,
  II495,
  II497,
  II498,
  II1184_1,
  II1184_2,
  II1121_1,
  II1121_2,
  II810_1,
  II500,
  II503,
  II504,
  II505,
  II506,
  II508,
  II509,
  II511,
  II512,
  II513,
  II514,
  II517,
  II519,
  II1140_1,
  II521,
  II523,
  II525,
  II526,
  II796_1,
  II529,
  II531,
  II532,
  II534,
  II535,
  II1207_1,
  II537,
  II1166_1,
  II539,
  II1166_2,
  II1034_1,
  II540,
  II543,
  II545,
  II547,
  II548,
  II551,
  II552,
  II553,
  II554,
  II555,
  II556,
  II559,
  II561,
  II562,
  II565,
  II566,
  II567,
  II568,
  II570,
  II571,
  II573,
  II575,
  II577,
  II579,
  II580,
  II582,
  II585,
  II587,
  II589,
  II1025_1,
  II590,
  II593,
  II595,
  II596,
  II599,
  II1176_1,
  II1176_2,
  II1044_1,
  II600,
  II609,
  II610,
  II612,
  II614,
  II624,
  II625,
  II634,
  II655,
  II657,
  II659,
  II660,
  II661,
  II662,
  II663,
  II665,
  II667,
  II669,
  II1132_1,
  II1132_2,
  II671,
  II673,
  II675,
  II676,
  II678,
  II680,
  II682,
  II684,
  II1160_1,
  II686,
  II689,
  II690,
  II691,
  II693,
  II695,
  II697,
  II699,
  II1151_1,
  II840_1,
  II840_2,
  II700,
  II702,
  II704,
  II706,
  II708,
  II711,
  II713,
  II715,
  II717,
  II719,
  II721,
  II963_1,
  II723,
  II725,
  II729,
  II731,
  II733,
  II735,
  II737,
  II738,
  II1170_1,
  II740,
  II742,
  II744,
  II746,
  II750,
  II1196_1,
  II767,
  II768,
  II769,
  II770,
  II771,
  II789_1,
  II777,
  II778,
  II779,
  II850_1,
  II850_2,
  II1083_1,
  II1180_1,
  II1180_2,
  II1056_1,
  II814_1,
  II1203_1,
  II1203_2,
  II1040_1,
  II861_1,
  II861_2,
  II1107_1,
  II1094_1,
  II1031_1,
  \[29] ,
  II1213_1,
  \[30] ,
  \[31] ,
  II966_1,
  \[32] ,
  II834_1,
  \[33] ,
  \[34] ,
  \[35] ,
  \[36] ,
  \[37] ,
  \[38] ,
  \[39] ,
  II881_1,
  II881_2,
  \[40] ,
  II1118_1,
  \[41] ,
  \[42] ,
  \[43] ,
  \[44] ,
  \[45] ,
  \[46] ,
  \[47] ,
  \[48] ,
  \[49] ,
  II1128_1,
  II873_1,
  \[50] ,
  II1080_1,
  \[51] ,
  \[52] ,
  \[53] ,
  \[54] ,
  \[55] ,
  II892_1,
  II892_2,
  \[56] ,
  \[57] ,
  \[58] ,
  \[59] ,
  II1157_1,
  II1216_1,
  II1216_2,
  \[60] ,
  \[61] ,
  II1148_1,
  \[62] ,
  \[63] ,
  \[64] ,
  II1103_1,
  \[65] ,
  II1103_2,
  \[66] ,
  \[67] ,
  \[68] ,
  \[69] ,
  II1091_1,
  \[70] ,
  II1113_1,
  \[71] ,
  \[72] ,
  \[73] ,
  II1210_1,
  \[74] ,
  \[75] ,
  \[76] ;
assign
  II829_1 = II575 | II547,
  \[77]  = II27,
  \[78]  = II28,
  II857_1 = II493 | Prog_0,
  \[79]  = II29,
  \[80]  = II30,
  II1037_1 = II336 | Prog_0,
  LoadOHHS1 = \[46] ,
  II2 = ~II769 | (~II771 | ~II711),
  II3 = ~II723 | ~II721,
  II4 = ~II551 | (~II381 | ~II725),
  II5 = ~II397 | (~II731 | (~II729 | ~II733)),
  II6 = ~II777 | (~II779 | ~II377),
  II7 = ~II311,
  II8 = ~II657 | ~II655,
  II9 = ~II659 | (~II661 | ~II377),
  II1028_1 = II493 | II367,
  II1188_1 = II376 & State_1,
  II1188_2 = II388 & II267,
  II910_1 = II360 & II277,
  GoBmHS1 = \[45] ,
  II1143_1 = II404 & II353,
  II1143_2 = II596 & II274,
  II1047_1 = II284 | II264,
  II1047_2 = Prog_0 | Rdy1BmHS1,
  GoRtHS1 = \[49] ,
  II896_1 = II320 | II279,
  II1125_1 = II561 | Rdy2RtHS1,
  SeFullIIHS1 = \[51] ,
  II1163_1 = II531 & II345,
  II1199_1 = II364 & II338,
  II1199_2 = II380 & II267,
  II1100_1 = II384 & WantBmHS1,
  II263 = ~Rdy1RtHS1,
  II264 = ~Rdy2RtHS1,
  II265 = ~Rdy1BmHS1,
  II266 = ~Rdy2BmHS1,
  II267 = ~IInDoneHS1,
  II269 = ~TpArrayHS1,
  II271 = ~WantBmHS1,
  II272 = ~WantRtHS1,
  II274 = ~FullOHS1,
  II275 = ~FullIIHS1,
  II276 = ~State_5,
  II277 = ~State_4,
  II278 = ~State_3,
  LxHIInHS1 = \[42] ,
  II279 = ~State_2,
  II280 = ~State_1,
  II281 = ~State_0,
  II282 = ~Prog_2,
  II283 = ~Prog_1,
  II284 = ~Prog_0,
  II1154_1 = II371 | II267,
  II287 = ~II789_1 & ~II750,
  II294 = ~II676 & (~II678 & ~II408),
  II295 = ~II680 & (~II682 & ~II376),
  II297 = ~II684 & (~II686 & ~II376),
  II1173_1 = II466 & II263,
  II300 = ~II810_1 & ~II700,
  II303 = ~II708 & ~II706,
  II1110_1 = II388 & II277,
  II1077_1 = II512 & II458,
  II311 = ~II744 & (~II746 & ~II742),
  II315 = ~II514 & ~II272,
  II317 = ~FullIIHS1 | ~FullOHS1,
  II318 = ~II277 | ~II834_1,
  II1136_1 = II590 & II282,
  II320 = ~II511 | ~II495,
  II322 = ~II323,
  II323 = ~II436 | (~II281 | ~State_4),
  II325 = ~II840_2 & ~II840_1,
  II326 = ~FullIIHS1 & ~FullOHS1,
  II327 = ~II326,
  II328 = ~II539 & (~II511 & ~II609),
  II329 = ~II328,
  II330 = ~II493 | ~WantBmHS1,
  II331 = ~II330,
  II333 = ~II850_2 & ~II850_1,
  II335 = ~II282 | ~II277,
  II336 = ~II357 | ~II473,
  II338 = ~II439 | ~II857_1,
  II339 = ~II338,
  II340 = ~II861_2 | ~II861_1,
  II341 = ~II340,
  II342 = ~II343,
  II343 = ~II482 | (~II394 | ~II276),
  II344 = ~II345,
  II345 = ~Rdy2RtHS1 | ~Rdy1RtHS1,
  II347 = ~II394 & ~State_3,
  II348 = ~II363 & ~II315,
  II350 = ~II477 & ~II325,
  II351 = ~II350,
  II353 = ~II873_1 & ~II344,
  II354 = ~II543 & ~II367,
  II355 = ~II354,
  II357 = ~Rdy2BmHS1 | ~Rdy1BmHS1,
  II358 = ~II359,
  II359 = ~II532 | (~II432 | ~Rdy1RtHS1),
  II360 = ~II881_2 | ~II881_1,
  II362 = ~II407 & ~State_0,
  II363 = ~II362,
  II364 = ~II525 & (~II379 & ~II274),
  II366 = ~II399 & (~II335 & ~State_0),
  ReWhBufHS1 = \[29] ,
  II367 = ~II366,
  II370 = ~II371,
  II371 = ~II382 | ~II279,
  II372 = ~II892_2 | ~II892_1,
  II374 = ~II461 | ~II896_1,
  II376 = ~II479 & ~II281,
  II377 = ~II376,
  II378 = ~II431 & ~FullIIHS1,
  II379 = ~II378,
  II380 = ~II381,
  II381 = ~II396 | ~State_3,
  II382 = ~II485 & (~Prog_2 & ~II276),
  II384 = ~II493 & (~II407 & ~II315),
  II386 = ~II280 & ~State_2,
  II388 = ~II459 & ~II320,
  II390 = ~II391,
  II391 = ~II910_1 & ~State_2,
  II393 = ~II283 | ~II282,
  II394 = ~II357 & (~II327 & ~State_0),
  II396 = ~II425 & ~II280,
  II397 = ~II396,
  II398 = ~II399,
  II399 = ~II436 | ~II284,
  II1087_1 = II526 | Prog_0,
  II403 = ~II494 | (~II434 | ~II634),
  II10 = ~II287,
  II404 = ~II421 & ~II284,
  II11 = ~II667 | (~II669 | ~II475),
  II405 = ~II404,
  II12 = ~II469 | ~II377,
  II13 = ~II415,
  II407 = ~II532 | ~II412,
  II14 = ~II673 | ~II671,
  II408 = ~II523 & (~II435 & ~II341),
  II15 = ~II675 | ~II796_1,
  II16 = ~II323,
  II17 = ~II294,
  II18 = ~II295,
  II19 = ~II323 | ~II371,
  II410 = ~II411,
  II411 = ~II416 | (~Prog_0 | ~II279),
  II412 = ~II437 & ~II282,
  II20 = ~II297,
  II414 = ~II521 & (~II425 & ~State_1),
  II21 = ~II691 | (~II693 | ~II689),
  II415 = ~II414,
  II22 = ~II481 | (~II697 | (~II695 | ~II699)),
  II416 = ~II535 & ~II461,
  II23 = ~II300,
  II24 = ~II326 & ~OutAvHS1,
  II418 = ~II485 & ~II279,
  II25 = ~II767 | ~II814_1,
  II26 = ~II303,
  II27 = ~II275 & ~OutAvHS1,
  II28 = ~FullIIHS1 & ~OutAvHS1,
  II29 = ~II441 & (~State_2 & ~II278),
  II421 = ~II422 | ~II274,
  II422 = ~II525 & ~II431,
  II423 = ~II422,
  II30 = ~II351 | ~II829_1,
  II424 = ~II425,
  II425 = ~II508 | (~II281 | ~State_2),
  II428 = ~II429,
  II429 = ~II450 | ~Prog_0,
  II430 = ~II451 & ~Prog_2,
  II431 = ~II430,
  II432 = ~II451 & ~II282,
  II434 = ~II503 & ~FullIIHS1,
  II435 = ~II434,
  II436 = ~II505 & ~State_1,
  II437 = ~II436,
  II439 = ~II514 | ~Prog_0,
  II440 = ~II509 & ~II495,
  II441 = ~II440,
  II442 = ~II509 & (~II347 & ~State_1),
  II444 = ~II445,
  II445 = ~II534 | ~II374,
  II446 = ~II447,
  II447 = ~II362 | ~Rdy2RtHS1,
  II449 = ~II450 | (~II318 | ~State_1),
  II450 = ~II505 & ~State_0,
  II451 = ~II450,
  II1193_1 = II521 & II424,
  II452 = ~II453,
  II453 = ~II504 | (~II327 | ~II277),
  II455 = ~II512 | ~II264,
  II457 = ~II506 | ~II266,
  II458 = ~II571 & ~II279,
  II459 = ~II458,
  II461 = ~II506 | ~II282,
  II463 = ~II963_1 & ~II390,
  II465 = ~II966_1 & ~II390,
  II466 = ~II503 & ~Rdy1BmHS1,
  II467 = ~II466,
  II468 = ~II487 & (~II386 & ~State_0),
  II469 = ~II468,
  II1097_1 = II556 & II317,
  II470 = ~II571 & (~II335 & ~II320),
  II473 = ~II266 | ~II265,
  II474 = ~II577 & ~II493,
  II475 = ~II474,
  II476 = ~II545 & ~II519,
  II477 = ~II476,
  II479 = ~II486 | ~II279,
  II481 = ~II486 | ~II372,
  II482 = ~II525 & (~State_2 & ~State_3),
  II485 = ~II548 | ~II277,
  II486 = ~II487,
  II487 = ~II508 | ~State_3,
  II489 = ~II570 | ~II506,
  II491 = ~II548 | ~State_5,
  II493 = ~II266 | ~Rdy1BmHS1,
  II494 = ~II495,
  II495 = ~II281 | ~II280,
  II497 = ~II457 | ~II455,
  II498 = ~II473 & ~II271,
  II1184_1 = II506 & II486,
  II1184_2 = II376 & II269,
  II1121_1 = II589 | State_0,
  II1121_2 = II559 | Rdy2BmHS1,
  II810_1 = II562 & II364,
  II500 = ~II453 & ~II281,
  II503 = ~II504 | ~II277,
  II504 = ~II505,
  II505 = ~II570 | ~II279,
  II506 = ~II281 & ~State_1,
  II508 = ~II509,
  II509 = ~II277 | ~II276,
  II511 = ~State_0 | ~State_1,
  II512 = ~State_0 & ~II280,
  II513 = ~II512,
  II514 = ~Rdy2RtHS1 & ~II263,
  II517 = ~II358 | ~II264,
  II519 = ~WantBmHS1 | ~Rdy2BmHS1,
  II1140_1 = II573 & II271,
  II521 = ~II278 | ~RtTSHS1,
  II523 = ~Prog_2 | ~II274,
  II525 = ~II280 | ~II277,
  NewTrHS1 = \[36] ,
  II526 = ~II416 & ~II370,
  II796_1 = II323 | II283,
  II529 = ~II489 | ~II399,
  II531 = ~II491 | ~II429,
  II532 = ~II327 & ~State_4,
  II534 = ~II571 & ~State_4,
  II535 = ~II534,
  II1207_1 = II579 | II519,
  II537 = ~Rdy2RtHS1 | ~II263,
  II1166_1 = II529 & II357,
  II539 = ~II274 | ~II263,
  II1166_2 = II452 & Prog_2,
  II1034_1 = II428 & II317,
  II540 = ~II449 & (~II263 & ~Rdy2RtHS1),
  II543 = ~Rdy2BmHS1 | ~II265,
  II545 = ~II362 | ~II272,
  II547 = ~II446 | ~WantRtHS1,
  II548 = ~II513 & ~State_3,
  II551 = ~II442 | ~II279,
  II552 = ~II553,
  II553 = ~II500 | ~State_1,
  II554 = ~II555,
  II555 = ~II1025_1 & ~II330,
  II556 = ~II355 | ~II1028_1,
  II559 = ~II1031_1 & ~II412,
  SeFullOHS1 = \[48] ,
  II561 = ~II1034_1 & ~II432,
  II562 = ~II439 | ~II1037_1,
  II565 = ~II1040_1 & ~II444,
  II566 = ~II567,
  II567 = ~II1044_1 & ~II388,
  II568 = ~II1047_2 | ~II1047_1,
  II570 = ~State_3 & ~II276,
  II571 = ~II570,
  II573 = ~II545 | ~II517,
  II575 = ~II284 | ~II271,
  II577 = ~II436 | (~II318 | ~State_0),
  II579 = ~II1056_1 & ~II446,
  II580 = ~II397 & ~II345,
  II582 = ~II517 & ~II331,
  II585 = ~II422 | ~II353,
  II587 = ~II317 | ~Prog_0,
  II589 = ~II482 | ~Prog_2,
  II1025_1 = II325 & Rdy2BmHS1,
  II590 = ~II539 & ~II429,
  II593 = ~II430 | ~II284,
  II595 = ~II274 | ~Rdy2BmHS1,
  II596 = ~II367 & ~II336,
  II599 = ~II354 | ~II275,
  II1176_1 = II566 & State_4,
  II1176_2 = II600 & Prog_0,
  II1044_1 = II570 & II497,
  II600 = ~II447 & ~II331,
  Mode0HS1 = \[40] ,
  II609 = ~II434 | ~II265,
  II610 = ~II284 & ~Prog_2,
  II612 = ~II274 & ~Rdy1RtHS1,
  II614 = ~II575 & ~II523,
  II624 = ~II511 & ~State_2,
  II625 = ~II624,
  II634 = ~II333 & ~II264,
  II655 = ~II1077_1 & ~II322,
  II657 = ~II1080_1 & ~II410,
  II659 = ~II1083_1 & ~II322,
  II660 = ~II469 | ~II1087_1,
  II661 = ~II660,
  II662 = ~II329 | ~II1091_1,
  II663 = ~II662,
  II665 = ~II1094_1 & ~II540,
  II667 = ~II1097_1 & ~II328,
  II669 = ~II1100_1 & ~II342,
  II1132_1 = II595 | II593,
  II1132_2 = II467 | II281,
  II671 = ~II1103_2 & ~II1103_1,
  II673 = ~II1107_1 & ~II410,
  II675 = ~II1110_1 & ~II470,
  II676 = ~II343 | ~II1113_1,
  II678 = ~II423 | ~II329,
  II680 = ~II381 | ~II445,
  II682 = ~II323 | ~II1118_1,
  II684 = ~II1121_2 | ~II1121_1,
  II1160_1 = II412 & II281,
  II686 = ~II441 | ~II1125_1,
  II689 = ~II1128_1 & ~II440,
  II690 = ~II1132_2 | ~II1132_1,
  II691 = ~II690,
  II693 = ~II1136_1 & ~II376,
  II695 = ~II328 & ~II408,
  II697 = ~II1140_1 & ~II384,
  II699 = ~II1143_2 & ~II1143_1,
  ShftIIRHS1 = \[35] ,
  Mode1HS1 = \[37] ,
  II1151_1 = II537 | II405,
  II840_1 = II284 & II283,
  II840_2 = Prog_0 & Prog_1,
  II700 = ~II351 | ~II403,
  II702 = ~II481 | ~II1148_1,
  II704 = ~II329 | ~II1151_1,
  II706 = ~II403 | ~II1154_1,
  II708 = ~II351 | ~II1157_1,
  II711 = ~II1160_1 & ~II388,
  II713 = ~II1163_1 & ~II470,
  II715 = ~II1166_2 & ~II1166_1,
  II717 = ~II1170_1 & ~II322,
  II719 = ~II1173_1 & ~II500,
  II721 = ~II1176_2 & ~II1176_1,
  II963_1 = II345 & II335,
  II723 = ~II1180_2 & ~II1180_1,
  II725 = ~II1184_2 & ~II1184_1,
  II729 = ~II1188_2 & ~II1188_1,
  II731 = ~II474 & ~II540,
  II733 = ~II1193_1 & ~II342,
  II735 = ~II1196_1 & ~II552,
  II737 = ~II1199_2 & ~II1199_1,
  II738 = ~II1203_2 | ~II1203_1,
  II1170_1 = II414 & II393,
  II740 = ~II477 | ~II1207_1,
  II742 = ~II551 | ~II1210_1,
  II744 = ~II553 | ~II1213_1,
  II746 = ~II1216_2 | ~II1216_1,
  II750 = ~II663 | ~II665,
  II1196_1 = II418 & II345,
  II767 = ~II702 & ~II704,
  II768 = ~II717 | ~II719,
  II769 = ~II768,
  Mode2HS1 = \[33] ,
  II770 = ~II713 | ~II715,
  II771 = ~II770,
  II789_1 = II580 & II278,
  II777 = ~II738 & ~II740,
  II778 = ~II735 | ~II737,
  II779 = ~II778,
  II850_1 = II612 & II610,
  II850_2 = II614 & WantRtHS1,
  II1083_1 = II506 & II458,
  II1180_1 = II322 & II267,
  II1180_2 = II554 & II348,
  LoadIIHHS1 = \[50] ,
  ActBmHS1 = \[44] ,
  II1056_1 = II358 & II280,
  ActRtHS1 = \[39] ,
  II814_1 = II355 | FullOHS1,
  II1203_1 = II491 | II463,
  II1203_2 = II577 | II543,
  II1040_1 = II322 & OutputHS1,
  II861_1 = II455 | II263,
  II861_2 = II457 | II265,
  II1107_1 = II382 & II284,
  II1094_1 = II582 & WantRtHS1,
  II1031_1 = II398 & II317,
  \[29]  = 0,
  TxHIInHS1 = \[41] ,
  II1213_1 = II547 | II498,
  \[30]  = 0,
  \[31]  = 0,
  II966_1 = II357 & II335,
  \[32]  = 0,
  II834_1 = II523 | FullIIHS1,
  \[33]  = 0,
  \[34]  = 0,
  \[35]  = 0,
  \[36]  = 0,
  \[37]  = 0,
  \[38]  = 0,
  \[39]  = 0,
  II881_1 = Prog_2 | IInDoneHS1,
  II881_2 = II326 | II282,
  \[40]  = 0,
  II1118_1 = II479 | State_1,
  \[41]  = 0,
  \[42]  = 0,
  \[43]  = 0,
  \[44]  = 0,
  TgWhBufHS1 = \[30] ,
  \[45]  = 0,
  \[46]  = 0,
  \[47]  = 0,
  \[48]  = 0,
  \[49]  = 0,
  II1128_1 = II568 & II378,
  II873_1 = II264 & II263,
  \[50]  = 0,
  II1080_1 = II382 & Prog_0,
  \[51]  = 0,
  SeOutAvHS1 = \[31] ,
  \[52]  = II2,
  \[53]  = II3,
  \[54]  = II4,
  \[55]  = II5,
  II892_1 = II495 | II279,
  II892_2 = II625 | II269,
  DumpIIHS1 = \[47] ,
  \[56]  = II6,
  \[57]  = II7,
  \[58]  = II8,
  \[59]  = II9,
  LdProgHS1 = \[32] ,
  II1157_1 = II599 | II274,
  II1216_1 = II537 | II449,
  II1216_2 = II489 | II465,
  \[60]  = II10,
  \[61]  = II11,
  II1148_1 = II565 | II267,
  \[62]  = II12,
  \[63]  = II13,
  \[64]  = II14,
  II1103_1 = II418 & State_5,
  \[65]  = II15,
  II1103_2 = II322 & Prog_0,
  \[66]  = II16,
  \[67]  = II17,
  \[68]  = II18,
  \[69]  = II19,
  II1091_1 = II587 | II585,
  ReRtTSHS1 = \[34] ,
  NewLineHS1 = \[43] ,
  \[70]  = II20,
  II1113_1 = II415 | II282,
  \[71]  = II21,
  \[72]  = II22,
  ShftORHS1 = \[38] ,
  \[73]  = II23,
  II1210_1 = II421 | II339,
  \[74]  = II24,
  \[75]  = II25,
  \[76]  = II26;
always begin
  \[8373]  = \[78] ;
  \[8374]  = \[77] ;
  \[8375]  = \[74] ;
  \[8376]  = \[79] ;
  \[8377]  = \[66] ;
  \[8378]  = \[63] ;
  \[8379]  = \[69] ;
  \[8380]  = \[62] ;
  \[8381]  = \[65] ;
  \[8382]  = \[68] ;
  \[8383]  = \[58] ;
  \[8384]  = \[64] ;
  \[8385]  = \[71] ;
  \[8386]  = \[70] ;
  \[8387]  = \[67] ;
  \[8388]  = \[59] ;
  \[8389]  = \[61] ;
  \[8390]  = \[72] ;
  \[8391]  = \[80] ;
  \[8392]  = \[75] ;
  \[8393]  = \[60] ;
  \[8394]  = \[73] ;
  \[8395]  = \[76] ;
  State_0 = \[57] ;
  State_1 = \[56] ;
  State_2 = \[55] ;
  State_3 = \[54] ;
  State_4 = \[53] ;
  State_5 = \[52] ;
end
initial begin
  \[8373]  = 0;
  \[8374]  = 0;
  \[8375]  = 0;
  \[8376]  = 0;
  \[8377]  = 0;
  \[8378]  = 0;
  \[8379]  = 0;
  \[8380]  = 0;
  \[8381]  = 0;
  \[8382]  = 0;
  \[8383]  = 0;
  \[8384]  = 0;
  \[8385]  = 0;
  \[8386]  = 0;
  \[8387]  = 0;
  \[8388]  = 0;
  \[8389]  = 0;
  \[8390]  = 0;
  \[8391]  = 0;
  \[8392]  = 0;
  \[8393]  = 0;
  \[8394]  = 0;
  \[8395]  = 0;
  State_0 = 0;
  State_1 = 0;
  State_2 = 0;
  State_3 = 0;
  State_4 = 0;
  State_5 = 0;
end
endmodule

