// IWLS benchmark module "clmB" printed on Wed May 29 22:05:43 2002
module clmb(\IN-i91 , \IN-i191 , \IN-i291 , \IN-i391 , \IN-i90 , \IN-i190 , \IN-i290 , \IN-i390 , \IN-i89 , \IN-i189 , \IN-i289 , \IN-i389 , \IN-i88 , \IN-i188 , \IN-i288 , \IN-i388 , \IN-i87 , \IN-i187 , \IN-i287 , \IN-i387 , \IN-i86 , \IN-i186 , \IN-i286 , \IN-i386 , \IN-i85 , \IN-i185 , \IN-i285 , \IN-i385 , \IN-i84 , \IN-i184 , \IN-i284 , \IN-i384 , \IN-i83 , \IN-i183 , \IN-i283 , \IN-i383 , \IN-i82 , \IN-i182 , \IN-i282 , \IN-i382 , \IN-i81 , \IN-i181 , \IN-i281 , \IN-i381 , \IN-i80 , \IN-i180 , \IN-i280 , \IN-i380 , \IN-i79 , \IN-i179 , \IN-i279 , \IN-i379 , \IN-i78 , \IN-i178 , \IN-i278 , \IN-i378 , \IN-i77 , \IN-i177 , \IN-i277 , \IN-i377 , \IN-i76 , \IN-i176 , \IN-i276 , \IN-i376 , \IN-i75 , \IN-i175 , \IN-i275 , \IN-i375 , \IN-i74 , \IN-i174 , \IN-i274 , \IN-i374 , \IN-i73 , \IN-i173 , \IN-i273 , \IN-i373 , \IN-i72 , \IN-i172 , \IN-i272 , \IN-i372 , \IN-i71 , \IN-i171 , \IN-i271 , \IN-i371 , \IN-i70 , \IN-i170 , \IN-i270 , \IN-i370 , \IN-i69 , \IN-i169 , \IN-i269 , \IN-i369 , \IN-i68 , \IN-i168 , \IN-i268 , \IN-i368 , \IN-i67 , \IN-i167 , \IN-i267 , \IN-i367 , \IN-i66 , \IN-i166 , \IN-i266 , \IN-i366 , \IN-i65 , \IN-i165 , \IN-i265 , \IN-i365 , \IN-i64 , \IN-i164 , \IN-i264 , \IN-i364 , \IN-i63 , \IN-i163 , \IN-i263 , \IN-i363 , \IN-i62 , \IN-i162 , \IN-i262 , \IN-i362 , \IN-i61 , \IN-i161 , \IN-i261 , \IN-i361 , \IN-i60 , \IN-i160 , \IN-i260 , \IN-i360 , \IN-i59 , \IN-i159 , \IN-i259 , \IN-i359 , \IN-i58 , \IN-i158 , \IN-i258 , \IN-i358 , \IN-i57 , \IN-i157 , \IN-i257 , \IN-i357 , \IN-i56 , \IN-i156 , \IN-i256 , \IN-i356 , \IN-i55 , \IN-i155 , \IN-i255 , \IN-i355 , \IN-i54 , \IN-i154 , \IN-i254 , \IN-i354 , \IN-i53 , \IN-i153 , \IN-i253 , \IN-i353 , \IN-i52 , \IN-i152 , \IN-i252 , \IN-i352 , \IN-i51 , \IN-i151 , \IN-i251 , \IN-i351 , \IN-i50 , \IN-i150 , \IN-i250 , \IN-i350 , \IN-i49 , \IN-i149 , \IN-i249 , \IN-i349 , \IN-i148 , \IN-i248 , \IN-i348 , \IN-i147 , \IN-i247 , \IN-i347 , \IN-i146 , \IN-i246 , \IN-i346 , \IN-i145 , \IN-i245 , \IN-i345 , \IN-i144 , \IN-i244 , \IN-i344 , \IN-i143 , \IN-i243 , \IN-i343 , \IN-i142 , \IN-i242 , \IN-i342 , \IN-i141 , \IN-i241 , \IN-i341 , \IN-i140 , \IN-i240 , \IN-i340 , \IN-i139 , \IN-i239 , \IN-i339 , \IN-i138 , \IN-i238 , \IN-i338 , \IN-i137 , \IN-i237 , \IN-i337 , \IN-i136 , \IN-i236 , \IN-i336 , \IN-i135 , \IN-i235 , \IN-i335 , \IN-i134 , \IN-i234 , \IN-i334 , \IN-i133 , \IN-i233 , \IN-i333 , \IN-i132 , \IN-i232 , \IN-i332 , \IN-i131 , \IN-i231 , \IN-i331 , \IN-i130 , \IN-i230 , \IN-i330 , \IN-i129 , \IN-i229 , \IN-i329 , \IN-i28 , \IN-i128 , \IN-i228 , \IN-i328 , i27, \IN-i127 , \IN-i227 , \IN-i327 , i26, \IN-i126 , \IN-i226 , \IN-i326 , i25, \IN-i125 , \IN-i225 , \IN-i325 , i24, \IN-i124 , \IN-i224 , \IN-i324 , i23, \IN-i123 , \IN-i223 , \IN-i323 , i22, \IN-i122 , \IN-i222 , \IN-i322 , i21, \IN-i121 , \IN-i221 , \IN-i321 , i20, \IN-i120 , \IN-i220 , \IN-i320 , i19, \IN-i119 , \IN-i219 , \IN-i319 , i18, \IN-i118 , \IN-i218 , \IN-i318 , i17, \IN-i117 , \IN-i217 , \IN-i317 , i16, \IN-i116 , \IN-i216 , \IN-i316 , \IN-i416 , i15, \IN-i115 , \IN-i215 , \IN-i315 , \IN-i415 , \IN-i114 , \IN-i214 , \IN-i314 , \IN-i414 , \IN-i113 , \IN-i213 , \IN-i313 , \IN-i413 , \IN-i112 , \IN-i212 , \IN-i312 , \IN-i412 , \IN-i111 , \IN-i211 , \IN-i311 , \IN-i411 , \IN-i110 , \IN-i210 , \IN-i310 , \IN-i410 , \IN-i109 , \IN-i209 , \IN-i309 , \IN-i409 , \IN-i108 , \IN-i208 , \IN-i308 , \IN-i408 , \IN-i107 , \IN-i207 , \IN-i307 , \IN-i407 , \IN-i106 , \IN-i206 , \IN-i306 , \IN-i406 , \IN-i105 , \IN-i205 , \IN-i305 , \IN-i405 , \IN-i104 , \IN-i204 , \IN-i304 , \IN-i404 , \IN-i103 , \IN-i203 , \IN-i303 , \IN-i403 , \IN-i102 , \IN-i202 , \IN-i302 , \IN-i402 , \IN-i101 , \IN-i201 , \IN-i301 , \IN-i401 , \IN-i100 , \IN-i200 , \IN-i300 , \IN-i400 , \IN-i99 , \IN-i199 , \IN-i299 , \IN-i399 , \IN-i98 , \IN-i198 , \IN-i298 , \IN-i398 , \IN-i97 , \IN-i197 , \IN-i297 , \IN-i397 , \IN-i96 , \IN-i196 , \IN-i296 , \IN-i396 , \IN-i95 , \IN-i195 , \IN-i295 , \IN-i395 , \IN-i94 , \IN-i194 , \IN-i294 , \IN-i394 , \IN-i93 , \IN-i193 , \IN-i293 , \IN-i393 , \IN-i92 , \IN-i192 , \IN-i292 , \IN-i392 , i91, i191, i291, i391, i90, i190, i290, i390, i89, i189, i289, i389, i88, i188, i288, i388, i87, i187, i287, i387, i86, i186, i286, i386, i85, i185, i285, i385, i84, i184, i284, i384, i83, i183, i283, i383, i82, i182, i282, i382, i81, i181, i281, i381, i80, i180, i280, i380, i79, i179, i279, i379, i78, i178, i278, i378, i77, i177, i277, i377, i76, i176, i276, i376, i75, i175, i275, i375, i74, i174, i274, i374, i73, i173, i273, i373, i72, i172, i272, i372, i71, i171, i271, i371, i70, i170, i270, i370, i69, i169, i269, i369, i68, i168, i268, i368, i67, i167, i267, i367, i66, i166, i266, i366, i65, i165, i265, i365, i64, i164, i264, i364, i63, i163, i263, i363, i62, i162, i262, i362, i61, i161, i261, i361, i60, i160, i260, i360, i59, i159, i259, i359, i58, i158, i258, i358, i57, i157, i257, i357, i56, i156, i256, i356, i55, i155, i255, i355, i54, i154, i254, i354, i53, i153, i253, i353, i52, i152, i252, i352, i51, i151, i251, i351, i50, i150, i250, i350, i49, i149, i249, i349, i148, i248, i348, i147, i247, i347, i146, i246, i346, i145, i245, i345, i144, i244, i344, i143, i243, i343, i142, i242, i342, i141, i241, i341, i140, i240, i340, i139, i239, i339, i138, i238, i338, i137, i237, i337, i136, i236, i336, i135, i235, i335, i134, i234, i334, i133, i233, i333, i132, i232, i332, i131, i231, i331, i130, i230, i330, i129, i229, i329, i28, i128, i228, i328, i127, i227, i327, i126, i226, i326, i125, i225, i325, i124, i224, i324, i123, i223, i323, i122, i222, i322, i121, i221, i321, i120, i220, i320, i119, i219, i319, i118, i218, i318, i117, i217, i317, i116, i216, i316, i416, i115, i215, i315, i415, i114, i214, i314, i414, i113, i213, i313, i413, i112, i212, i312, i412, i111, i211, i311, i411, i110, i210, i310, i410, i109, i209, i309, i409, i108, i208, i308, i408, i107, i207, i307, i407, i106, i206, i306, i406, i105, i205, i305, i405, i104, i204, i304, i404, i103, i203, i303, i403, i102, i202, i302, i402, i101, i201, i301, i401, i100, i200, i300, i400, i99, i199, i299, i399, i98, i198, i298, i398, i97, i197, i297, i397, i96, i196, i296, i396, i95, i195, i295, i395, i94, i194, i294, i394, i93, i193, i293, i393, i92, i192, i292, i392);
input
  \IN-i28 ,
  \IN-i49 ,
  \IN-i50 ,
  \IN-i51 ,
  \IN-i52 ,
  \IN-i53 ,
  \IN-i54 ,
  \IN-i55 ,
  \IN-i56 ,
  \IN-i57 ,
  \IN-i58 ,
  \IN-i59 ,
  \IN-i60 ,
  \IN-i61 ,
  \IN-i62 ,
  \IN-i63 ,
  \IN-i64 ,
  \IN-i65 ,
  \IN-i66 ,
  \IN-i67 ,
  \IN-i68 ,
  \IN-i69 ,
  \IN-i70 ,
  \IN-i71 ,
  \IN-i72 ,
  \IN-i73 ,
  \IN-i74 ,
  \IN-i75 ,
  \IN-i76 ,
  \IN-i77 ,
  \IN-i78 ,
  \IN-i79 ,
  \IN-i80 ,
  \IN-i81 ,
  \IN-i82 ,
  \IN-i83 ,
  \IN-i84 ,
  \IN-i85 ,
  \IN-i86 ,
  \IN-i87 ,
  \IN-i88 ,
  \IN-i89 ,
  \IN-i90 ,
  \IN-i91 ,
  \IN-i92 ,
  \IN-i93 ,
  \IN-i94 ,
  \IN-i95 ,
  \IN-i96 ,
  \IN-i97 ,
  \IN-i98 ,
  \IN-i99 ,
  i15,
  i16,
  i17,
  i18,
  i19,
  i20,
  i21,
  i22,
  i23,
  i24,
  i25,
  i26,
  i27,
  \IN-i110 ,
  \IN-i111 ,
  \IN-i112 ,
  \IN-i113 ,
  \IN-i114 ,
  \IN-i115 ,
  \IN-i116 ,
  \IN-i117 ,
  \IN-i118 ,
  \IN-i119 ,
  \IN-i120 ,
  \IN-i121 ,
  \IN-i122 ,
  \IN-i123 ,
  \IN-i124 ,
  \IN-i125 ,
  \IN-i126 ,
  \IN-i127 ,
  \IN-i128 ,
  \IN-i129 ,
  \IN-i130 ,
  \IN-i131 ,
  \IN-i132 ,
  \IN-i133 ,
  \IN-i134 ,
  \IN-i135 ,
  \IN-i136 ,
  \IN-i137 ,
  \IN-i138 ,
  \IN-i139 ,
  \IN-i140 ,
  \IN-i141 ,
  \IN-i142 ,
  \IN-i143 ,
  \IN-i144 ,
  \IN-i145 ,
  \IN-i146 ,
  \IN-i147 ,
  \IN-i148 ,
  \IN-i149 ,
  \IN-i100 ,
  \IN-i101 ,
  \IN-i102 ,
  \IN-i103 ,
  \IN-i104 ,
  \IN-i105 ,
  \IN-i106 ,
  \IN-i107 ,
  \IN-i108 ,
  \IN-i109 ,
  \IN-i190 ,
  \IN-i191 ,
  \IN-i192 ,
  \IN-i193 ,
  \IN-i194 ,
  \IN-i195 ,
  \IN-i196 ,
  \IN-i197 ,
  \IN-i198 ,
  \IN-i199 ,
  \IN-i150 ,
  \IN-i151 ,
  \IN-i152 ,
  \IN-i153 ,
  \IN-i154 ,
  \IN-i155 ,
  \IN-i156 ,
  \IN-i157 ,
  \IN-i158 ,
  \IN-i159 ,
  \IN-i160 ,
  \IN-i161 ,
  \IN-i162 ,
  \IN-i163 ,
  \IN-i164 ,
  \IN-i165 ,
  \IN-i166 ,
  \IN-i167 ,
  \IN-i168 ,
  \IN-i169 ,
  \IN-i170 ,
  \IN-i171 ,
  \IN-i172 ,
  \IN-i173 ,
  \IN-i174 ,
  \IN-i175 ,
  \IN-i176 ,
  \IN-i177 ,
  \IN-i178 ,
  \IN-i179 ,
  \IN-i180 ,
  \IN-i181 ,
  \IN-i182 ,
  \IN-i183 ,
  \IN-i184 ,
  \IN-i185 ,
  \IN-i186 ,
  \IN-i187 ,
  \IN-i188 ,
  \IN-i189 ,
  \IN-i210 ,
  \IN-i211 ,
  \IN-i212 ,
  \IN-i213 ,
  \IN-i214 ,
  \IN-i215 ,
  \IN-i216 ,
  \IN-i217 ,
  \IN-i218 ,
  \IN-i219 ,
  \IN-i220 ,
  \IN-i221 ,
  \IN-i222 ,
  \IN-i223 ,
  \IN-i224 ,
  \IN-i225 ,
  \IN-i226 ,
  \IN-i227 ,
  \IN-i228 ,
  \IN-i229 ,
  \IN-i230 ,
  \IN-i231 ,
  \IN-i232 ,
  \IN-i233 ,
  \IN-i234 ,
  \IN-i235 ,
  \IN-i236 ,
  \IN-i237 ,
  \IN-i238 ,
  \IN-i239 ,
  \IN-i240 ,
  \IN-i241 ,
  \IN-i242 ,
  \IN-i243 ,
  \IN-i244 ,
  \IN-i245 ,
  \IN-i246 ,
  \IN-i247 ,
  \IN-i248 ,
  \IN-i249 ,
  \IN-i200 ,
  \IN-i201 ,
  \IN-i202 ,
  \IN-i203 ,
  \IN-i204 ,
  \IN-i205 ,
  \IN-i206 ,
  \IN-i207 ,
  \IN-i208 ,
  \IN-i209 ,
  \IN-i290 ,
  \IN-i291 ,
  \IN-i292 ,
  \IN-i293 ,
  \IN-i294 ,
  \IN-i295 ,
  \IN-i296 ,
  \IN-i297 ,
  \IN-i298 ,
  \IN-i299 ,
  \IN-i250 ,
  \IN-i251 ,
  \IN-i252 ,
  \IN-i253 ,
  \IN-i254 ,
  \IN-i255 ,
  \IN-i256 ,
  \IN-i257 ,
  \IN-i258 ,
  \IN-i259 ,
  \IN-i260 ,
  \IN-i261 ,
  \IN-i262 ,
  \IN-i263 ,
  \IN-i264 ,
  \IN-i265 ,
  \IN-i266 ,
  \IN-i267 ,
  \IN-i268 ,
  \IN-i269 ,
  \IN-i270 ,
  \IN-i271 ,
  \IN-i272 ,
  \IN-i273 ,
  \IN-i274 ,
  \IN-i275 ,
  \IN-i276 ,
  \IN-i277 ,
  \IN-i278 ,
  \IN-i279 ,
  \IN-i280 ,
  \IN-i281 ,
  \IN-i282 ,
  \IN-i283 ,
  \IN-i284 ,
  \IN-i285 ,
  \IN-i286 ,
  \IN-i287 ,
  \IN-i288 ,
  \IN-i289 ,
  \IN-i310 ,
  \IN-i311 ,
  \IN-i312 ,
  \IN-i313 ,
  \IN-i314 ,
  \IN-i315 ,
  \IN-i316 ,
  \IN-i317 ,
  \IN-i318 ,
  \IN-i319 ,
  \IN-i320 ,
  \IN-i321 ,
  \IN-i322 ,
  \IN-i323 ,
  \IN-i324 ,
  \IN-i325 ,
  \IN-i326 ,
  \IN-i327 ,
  \IN-i328 ,
  \IN-i329 ,
  \IN-i330 ,
  \IN-i331 ,
  \IN-i332 ,
  \IN-i333 ,
  \IN-i334 ,
  \IN-i335 ,
  \IN-i336 ,
  \IN-i337 ,
  \IN-i338 ,
  \IN-i339 ,
  \IN-i340 ,
  \IN-i341 ,
  \IN-i342 ,
  \IN-i343 ,
  \IN-i344 ,
  \IN-i345 ,
  \IN-i346 ,
  \IN-i347 ,
  \IN-i348 ,
  \IN-i349 ,
  \IN-i300 ,
  \IN-i301 ,
  \IN-i302 ,
  \IN-i303 ,
  \IN-i304 ,
  \IN-i305 ,
  \IN-i306 ,
  \IN-i307 ,
  \IN-i308 ,
  \IN-i309 ,
  \IN-i390 ,
  \IN-i391 ,
  \IN-i392 ,
  \IN-i393 ,
  \IN-i394 ,
  \IN-i395 ,
  \IN-i396 ,
  \IN-i397 ,
  \IN-i398 ,
  \IN-i399 ,
  \IN-i350 ,
  \IN-i351 ,
  \IN-i352 ,
  \IN-i353 ,
  \IN-i354 ,
  \IN-i355 ,
  \IN-i356 ,
  \IN-i357 ,
  \IN-i358 ,
  \IN-i359 ,
  \IN-i360 ,
  \IN-i361 ,
  \IN-i362 ,
  \IN-i363 ,
  \IN-i364 ,
  \IN-i365 ,
  \IN-i366 ,
  \IN-i367 ,
  \IN-i368 ,
  \IN-i369 ,
  \IN-i370 ,
  \IN-i371 ,
  \IN-i372 ,
  \IN-i373 ,
  \IN-i374 ,
  \IN-i375 ,
  \IN-i376 ,
  \IN-i377 ,
  \IN-i378 ,
  \IN-i379 ,
  \IN-i380 ,
  \IN-i381 ,
  \IN-i382 ,
  \IN-i383 ,
  \IN-i384 ,
  \IN-i385 ,
  \IN-i386 ,
  \IN-i387 ,
  \IN-i388 ,
  \IN-i389 ,
  \IN-i410 ,
  \IN-i411 ,
  \IN-i412 ,
  \IN-i413 ,
  \IN-i414 ,
  \IN-i415 ,
  \IN-i416 ,
  \IN-i400 ,
  \IN-i401 ,
  \IN-i402 ,
  \IN-i403 ,
  \IN-i404 ,
  \IN-i405 ,
  \IN-i406 ,
  \IN-i407 ,
  \IN-i408 ,
  \IN-i409 ;
output
  i100,
  i101,
  i102,
  i103,
  i104,
  i105,
  i106,
  i107,
  i108,
  i109,
  i110,
  i111,
  i112,
  i113,
  i114,
  i115,
  i116,
  i117,
  i118,
  i119,
  i120,
  i121,
  i122,
  i123,
  i124,
  i125,
  i126,
  i127,
  i128,
  i129,
  i130,
  i131,
  i132,
  i133,
  i134,
  i135,
  i136,
  i137,
  i138,
  i139,
  i140,
  i141,
  i142,
  i143,
  i144,
  i145,
  i146,
  i147,
  i148,
  i149,
  i150,
  i151,
  i152,
  i153,
  i154,
  i155,
  i156,
  i157,
  i158,
  i159,
  i160,
  i161,
  i162,
  i163,
  i164,
  i165,
  i166,
  i167,
  i168,
  i169,
  i170,
  i171,
  i172,
  i173,
  i174,
  i175,
  i176,
  i177,
  i178,
  i179,
  i180,
  i181,
  i182,
  i183,
  i184,
  i185,
  i186,
  i187,
  i188,
  i189,
  i190,
  i191,
  i192,
  i193,
  i194,
  i195,
  i196,
  i197,
  i198,
  i199,
  i200,
  i201,
  i202,
  i203,
  i204,
  i205,
  i206,
  i207,
  i208,
  i209,
  i210,
  i211,
  i212,
  i213,
  i214,
  i215,
  i216,
  i217,
  i218,
  i219,
  i220,
  i221,
  i222,
  i223,
  i224,
  i225,
  i226,
  i227,
  i228,
  i229,
  i230,
  i231,
  i232,
  i233,
  i234,
  i235,
  i236,
  i237,
  i238,
  i239,
  i240,
  i241,
  i242,
  i243,
  i244,
  i245,
  i246,
  i247,
  i248,
  i249,
  i250,
  i251,
  i252,
  i253,
  i254,
  i255,
  i256,
  i257,
  i258,
  i259,
  i260,
  i261,
  i262,
  i263,
  i264,
  i265,
  i266,
  i267,
  i268,
  i269,
  i270,
  i271,
  i272,
  i273,
  i274,
  i275,
  i276,
  i277,
  i278,
  i279,
  i280,
  i281,
  i282,
  i283,
  i284,
  i285,
  i286,
  i287,
  i288,
  i289,
  i290,
  i291,
  i292,
  i293,
  i294,
  i295,
  i296,
  i297,
  i298,
  i299,
  i300,
  i301,
  i302,
  i303,
  i304,
  i305,
  i306,
  i307,
  i308,
  i309,
  i310,
  i311,
  i312,
  i313,
  i314,
  i315,
  i316,
  i317,
  i318,
  i319,
  i320,
  i321,
  i322,
  i323,
  i324,
  i325,
  i326,
  i327,
  i328,
  i329,
  i330,
  i331,
  i332,
  i333,
  i334,
  i335,
  i336,
  i337,
  i338,
  i339,
  i340,
  i341,
  i342,
  i343,
  i344,
  i345,
  i346,
  i347,
  i348,
  i349,
  i350,
  i351,
  i352,
  i353,
  i354,
  i355,
  i356,
  i357,
  i358,
  i359,
  i360,
  i361,
  i362,
  i363,
  i364,
  i365,
  i366,
  i367,
  i368,
  i369,
  i370,
  i371,
  i372,
  i373,
  i374,
  i375,
  i376,
  i377,
  i378,
  i379,
  i380,
  i381,
  i382,
  i383,
  i384,
  i385,
  i386,
  i387,
  i388,
  i389,
  i390,
  i391,
  i392,
  i393,
  i394,
  i395,
  i396,
  i397,
  i398,
  i399,
  i400,
  i401,
  i402,
  i403,
  i404,
  i405,
  i406,
  i407,
  i408,
  i409,
  i410,
  i411,
  i412,
  i413,
  i414,
  i415,
  i416,
  i28,
  i49,
  i50,
  i51,
  i52,
  i53,
  i54,
  i55,
  i56,
  i57,
  i58,
  i59,
  i60,
  i61,
  i62,
  i63,
  i64,
  i65,
  i66,
  i67,
  i68,
  i69,
  i70,
  i71,
  i72,
  i73,
  i74,
  i75,
  i76,
  i77,
  i78,
  i79,
  i80,
  i81,
  i82,
  i83,
  i84,
  i85,
  i86,
  i87,
  i88,
  i89,
  i90,
  i91,
  i92,
  i93,
  i94,
  i95,
  i96,
  i97,
  i98,
  i99;
reg
  i2,
  i3,
  i4,
  i5,
  i6,
  i7,
  i8,
  i9,
  i10,
  i11,
  i12,
  i13,
  i14,
  i29,
  i30,
  i31,
  i32,
  i33,
  i34,
  i35,
  i36,
  i37,
  i38,
  i39,
  i40,
  i41,
  i42,
  i43,
  i44,
  i45,
  i46,
  i47,
  i48;
wire
  v5374,
  v5375,
  v5376,
  v5377,
  v5378,
  v5379,
  v5380,
  v5381,
  v5382,
  v5383,
  v5384,
  v5385,
  v5386,
  v5387,
  v5388,
  v5389,
  v5390,
  v5391,
  v5392,
  v5393,
  v5394,
  v5395,
  v5396,
  v5397,
  v5398,
  v5399,
  v5400,
  v5401,
  v5402,
  v5403,
  v5404,
  v5405,
  v5406,
  v5407,
  v5408,
  v5409,
  v5410,
  v5411,
  v5412,
  v5413,
  v5414,
  v5415,
  v5416,
  v5417,
  v5418,
  v5419,
  v5420,
  v5421,
  v5422,
  v5423,
  v5424,
  v5425,
  v5426,
  v5427,
  v5428,
  v5429,
  v5430,
  v5431,
  v5432,
  v5433,
  v5434,
  v5435,
  v5436,
  v5437,
  v5438,
  v5439,
  v5440,
  v5441,
  v5442,
  v5443,
  v5444,
  v5445,
  v5446,
  v5447,
  v5448,
  v5449,
  v5450,
  v5451,
  v5452,
  v5453,
  v5454,
  v5455,
  v5456,
  v5457,
  v5458,
  v5459,
  v5460,
  v5461,
  v5462,
  v5463,
  v5464,
  v5465,
  v5466,
  v5467,
  v5468,
  v5469,
  v5470,
  v5471,
  v5472,
  v5473,
  v5474,
  v5475,
  v5476,
  v5477,
  v5478,
  v5479,
  v5480,
  v5481,
  v5482,
  v5483,
  v5484,
  v5485,
  v5486,
  v5487,
  v5488,
  v5489,
  v5490,
  v5491,
  v5492,
  v5493,
  v5494,
  v5495,
  v5496,
  v5497,
  v5498,
  v5499,
  v5500,
  v5501,
  v5502,
  v5503,
  v5504,
  v5505,
  v5506,
  v5507,
  v5508,
  v5509,
  v5510,
  v5511,
  v5512,
  v5513,
  v5514,
  v5515,
  v5516,
  v5517,
  v5518,
  v5519,
  v5520,
  v5521,
  v5522,
  v5523,
  v5524,
  v5525,
  v5526,
  v5527,
  v5528,
  v5529,
  v5530,
  v5531,
  v5532,
  v5533,
  v5534,
  v5535,
  v5536,
  v5537,
  v5538,
  v5539,
  v5540,
  v5541,
  v5542,
  v5543,
  v5544,
  v5545,
  v5546,
  v5547,
  v5548,
  v5549,
  v5550,
  v5551,
  v5552,
  v5553,
  v5554,
  v5555,
  v5556,
  v5557,
  v5558,
  v5559,
  v5560,
  v5561,
  v5562,
  v5563,
  v5564,
  v5565,
  v5566,
  v5567,
  v5568,
  v5569,
  v5570,
  v5571,
  v5572,
  v5573,
  v5574,
  v5575,
  v5576,
  v5577,
  v5578,
  v5579,
  v5580,
  v5581,
  v5582,
  v5583,
  v5584,
  v5585,
  v5586,
  v5587,
  v5588,
  v5589,
  v5590,
  v5591,
  v5592,
  v5593,
  v5594,
  v5595,
  v5596,
  v5597,
  v5598,
  v5599,
  v5600,
  v5601,
  v5602,
  v5603,
  v5604,
  v5605,
  v5606,
  v5607,
  v5608,
  v5609,
  v5610,
  v5611,
  v5612,
  v5613,
  v5614,
  v5615,
  v5616,
  v5617,
  v5618,
  v5619,
  v5620,
  v5621,
  v5622,
  v5623,
  v5624,
  v5625,
  v5626,
  v5627,
  v5628,
  v5629,
  v5630,
  v5631,
  v5632,
  v5633,
  v5634,
  v5635,
  v5636,
  v5637,
  v5638,
  v5639,
  v5640,
  v5641,
  v5642,
  v5643,
  v5644,
  v5645,
  v5646,
  v5647,
  v5648,
  v5649,
  v5650,
  v5651,
  v5652,
  v5653,
  v5654,
  v5655,
  v5656,
  v5657,
  v5658,
  v5659,
  v5660,
  v5661,
  v5662,
  v5663,
  v5664,
  v5665,
  v5666,
  v5667,
  v5668,
  v5669,
  v5670,
  v5671,
  v5672,
  v5673,
  v5674,
  v5675,
  v5676,
  v5677,
  v5678,
  v5679,
  v5680,
  v5681,
  v5682,
  v5683,
  v5684,
  v5685,
  v5686,
  v5687,
  v5688,
  v5689,
  v5690,
  v5691,
  v5692,
  v5693,
  v5694,
  v5695,
  v5696,
  v5697,
  v5698,
  v5699,
  v5700,
  v5701,
  v5702,
  v5703,
  v5704,
  v5705,
  v5706,
  v5707,
  v5708,
  v5709,
  v5710,
  v5711,
  v5712,
  v5713,
  v5714,
  v5715,
  v5716,
  v5717,
  v5718,
  v5719,
  v5720,
  v5721,
  v5722,
  v5723,
  v5724,
  v5725,
  v5726,
  v5727,
  v5728,
  v5729,
  v5730,
  v5731,
  v5732,
  v5733,
  v5734,
  v5735,
  v5736,
  v5737,
  v5738,
  v5739,
  v5740,
  v5741,
  v5742,
  v5743,
  v5744,
  v5745,
  v5746,
  v5747,
  v5748,
  v5749,
  v5750,
  v5751,
  v5752,
  v5753,
  v5754,
  v5755,
  v5756,
  v5757,
  v5758,
  v5759,
  v5760,
  v5761,
  v5762,
  v5763,
  v5764,
  v5765,
  v5766,
  v5767,
  v5768,
  v5769,
  v5770,
  v5771,
  v5772,
  v5773,
  v5774,
  v5775,
  v5776,
  v5777,
  v5778,
  v5779,
  v5780,
  v5781,
  v5782,
  v5783,
  v5784,
  v5785,
  v5786,
  v5787,
  v5788,
  v5789,
  v5790,
  v5791,
  v5792,
  v5793,
  v5794,
  v5795,
  v5796,
  v5797,
  v5798,
  v5799,
  v5800,
  v5801,
  v5802,
  v5803,
  v5804,
  v5805,
  v5806,
  v5807,
  v5808,
  v5809,
  v5810,
  v5811,
  v5812,
  v5813,
  v5814,
  v5815,
  v5816,
  v5817,
  v5818,
  v5819,
  v5820,
  v5821,
  v5822,
  v5823,
  v5824,
  v5825,
  v5826,
  v5827,
  v5828,
  v5829,
  v5830,
  v5831,
  v5832,
  v5833,
  v5834,
  v5835,
  v5836,
  v5837,
  v5838,
  v5839,
  v5840,
  v5841,
  v5842,
  v5843,
  v5844,
  v5845,
  v5846,
  v5847,
  v5848,
  v5849,
  v5850,
  v5851,
  v5852,
  v5853,
  v5854,
  v5855,
  v5856,
  v5857,
  v5858,
  v5859,
  v5860,
  v5861,
  v5862,
  v5863,
  v5864,
  v5865,
  v5866,
  v5867,
  v5868,
  v5869,
  v5870,
  v5871,
  v5872,
  v5873,
  v5874,
  v5875,
  v5876,
  v5877,
  v5878,
  v5879,
  v5880,
  v5881,
  v5882,
  v5883,
  v5884,
  v5885,
  v5886,
  v5887,
  v5888,
  v5889,
  v5890,
  v5891,
  v5892,
  v5893,
  v5894,
  v5895,
  v5896,
  v5897,
  v5898,
  v5899,
  v5900,
  v5901,
  v5902,
  v5903,
  v5904,
  v5905,
  v5906,
  v5907,
  v5908,
  v5909,
  v5910,
  v5911,
  v5912,
  v5913,
  v5914,
  v5915,
  v5916,
  v5917,
  v5918,
  v5919,
  v5920,
  v5921,
  \[402] ,
  v5922,
  v5923,
  v5924,
  v5925,
  v5926,
  v5927,
  v5928,
  v5929,
  v5930,
  v5931,
  \[403] ,
  v5932,
  v5933,
  v5934,
  v5935,
  v5936,
  v5937,
  v5938,
  v5939,
  v5940,
  v5941,
  \[404] ,
  v5942,
  v5943,
  v5944,
  v5945,
  v5946,
  v5947,
  v5948,
  v5949,
  v5950,
  v5951,
  \[405] ,
  v5952,
  v5953,
  v5954,
  v5955,
  v5956,
  v5957,
  v5958,
  v5959,
  v5960,
  v5961,
  \[406] ,
  v5962,
  v5963,
  v5964,
  v5965,
  v5966,
  v5967,
  v5968,
  v5969,
  v5970,
  v5971,
  \[407] ,
  v5972,
  v5973,
  v5974,
  v5975,
  v5976,
  v5977,
  v5978,
  v5979,
  v5980,
  v5981,
  \[408] ,
  v5982,
  v5983,
  v5984,
  v5985,
  v5986,
  v5987,
  v5988,
  v5989,
  v5990,
  v5991,
  \[409] ,
  v5992,
  v5993,
  v5994,
  v5995,
  v5996,
  v5997,
  v5998,
  v5999,
  \[410] ,
  \[411] ,
  \[412] ,
  \[413] ,
  \[414] ,
  \[415] ,
  \[416] ,
  \[417] ,
  \[418] ,
  \[419] ,
  \[420] ,
  v2,
  v3,
  v4,
  v5,
  v6,
  v7,
  v8,
  v9,
  \[421] ,
  \[422] ,
  \[423] ,
  \[424] ,
  \[425] ,
  \[426] ,
  \[427] ,
  \[428] ,
  \[429] ,
  \[430] ,
  \[431] ,
  \[432] ,
  \[433] ,
  \[434] ,
  v6000,
  v6001,
  v6002,
  v6003,
  v6004,
  v6005,
  v6006,
  v6007,
  v6008,
  v6009,
  v6010,
  v6011,
  v6012,
  v6013,
  v6014,
  v6015,
  v6016,
  v6017,
  v6018,
  v6019,
  v6020,
  v6021,
  v6022,
  v6023,
  v6024,
  v6025,
  v6026,
  v6027,
  v6028,
  v6029,
  v6030,
  v6031,
  v6032,
  v6033,
  v6034,
  v6035,
  v6036,
  v6037,
  v6038,
  v6039,
  v6040,
  v6041,
  v6042,
  v6043,
  v6044,
  v6045,
  v6046,
  v6047,
  v6048,
  v6049,
  v6050,
  v6051,
  v6052,
  v6053,
  v6054,
  v6055,
  v6056,
  v6057,
  v6058,
  v6059,
  v6060,
  v6061,
  v6062,
  v6063,
  v6064,
  v6065,
  v6066,
  v6067,
  v6068,
  v6069,
  v6070,
  v6071,
  v6072,
  v6073,
  v6074,
  v6075,
  v6076,
  v6077,
  v6078,
  v6079,
  v6080,
  v6081,
  v6082,
  v6083,
  v6084,
  v6085,
  v6086,
  v6087,
  v6088,
  v6089,
  v6090,
  v6091,
  v6092,
  v6093,
  v6094,
  v6095,
  v6096,
  v6097,
  v6098,
  v6099,
  v6100,
  v6101,
  v6102,
  v6103,
  v6104,
  v6105,
  v6106,
  v6107,
  v6108,
  v6109,
  v6110,
  v6111,
  v6112,
  v6113,
  v6114,
  v6115,
  v6116,
  v6117,
  v6118,
  v6119,
  v6120,
  v6121,
  v6122,
  v6123,
  v6124,
  v6125,
  v6126,
  v6127,
  v6128,
  v6129,
  v6130,
  v6131,
  v6132,
  v6133,
  v6134,
  v6135,
  v6136,
  v6137,
  v6138,
  v6139,
  v6140,
  v6141,
  v6142,
  v6143,
  v6144,
  v6145,
  v6146,
  v6147,
  v6148,
  v6149,
  v6150,
  v6151,
  v6152,
  v6153,
  v6154,
  v6155,
  v6156,
  v6157,
  v6158,
  v6159,
  v6160,
  v6161,
  v6162,
  v6163,
  v6164,
  v6165,
  v6166,
  v6167,
  v6168,
  v6169,
  v6170,
  v6171,
  v6172,
  v6173,
  v6174,
  v6175,
  v6176,
  v6177,
  v6178,
  v6179,
  v6180,
  v6181,
  v6182,
  v6183,
  v6184,
  v6185,
  v6186,
  v6187,
  v6188,
  v6189,
  v6190,
  v6191,
  v6192,
  v6193,
  v6194,
  v6195,
  v6196,
  v6197,
  v6198,
  v6199,
  v6200,
  v6201,
  v6202,
  v6203,
  v6204,
  v6205,
  v6206,
  v6207,
  v6208,
  v6209,
  v6210,
  v6211,
  v6212,
  v6213,
  v6214,
  v6215,
  v6216,
  v6217,
  v6218,
  v6219,
  v6220,
  v6221,
  v6222,
  v6223,
  v6224,
  v6225,
  v6226,
  v6227,
  v6228,
  v6229,
  v6230,
  v6231,
  v6232,
  v6233,
  v6234,
  v6235,
  v6236,
  v6237,
  v6238,
  v6239,
  v6240,
  v6241,
  v6242,
  v6243,
  v6244,
  v6245,
  v6246,
  v6247,
  v6248,
  v6249,
  v6250,
  v6251,
  v6252,
  v6253,
  v6254,
  v6255,
  v6256,
  v6257,
  v6258,
  v6259,
  v6260,
  v6261,
  v6262,
  v6263,
  v6264,
  v6265,
  v6266,
  v6267,
  v6268,
  v6269,
  v6270,
  v6271,
  v6272,
  v6273,
  v6274,
  v6275,
  v6276,
  v6277,
  v6278,
  v6279,
  v6280,
  v6281,
  v6282,
  v6283,
  v6284,
  v6285,
  v6286,
  v6287,
  v6288,
  v6289,
  v6290,
  v6291,
  v6292,
  v6293,
  v6294,
  v6295,
  v6296,
  v6297,
  v6298,
  v6299,
  v6300,
  v6301,
  v6302,
  v6303,
  v6304,
  v6305,
  v6306,
  v6307,
  v6308,
  v6309,
  v6310,
  v6311,
  v6312,
  v6313,
  v6314,
  v6315,
  v6316,
  v6317,
  v6318,
  v6319,
  v6320,
  v6321,
  v6322,
  v6323,
  v6324,
  v6325,
  v6326,
  v6327,
  v6328,
  v6329,
  v6330,
  v6331,
  v6332,
  v6333,
  v6334,
  v6335,
  v6336,
  v6337,
  v6338,
  v6339,
  v6340,
  v6341,
  v6342,
  v6343,
  v6344,
  v6345,
  v6346,
  v6347,
  v6348,
  v6349,
  v6350,
  v6351,
  v6352,
  v6353,
  v6354,
  v6355,
  v6356,
  v6357,
  v6358,
  v6359,
  v6360,
  v6361,
  v6362,
  v6363,
  v6364,
  v6365,
  v6366,
  v6367,
  v6368,
  v6369,
  v6370,
  v6371,
  v6372,
  v6373,
  v6374,
  v6375,
  v6376,
  v6377,
  v6378,
  v6379,
  v6380,
  v6381,
  v6382,
  v6383,
  v6384,
  v6385,
  v6386,
  v6387,
  v6388,
  v6389,
  v6390,
  v6391,
  v6392,
  v6393,
  v6394,
  v6395,
  v6396,
  v6397,
  v6398,
  v6399,
  v6400,
  v6401,
  v6402,
  v6403,
  v6404,
  v6405,
  v6406,
  v6407,
  v6408,
  v6409,
  v6410,
  v6411,
  v6412,
  v6413,
  v6414,
  v6415,
  v6416,
  v6417,
  v6418,
  v6419,
  v6420,
  v6421,
  v6422,
  v6423,
  v6424,
  v6425,
  v6426,
  v6427,
  v6428,
  v6429,
  v6430,
  v6431,
  v6432,
  v6433,
  v6434,
  v6435,
  v6436,
  v6437,
  v6438,
  v6439,
  v6440,
  v6441,
  v6442,
  v6443,
  v6444,
  v6445,
  v6446,
  v6447,
  v6448,
  v6449,
  v6450,
  v6451,
  v6452,
  v6453,
  v6454,
  v6455,
  v6456,
  v6457,
  v6458,
  v6459,
  v6460,
  v6461,
  v6462,
  v6463,
  v6464,
  v6465,
  v6466,
  v6467,
  v6468,
  v6469,
  v6470,
  v6471,
  v6472,
  v6473,
  v6474,
  v6475,
  v6476,
  v6477,
  v6478,
  v6479,
  v6480,
  v6481,
  v6482,
  v6483,
  v6484,
  v6485,
  v6486,
  v6487,
  v6488,
  v6489,
  v6490,
  v6491,
  v6492,
  v6493,
  v6494,
  v6495,
  v6496,
  v6497,
  v6498,
  v6499,
  v6500,
  v6501,
  v6502,
  v6503,
  v6504,
  v6505,
  v6506,
  v6507,
  v6508,
  v6509,
  v6510,
  v6511,
  v6512,
  v6513,
  v6514,
  v6515,
  v6516,
  v6517,
  v6518,
  v6519,
  v6520,
  v6521,
  v6522,
  v6523,
  v6524,
  v6525,
  v6526,
  v6527,
  v6528,
  v6529,
  v6530,
  v6531,
  v6532,
  v6533,
  v6534,
  v6535,
  v6536,
  v6537,
  v6538,
  v6539,
  v6540,
  v6541,
  v6542,
  v6543,
  v6544,
  v6545,
  v6546,
  v6547,
  v6548,
  v6549,
  v6550,
  v6551,
  v6552,
  v6553,
  v6554,
  v6555,
  v6556,
  v6557,
  v6558,
  v6559,
  v6560,
  v6561,
  v6562,
  v6563,
  v6564,
  v6565,
  v6566,
  v6567,
  v6568,
  v6569,
  v6570,
  v6571,
  v6572,
  v6573,
  v6574,
  v6575,
  v6576,
  v6577,
  v6578,
  v6579,
  v6580,
  v6581,
  v6582,
  v6583,
  v6584,
  v6585,
  v6586,
  v6587,
  v6588,
  v6589,
  v6590,
  v6591,
  v6592,
  v6593,
  v6594,
  v6595,
  v6596,
  v6597,
  v6598,
  v6599,
  v6600,
  v6601,
  v6602,
  v6603,
  v6604,
  v6605,
  v6606,
  v6607,
  v6608,
  v6609,
  v6610,
  v6611,
  v6612,
  v6613,
  v6614,
  v6615,
  v6616,
  v6617,
  v6618,
  v6619,
  v6620,
  v6621,
  v6622,
  v6623,
  v6624,
  v6625,
  v6626,
  v6627,
  v6628,
  v6629,
  v6630,
  v6631,
  v6632,
  v6633,
  v6634,
  v6635,
  v6636,
  v6637,
  v6638,
  v6639,
  v6640,
  v6641,
  v6642,
  v6643,
  v6644,
  v6645,
  v6646,
  v6647,
  v6648,
  v6649,
  v6650,
  v6651,
  v6652,
  v6653,
  v6654,
  v6655,
  v6656,
  v6657,
  v6658,
  v6659,
  v6660,
  v6661,
  v6662,
  v6663,
  v6664,
  v6665,
  v6666,
  v6667,
  v6668,
  v6669,
  v6670,
  v6671,
  v6672,
  v6673,
  v6674,
  v6675,
  v6676,
  v6677,
  v6678,
  v6679,
  v6680,
  v6681,
  v6682,
  v6683,
  v6684,
  v6685,
  v6686,
  v6687,
  v6688,
  v6689,
  v6690,
  v6691,
  v6692,
  v6693,
  v6694,
  v6695,
  v6696,
  v6697,
  v6698,
  v6699,
  v6700,
  v6701,
  v6702,
  v6703,
  v6704,
  v6705,
  v6706,
  v6707,
  v6708,
  v6709,
  v6710,
  v6711,
  v6712,
  v6713,
  v6714,
  v6715,
  v6716,
  v6717,
  v6718,
  v6719,
  v6720,
  v6721,
  v6722,
  v6723,
  v6724,
  v6725,
  v6726,
  v6727,
  v6728,
  v6729,
  v6730,
  v6731,
  v6732,
  v6733,
  v6734,
  v6735,
  v6736,
  v6737,
  v6738,
  v6739,
  v6740,
  v6741,
  v6742,
  v6743,
  v6744,
  v6745,
  v6746,
  v6747,
  v6748,
  v6749,
  v6750,
  v6751,
  v6752,
  v6753,
  v6754,
  v6755,
  v6756,
  v6757,
  v6758,
  v6759,
  v6760,
  v6761,
  v6762,
  v6763,
  v6764,
  v6765,
  v6766,
  v6767,
  v6768,
  v6769,
  v6770,
  v6771,
  v6772,
  v6773,
  v6774,
  v6775,
  v6776,
  v6777,
  v6778,
  v6779,
  v6780,
  v6781,
  v6782,
  v6783,
  v6784,
  v6785,
  v6786,
  v6787,
  v6788,
  v6789,
  v6790,
  v6791,
  v6792,
  v6793,
  v6794,
  v6795,
  v6796,
  v6797,
  v6798,
  v6799,
  v6800,
  v6801,
  v6802,
  v6803,
  v6804,
  v6805,
  v6806,
  v6807,
  v6808,
  v6809,
  v6810,
  v6811,
  v6812,
  v6813,
  v6814,
  v6815,
  v6816,
  v6817,
  v6818,
  v6819,
  v6820,
  v6821,
  v6822,
  v6823,
  v6824,
  v6825,
  v6826,
  v6827,
  v6828,
  v6829,
  v6830,
  v6831,
  v6832,
  v6833,
  v6834,
  v6835,
  v6836,
  v6837,
  v6838,
  v6839,
  v6840,
  v6841,
  v6842,
  v6843,
  v6844,
  v6845,
  v6846,
  v6847,
  v6848,
  v6849,
  v6850,
  v6851,
  v6852,
  v6853,
  v6854,
  v6855,
  v6856,
  v6857,
  v6858,
  v6859,
  v6860,
  v6861,
  v6862,
  v6863,
  v6864,
  v6865,
  v6866,
  v6867,
  v6868,
  v6869,
  v6870,
  v6871,
  v6872,
  v6873,
  v6874,
  v6875,
  v6876,
  v6877,
  v6878,
  v6879,
  v6880,
  v6881,
  v6882,
  v6883,
  v6884,
  v6885,
  v6886,
  v6887,
  v6888,
  v6889,
  v6890,
  v6891,
  v6892,
  v6893,
  v6894,
  v6895,
  v6896,
  v6897,
  v6898,
  v6899,
  v6900,
  v6901,
  v6902,
  v6903,
  v6904,
  v6905,
  v6906,
  v6907,
  v6908,
  v6909,
  v6910,
  v6911,
  v6912,
  v6913,
  v6914,
  v6915,
  v6916,
  v6917,
  v6918,
  v6919,
  v6920,
  v6921,
  v6922,
  v6923,
  v6924,
  v6925,
  v6926,
  v6927,
  v6928,
  v6929,
  v6930,
  v6931,
  v6932,
  v6933,
  v6934,
  v6935,
  v6936,
  v6937,
  v6938,
  v6939,
  v6940,
  v6941,
  v6942,
  v6943,
  v6944,
  v6945,
  v6946,
  v6947,
  v6948,
  v6949,
  v6950,
  v6951,
  v6952,
  v6953,
  v6954,
  v6955,
  v6956,
  v6957,
  v6958,
  v6959,
  v6960,
  v6961,
  v6962,
  v6963,
  v6964,
  v6965,
  v6966,
  v6967,
  v6968,
  v6969,
  v6970,
  v6971,
  v6972,
  v6973,
  v6974,
  v6975,
  v6976,
  v6977,
  v6978,
  v6979,
  v6980,
  v6981,
  v6982,
  v6983,
  v6984,
  v6985,
  v6986,
  v6987,
  v6988,
  v6989,
  v6990,
  v6991,
  v6992,
  v6993,
  v6994,
  v6995,
  v6996,
  v6997,
  v6998,
  v6999,
  v7000,
  v7001,
  v7002,
  v7003,
  v7004,
  v7005,
  v7006,
  v7007,
  v7008,
  v7009,
  v7010,
  v7011,
  v7012,
  v7013,
  v7014,
  v7015,
  v7016,
  v7017,
  v7018,
  v7019,
  v7020,
  v7021,
  v7022,
  v7023,
  v7024,
  v7025,
  v7026,
  v7027,
  v7028,
  v7029,
  v7030,
  v7031,
  v7032,
  v7033,
  v7034,
  v7035,
  v7036,
  v7037,
  v7038,
  v7039,
  v7040,
  v7041,
  v7042,
  v7043,
  v7044,
  v7045,
  v7046,
  v7047,
  v7048,
  v7049,
  v7050,
  v7051,
  v7052,
  v7053,
  v7054,
  v7055,
  v7056,
  v7057,
  v7058,
  v7059,
  v7060,
  v7061,
  v7062,
  v7063,
  v7064,
  v7065,
  v7066,
  v7067,
  v7068,
  v7069,
  v7070,
  v7071,
  v7072,
  v7073,
  v7074,
  v7075,
  v7076,
  v7077,
  v7078,
  v7079,
  v7080,
  v7081,
  v7082,
  v7083,
  v7084,
  v7085,
  v7086,
  v7087,
  v7088,
  v7089,
  v7090,
  v7091,
  v7092,
  v7093,
  v7094,
  v7095,
  v7096,
  v7097,
  v7098,
  v7099,
  v7100,
  v7101,
  v7102,
  v7103,
  v7104,
  v7105,
  v7106,
  v7107,
  v7108,
  v7109,
  v7110,
  v7111,
  v7112,
  v7113,
  v7114,
  v7115,
  v7116,
  v7117,
  v7118,
  v7119,
  v7120,
  v7121,
  v7122,
  v7123,
  v7124,
  v7125,
  v7126,
  v7127,
  v7128,
  v7129,
  v7130,
  v7131,
  v7132,
  v7133,
  v7134,
  v7135,
  v7136,
  v7137,
  v7138,
  v7139,
  v7140,
  v7141,
  v7142,
  v7143,
  v7144,
  v7145,
  v7146,
  v7147,
  v7148,
  v7149,
  v7150,
  v7151,
  v7152,
  v7153,
  v7154,
  v7155,
  v7156,
  v7157,
  v7158,
  v7159,
  v7160,
  v7161,
  v7162,
  v7163,
  v7164,
  v7165,
  v7166,
  v7167,
  v7168,
  v7169,
  v7170,
  v7171,
  v7172,
  v7173,
  v7174,
  v7175,
  v7176,
  v7177,
  v7178,
  v7179,
  v7180,
  v7181,
  v7182,
  v7183,
  v7184,
  v7185,
  v7186,
  v7187,
  v7188,
  v7189,
  v7190,
  v7191,
  v7192,
  v7193,
  v7194,
  v7195,
  v7196,
  v7197,
  v7198,
  v7199,
  v7200,
  v7201,
  v7202,
  v7203,
  v7204,
  v7205,
  v7206,
  v7207,
  v7208,
  v7209,
  v7210,
  v7211,
  v7212,
  v7213,
  v7214,
  v7215,
  v7216,
  v7217,
  v7218,
  v7219,
  v7220,
  v7221,
  v7222,
  v7223,
  v7224,
  v7225,
  v7226,
  v7227,
  v7228,
  v7229,
  v7230,
  v7231,
  v7232,
  v7233,
  v7234,
  v7235,
  v7236,
  v7237,
  v7238,
  v7239,
  v7240,
  v7241,
  v7242,
  v7243,
  v7244,
  v7245,
  v7246,
  v7247,
  v7248,
  v7249,
  v7250,
  v7251,
  v7252,
  v7253,
  v7254,
  v7255,
  v7256,
  v7257,
  v7258,
  v7259,
  v7260,
  v7261,
  v7262,
  v7263,
  v7264,
  v7265,
  v7266,
  v7267,
  v7268,
  v7269,
  v7270,
  v7271,
  v7272,
  v7273,
  v7274,
  v7275,
  v7276,
  v7277,
  v7278,
  v7279,
  v7280,
  v7281,
  v7282,
  v7283,
  v7284,
  v7285,
  v7286,
  v7287,
  v7288,
  v7289,
  v7290,
  v7291,
  v7292,
  v7293,
  v7294,
  v7295,
  v7296,
  v7297,
  v7298,
  v7299,
  v7300,
  v7301,
  v7302,
  v7303,
  v7304,
  v7305,
  v7306,
  v7307,
  v7308,
  v7309,
  v7310,
  v7311,
  v7312,
  v7313,
  v7314,
  v7315,
  v7316,
  v7317,
  v7318,
  v7319,
  v7320,
  v7321,
  v7322,
  v7323,
  v7324,
  v7325,
  v7326,
  v7327,
  v7328,
  v7329,
  v7330,
  v7331,
  v7332,
  v7333,
  v7334,
  v7335,
  v7336,
  v7337,
  v7338,
  v7339,
  v7340,
  v7341,
  v7342,
  v7343,
  v7344,
  v7345,
  v7346,
  v7347,
  v7348,
  v7349,
  v7350,
  v7351,
  v7352,
  v7353,
  v7354,
  v7355,
  v7356,
  v7357,
  v7358,
  v7359,
  v7360,
  v7361,
  v7362,
  v7363,
  v7364,
  v7365,
  v7366,
  v7367,
  v7368,
  v7369,
  v7370,
  v7371,
  v7372,
  v7373,
  v7374,
  v7375,
  v7376,
  v7377,
  v7378,
  v7379,
  v7380,
  v7381,
  v7382,
  v7383,
  v7384,
  v7385,
  v7386,
  v7387,
  v7388,
  v7389,
  v7390,
  v7391,
  v7392,
  v7393,
  v7394,
  v7395,
  v7396,
  v7397,
  v7398,
  v7399,
  v7400,
  v7401,
  v7402,
  v7403,
  v7404,
  v7405,
  v7406,
  v7407,
  v7408,
  v7409,
  v7410,
  v7411,
  v7412,
  v7413,
  v7414,
  v7415,
  v7416,
  v7417,
  v7418,
  v7419,
  v7420,
  v7421,
  v7422,
  v7423,
  v7424,
  v7425,
  v7426,
  v7427,
  v7428,
  v7429,
  v7430,
  v7431,
  v7432,
  v7433,
  v7434,
  v7435,
  v7436,
  v7437,
  v7438,
  v7439,
  v7440,
  v7441,
  v7442,
  v7443,
  v7444,
  v7445,
  v7446,
  v7447,
  v7448,
  v7449,
  v7450,
  v7451,
  v7452,
  v7453,
  v7454,
  v7455,
  v7456,
  v7457,
  v7458,
  v7459,
  v7460,
  v7461,
  v7462,
  v7463,
  v7464,
  v7465,
  v7466,
  v7467,
  v7468,
  v7469,
  v7470,
  v7471,
  v7472,
  v7473,
  v7474,
  v7475,
  v7476,
  v7477,
  v7478,
  v7479,
  v7480,
  v7481,
  v7482,
  v7483,
  v7484,
  v7485,
  v7486,
  v7487,
  v7488,
  v7489,
  v7490,
  v7491,
  v7492,
  v7493,
  v7494,
  v7495,
  v7496,
  v7497,
  v7498,
  v7499,
  v7500,
  v7501,
  v7502,
  v7503,
  v7504,
  v7505,
  v7506,
  v7507,
  v7508,
  v7509,
  v7510,
  v7511,
  v7512,
  v7513,
  v7514,
  v7515,
  v7516,
  v7517,
  v7518,
  v7519,
  v7520,
  v7521,
  v7522,
  v7523,
  v7524,
  v7525,
  v7526,
  v7527,
  v7528,
  v7529,
  v7530,
  v7531,
  v7532,
  v7533,
  v7534,
  v7535,
  v7536,
  v7537,
  v7538,
  v7539,
  v7540,
  v7541,
  v7542,
  v7543,
  v7544,
  v7545,
  v7546,
  v7547,
  v7548,
  v7549,
  v7550,
  v7551,
  v7552,
  v7553,
  v7554,
  v7555,
  v7556,
  v7557,
  v7558,
  v7559,
  v7560,
  v7561,
  v7562,
  v7563,
  v7564,
  v7565,
  v7566,
  v7567,
  v7568,
  v7569,
  v7570,
  v7571,
  v7572,
  v7573,
  v7574,
  v7575,
  v7576,
  v7577,
  v7578,
  v7579,
  v7580,
  v7581,
  v7582,
  v7583,
  v7584,
  v7585,
  v7586,
  v7587,
  v7588,
  v7589,
  v7590,
  v7591,
  v7592,
  v7593,
  v7594,
  v7595,
  v7596,
  v7597,
  v7598,
  v7599,
  v7600,
  v7601,
  v7602,
  v7603,
  v7604,
  v7605,
  v7606,
  v7607,
  v7608,
  v7609,
  v7610,
  v7611,
  v7612,
  v7613,
  v7614,
  v7615,
  v7616,
  v7617,
  v7618,
  v7619,
  v7620,
  v7621,
  v7622,
  v7623,
  v7624,
  v7625,
  v7626,
  v7627,
  v7628,
  v7629,
  v7630,
  v7631,
  v7632,
  v7633,
  v7634,
  v7635,
  v7636,
  v7637,
  v7638,
  v7639,
  v7640,
  v7641,
  v7642,
  v7643,
  v7644,
  v7645,
  v7646,
  v7647,
  v7648,
  v7649,
  v7650,
  v7651,
  v7652,
  v7653,
  v7654,
  v7655,
  v7656,
  v7657,
  v7658,
  v7659,
  v7660,
  v7661,
  v7662,
  v7663,
  v7664,
  v7665,
  v7666,
  v7667,
  v7668,
  v7669,
  v7670,
  v7671,
  v7672,
  v7673,
  v7674,
  v7675,
  v7676,
  v7677,
  v7678,
  v7679,
  v7680,
  v7681,
  v7682,
  v7683,
  v7684,
  v7685,
  v7686,
  v7687,
  v7688,
  v7689,
  v7690,
  v7691,
  v7692,
  v7693,
  v7694,
  v7695,
  v7696,
  v7697,
  v7698,
  v7699,
  v7700,
  v7701,
  v7702,
  v7703,
  v7704,
  v7705,
  v7706,
  v7707,
  v7708,
  v7709,
  v7710,
  v7711,
  v7712,
  v7713,
  v7714,
  v7715,
  v7716,
  v7717,
  v7718,
  v7719,
  v7720,
  v7721,
  v7722,
  v7723,
  v7724,
  v7725,
  v7726,
  v7727,
  v7728,
  v7729,
  v7730,
  v7731,
  v7732,
  v7733,
  v7734,
  v7735,
  v7736,
  v7737,
  v7738,
  v7739,
  v7740,
  v7741,
  v7742,
  v7743,
  v7744,
  v7745,
  v7746,
  v7747,
  v7748,
  v7749,
  v7750,
  v7751,
  v7752,
  v7753,
  v7754,
  v7755,
  v7756,
  v7757,
  v7758,
  v7759,
  v7760,
  v7761,
  v7762,
  v7763,
  v7764,
  v7765,
  v7766,
  v7767,
  v7768,
  v7769,
  v7770,
  v7771,
  v7772,
  v7773,
  v7774,
  v7775,
  v7776,
  v7777,
  v7778,
  v7779,
  v7780,
  v7781,
  v7782,
  v7783,
  v7784,
  v7785,
  v7786,
  v7787,
  v7788,
  v7789,
  v7790,
  v7791,
  v7792,
  v7793,
  v7794,
  v7795,
  v7796,
  v7797,
  v7798,
  v7799,
  v7800,
  v7801,
  v7802,
  v7803,
  v7804,
  v7805,
  v7806,
  v7807,
  v7808,
  v7809,
  v7810,
  v7811,
  v7812,
  v7813,
  v7814,
  v7815,
  v7816,
  v7817,
  v7818,
  v7819,
  v7820,
  v7821,
  v7822,
  v7823,
  v7824,
  v7825,
  v7826,
  v7827,
  v7828,
  v7829,
  v7830,
  v7831,
  v7832,
  v7833,
  v7834,
  v7835,
  v7836,
  v7837,
  v7838,
  v7839,
  v7840,
  v7841,
  v7842,
  v7843,
  v7844,
  v7845,
  v7846,
  v7847,
  v7848,
  v7849,
  v7850,
  v7851,
  v7852,
  v7853,
  v7854,
  v7855,
  v7856,
  v7857,
  v7858,
  v7859,
  v7860,
  v7861,
  v7862,
  v7863,
  v7864,
  v7865,
  v7866,
  v7867,
  v7868,
  v7869,
  v7870,
  v7871,
  v7872,
  v7873,
  v7874,
  v7875,
  v7876,
  v7877,
  v7878,
  v7879,
  v7880,
  v7881,
  v7882,
  v7883,
  v7884,
  v7885,
  v7886,
  v7887,
  v7888,
  v7889,
  v7890,
  v7891,
  v7892,
  v7893,
  v7894,
  v7895,
  v7896,
  v7897,
  v7898,
  v7899,
  v7900,
  v7901,
  v7902,
  v7903,
  v7904,
  v7905,
  v7906,
  v7907,
  v7908,
  v7909,
  v7910,
  v7911,
  v7912,
  v7913,
  v7914,
  v7915,
  v7916,
  v7917,
  v7918,
  v7919,
  v7920,
  v7921,
  v7922,
  v7923,
  v7924,
  v7925,
  v7926,
  v7927,
  v7928,
  v7929,
  v7930,
  v7931,
  v7932,
  v7933,
  v7934,
  v7935,
  v7936,
  v7937,
  v7938,
  v7939,
  v7940,
  v7941,
  v7942,
  v7943,
  v7944,
  v7945,
  v7946,
  v7947,
  v7948,
  v7949,
  v7950,
  v7951,
  v7952,
  v7953,
  v7954,
  v7955,
  v7956,
  v7957,
  v7958,
  v7959,
  v7960,
  v7961,
  v7962,
  v7963,
  v7964,
  v7965,
  v7966,
  v7967,
  v7968,
  v7969,
  v7970,
  v7971,
  v7972,
  v7973,
  v7974,
  v7975,
  v7976,
  v7977,
  v7978,
  v7979,
  v7980,
  v7981,
  v7982,
  v7983,
  v7984,
  v7985,
  v7986,
  v7987,
  v7988,
  v7989,
  v7990,
  v7991,
  v7992,
  v7993,
  v7994,
  v7995,
  v7996,
  v7997,
  v7998,
  v7999,
  v8000,
  v8001,
  v8002,
  v8003,
  v8004,
  v8005,
  v8006,
  v8007,
  v8008,
  v8009,
  v8010,
  v8011,
  v8012,
  v8013,
  v8014,
  v8015,
  v8016,
  v8017,
  v8018,
  v8019,
  v8020,
  v8021,
  v8022,
  v8023,
  v8024,
  v8025,
  v8026,
  v8027,
  v8028,
  v8029,
  v8030,
  v8031,
  v8032,
  v8033,
  v8034,
  v8035,
  v8036,
  v8037,
  v8038,
  v8039,
  v8040,
  v8041,
  v8042,
  v8043,
  v8044,
  v8045,
  v8046,
  v8047,
  v8048,
  v8049,
  v8050,
  v8051,
  v8052,
  v8053,
  v8054,
  v8055,
  v8056,
  v8057,
  v8058,
  v8059,
  v8060,
  v8061,
  v8062,
  v8063,
  v8064,
  v8065,
  v8066,
  v8067,
  v8068,
  v8069,
  v8070,
  v8071,
  v8072,
  v8073,
  v8074,
  v8075,
  v8076,
  v8077,
  v8078,
  v8079,
  v8080,
  v8081,
  v8082,
  v8083,
  v8084,
  v8085,
  v8086,
  v8087,
  v8088,
  v8089,
  v8090,
  v8091,
  v8092,
  v8093,
  v8094,
  v8095,
  v8096,
  v8097,
  v8098,
  v8099,
  v8100,
  v8101,
  v8102,
  v8103,
  v8104,
  v8105,
  v8106,
  v8107,
  v8108,
  v8109,
  v8110,
  v8111,
  v8112,
  v8113,
  v8114,
  v8115,
  v8116,
  v8117,
  v8118,
  v8119,
  v8120,
  v8121,
  v8122,
  v8123,
  v8124,
  v8125,
  v8126,
  v8127,
  v8128,
  v8129,
  v8130,
  v8131,
  v8132,
  v8133,
  v8134,
  v8135,
  v8136,
  v8137,
  v8138,
  v8139,
  v8140,
  v8141,
  v8142,
  v8143,
  v8144,
  v8145,
  v8146,
  v8147,
  v8148,
  v8149,
  v8150,
  v8151,
  v8152,
  v8153,
  v8154,
  v8155,
  v8156,
  v8157,
  v8158,
  v8159,
  v8160,
  v8161,
  v8162,
  v8163,
  v8164,
  v8165,
  v8166,
  v8167,
  v8168,
  v8169,
  v8170,
  v8171,
  v8172,
  v8173,
  v8174,
  v8175,
  v8176,
  v8177,
  v8178,
  v8179,
  v8180,
  v8181,
  v8182,
  v8183,
  v8184,
  v8185,
  v8186,
  v8187,
  v8188,
  v8189,
  v8190,
  v8191,
  v8192,
  v8193,
  v8194,
  v8195,
  v8196,
  v8197,
  v8198,
  v8199,
  v8200,
  v8201,
  v8202,
  v8203,
  v8204,
  v8205,
  v8206,
  v8207,
  v8208,
  v8209,
  v8210,
  v8211,
  v8212,
  v8213,
  v8214,
  v8215,
  v8216,
  v8217,
  v8218,
  v8219,
  v8220,
  v8221,
  v8222,
  v8223,
  v8224,
  v8225,
  v8226,
  v8227,
  v8228,
  v8229,
  v8230,
  v8231,
  v8232,
  v8233,
  v8234,
  v8235,
  v8236,
  v8237,
  v8238,
  v8239,
  v8240,
  v8241,
  v8242,
  v8243,
  v8244,
  v8245,
  v8246,
  v8247,
  v8248,
  v8249,
  v8250,
  v8251,
  v8252,
  v8253,
  v8254,
  v8255,
  v8256,
  v8257,
  v8258,
  v8259,
  v8260,
  v8261,
  v8262,
  v8263,
  v8264,
  v8265,
  v8266,
  v8267,
  v8268,
  v8269,
  v8270,
  v8271,
  v8272,
  v8273,
  v8274,
  v8275,
  v8276,
  v8277,
  v8278,
  v8279,
  v8280,
  v8281,
  v8282,
  v8283,
  v8284,
  v8285,
  v8286,
  v8287,
  v8288,
  v8289,
  v8290,
  v8291,
  v8292,
  v8293,
  v8294,
  v8295,
  v8296,
  v8297,
  v8298,
  v8299,
  v8300,
  v8301,
  v8302,
  v8303,
  v8304,
  v8305,
  v8306,
  v8307,
  v8308,
  v8309,
  v8310,
  v8311,
  v8312,
  v8313,
  v8314,
  v8315,
  v8316,
  v8317,
  v8318,
  v8319,
  v8320,
  v8321,
  v8322,
  v8323,
  v8324,
  v8325,
  v8326,
  v8327,
  v8328,
  v8329,
  v8330,
  v8331,
  v8332,
  v8333,
  v8334,
  v8335,
  v8336,
  v8337,
  v8338,
  v8339,
  v8340,
  v8341,
  v8342,
  v8343,
  v8344,
  v8345,
  v8346,
  v8347,
  v8348,
  v8349,
  v8350,
  v8351,
  v8352,
  v8353,
  v8354,
  v8355,
  v8356,
  v8357,
  v8358,
  v8359,
  v8360,
  v8361,
  v8362,
  v8363,
  v8364,
  v8365,
  v8366,
  v8367,
  v8368,
  v8369,
  v8370,
  v8371,
  v8372,
  v8373,
  v8374,
  v8375,
  v8376,
  v8377,
  v8378,
  v8379,
  v8380,
  v8381,
  v8382,
  v8383,
  v8384,
  v8385,
  v8386,
  v8387,
  v8388,
  v8389,
  v8390,
  v8391,
  v8392,
  v8393,
  v8394,
  v8395,
  v8396,
  v8397,
  v8398,
  v8399,
  v100,
  v101,
  v102,
  v103,
  v104,
  v105,
  v106,
  v107,
  v108,
  v109,
  v110,
  v111,
  v112,
  v113,
  v114,
  v115,
  v116,
  v117,
  v118,
  v119,
  v120,
  v121,
  v122,
  v123,
  v124,
  v125,
  v126,
  v127,
  v128,
  v129,
  v130,
  v131,
  v132,
  v133,
  v134,
  v135,
  v136,
  v137,
  v138,
  v139,
  v8400,
  v8401,
  v8402,
  v8403,
  v8404,
  v8405,
  v8406,
  v140,
  v8407,
  v141,
  v8408,
  v142,
  v8409,
  v143,
  v144,
  v145,
  v146,
  v147,
  v148,
  v149,
  v8410,
  v8411,
  v8412,
  v8413,
  v8414,
  v8415,
  v8416,
  v150,
  v8417,
  v151,
  v8418,
  v152,
  v8419,
  v153,
  v154,
  v155,
  v156,
  v157,
  v158,
  v159,
  v8420,
  v8421,
  v8422,
  v8423,
  v8424,
  v8425,
  v8426,
  v160,
  v8427,
  v161,
  v8428,
  v162,
  v8429,
  v163,
  v164,
  v165,
  v166,
  v167,
  v168,
  v169,
  v8430,
  v8431,
  v8432,
  v8433,
  v8434,
  v8435,
  v8436,
  v170,
  v8437,
  v171,
  v8438,
  v172,
  v8439,
  v173,
  v174,
  v175,
  v176,
  v177,
  v178,
  v179,
  v8440,
  v8441,
  v8442,
  v8443,
  v8444,
  v8445,
  v8446,
  v180,
  v8447,
  v181,
  v8448,
  v182,
  v8449,
  v183,
  v184,
  v185,
  v186,
  v187,
  v188,
  v189,
  v8450,
  v8451,
  v8452,
  v8453,
  v8454,
  v8455,
  v8456,
  v190,
  v8457,
  v191,
  v8458,
  v192,
  v8459,
  v193,
  v194,
  v195,
  v196,
  v197,
  v198,
  v199,
  v8460,
  v8461,
  v8462,
  v8463,
  v8464,
  v8465,
  v8466,
  v8467,
  v8468,
  v8469,
  v8470,
  v8471,
  v8472,
  v8473,
  v8474,
  v8475,
  v8476,
  v8477,
  v8478,
  v8479,
  v8480,
  v8481,
  v8482,
  v8483,
  v8484,
  v8485,
  v8486,
  v8487,
  v8488,
  v8489,
  v8490,
  v8491,
  v8492,
  v8493,
  v8494,
  v8495,
  v8496,
  v8497,
  v8498,
  v8499,
  v200,
  v201,
  v202,
  v203,
  v204,
  v205,
  v206,
  v207,
  v208,
  v209,
  v210,
  v211,
  v212,
  v213,
  v214,
  v215,
  v216,
  v217,
  v218,
  v219,
  v220,
  v221,
  v222,
  v223,
  v224,
  v225,
  v226,
  v227,
  v228,
  v229,
  v230,
  v231,
  v232,
  v233,
  v234,
  v235,
  v236,
  v237,
  v238,
  v239,
  v8500,
  v8501,
  v8502,
  v8503,
  v8504,
  v8505,
  v8506,
  v240,
  v8507,
  v241,
  v8508,
  v242,
  v8509,
  v243,
  v244,
  v245,
  v246,
  v247,
  v248,
  v249,
  v8510,
  v8511,
  v8512,
  v8513,
  v8514,
  v8515,
  v8516,
  v250,
  v8517,
  v251,
  v8518,
  v252,
  v8519,
  v253,
  v254,
  v255,
  v256,
  v257,
  v258,
  v259,
  v8520,
  v8521,
  v8522,
  v8523,
  v8524,
  v8525,
  v8526,
  v260,
  v8527,
  v261,
  v8528,
  v262,
  v8529,
  v263,
  v264,
  v265,
  v266,
  v267,
  v268,
  v269,
  v8530,
  v8531,
  v8532,
  v8533,
  v8534,
  v8535,
  v8536,
  v270,
  v8537,
  v271,
  v8538,
  v272,
  v8539,
  v273,
  v274,
  v275,
  v276,
  v277,
  v278,
  v279,
  v8540,
  v8541,
  v8542,
  v8543,
  v8544,
  v8545,
  v8546,
  v280,
  v8547,
  v281,
  v8548,
  v282,
  v8549,
  v283,
  v284,
  v285,
  v286,
  v287,
  v288,
  v289,
  v8550,
  v8551,
  v8552,
  v8553,
  v8554,
  v8555,
  v8556,
  v290,
  v8557,
  v291,
  v8558,
  v292,
  v8559,
  v293,
  v294,
  v295,
  v296,
  v297,
  v298,
  v299,
  v8560,
  v8561,
  v8562,
  v8563,
  v8564,
  v8565,
  v8566,
  v8567,
  v8568,
  v8569,
  v8570,
  v8571,
  v8572,
  v8573,
  v8574,
  v8575,
  v8576,
  v8577,
  v8578,
  v8579,
  v8580,
  v8581,
  v8582,
  v8583,
  v8584,
  v8585,
  v8586,
  v8587,
  v8588,
  v8589,
  v8590,
  v8591,
  v8592,
  v8593,
  v8594,
  v8595,
  v8596,
  v8597,
  v8598,
  v8599,
  v300,
  v301,
  v302,
  v303,
  v304,
  v305,
  v306,
  v307,
  v308,
  v309,
  v310,
  v311,
  v312,
  v313,
  v314,
  v315,
  v316,
  v317,
  v318,
  v319,
  v320,
  v321,
  v322,
  v323,
  v324,
  v325,
  v326,
  v327,
  v328,
  v329,
  v330,
  v331,
  v332,
  v333,
  v334,
  v335,
  v336,
  v337,
  v338,
  v339,
  v8600,
  v8601,
  v8602,
  v8603,
  v8604,
  v8605,
  v8606,
  v340,
  v8607,
  v341,
  v8608,
  v342,
  v8609,
  v343,
  v344,
  v345,
  v346,
  v347,
  v348,
  v349,
  v8610,
  v8611,
  v8612,
  v8613,
  v8614,
  v8615,
  v8616,
  v350,
  v8617,
  v351,
  v8618,
  v352,
  v8619,
  v353,
  v354,
  v355,
  v356,
  v357,
  v358,
  v359,
  v8620,
  v8621,
  v8622,
  v8623,
  v8624,
  v8625,
  v8626,
  v360,
  v8627,
  v361,
  v8628,
  v362,
  v8629,
  v363,
  v364,
  v365,
  v366,
  v367,
  v368,
  v369,
  v8630,
  v8631,
  v8632,
  v8633,
  v8634,
  v8635,
  v8636,
  v370,
  v8637,
  v371,
  v8638,
  v372,
  v8639,
  v373,
  v374,
  v375,
  v376,
  v377,
  v378,
  v379,
  v8640,
  v8641,
  v8642,
  v8643,
  v8644,
  v8645,
  v8646,
  v380,
  v8647,
  v381,
  v8648,
  v382,
  v8649,
  v383,
  v384,
  v385,
  v386,
  v387,
  v388,
  v389,
  v8650,
  v8651,
  v8652,
  v8653,
  v8654,
  v8655,
  v8656,
  v390,
  v8657,
  v391,
  v8658,
  v392,
  v8659,
  v393,
  v394,
  v395,
  v396,
  v397,
  v398,
  v399,
  v8660,
  v8661,
  v8662,
  v8663,
  v8664,
  v8665,
  v8666,
  v8667,
  v8668,
  v8669,
  v8670,
  v8671,
  v8672,
  v8673,
  v8674,
  v8675,
  v8676,
  v8677,
  v8678,
  v8679,
  v8680,
  v8681,
  v8682,
  v8683,
  v8684,
  v8685,
  v8686,
  v8687,
  v8688,
  v8689,
  v8690,
  v8691,
  v8692,
  v8693,
  v8694,
  v8695,
  v8696,
  v8697,
  v8698,
  v8699,
  v400,
  v401,
  v402,
  v403,
  v404,
  v405,
  v406,
  v407,
  v408,
  v409,
  v410,
  v411,
  v412,
  v413,
  v414,
  v415,
  v416,
  v417,
  v418,
  v419,
  v420,
  v421,
  v422,
  v423,
  v424,
  v425,
  v426,
  v427,
  v428,
  v429,
  v430,
  v431,
  v432,
  v433,
  v434,
  v435,
  v436,
  v437,
  v438,
  v439,
  v8700,
  v8701,
  v8702,
  v8703,
  v8704,
  v8705,
  v8706,
  v440,
  v8707,
  v441,
  v8708,
  v442,
  v8709,
  v443,
  v444,
  v445,
  v446,
  v447,
  v448,
  v449,
  v8710,
  v8711,
  v8712,
  v8713,
  v8714,
  v8715,
  v8716,
  v450,
  v8717,
  v451,
  v8718,
  v452,
  v8719,
  v453,
  v454,
  v455,
  v456,
  v457,
  v458,
  v459,
  v8720,
  v8721,
  v8722,
  v8723,
  v8724,
  v8725,
  v8726,
  v460,
  v8727,
  v461,
  v8728,
  v462,
  v8729,
  v463,
  v464,
  v465,
  v466,
  v467,
  v468,
  v469,
  v8730,
  v8731,
  v8732,
  v8733,
  v8734,
  v8735,
  v8736,
  v470,
  v8737,
  v471,
  v8738,
  v472,
  v8739,
  v473,
  v474,
  v475,
  v476,
  v477,
  v478,
  v479,
  v8740,
  v8741,
  v8742,
  v8743,
  v8744,
  v8745,
  v8746,
  v480,
  v8747,
  v481,
  v8748,
  v482,
  v8749,
  v483,
  v484,
  v485,
  v486,
  v487,
  v488,
  v489,
  v8750,
  v8751,
  v8752,
  v8753,
  v8754,
  v8755,
  v8756,
  v490,
  v8757,
  v491,
  v8758,
  v492,
  v8759,
  v493,
  v494,
  v495,
  v496,
  v497,
  v498,
  v499,
  v8760,
  v8761,
  v8762,
  v8763,
  v8764,
  v8765,
  v8766,
  v8767,
  v8768,
  v8769,
  v8770,
  v8771,
  v8772,
  v8773,
  v8774,
  v8775,
  v8776,
  v8777,
  v8778,
  v8779,
  v8780,
  v8781,
  v8782,
  v8783,
  v8784,
  v8785,
  v8786,
  v8787,
  v8788,
  v8789,
  v8790,
  v8791,
  v8792,
  v8793,
  v8794,
  v8795,
  v8796,
  v8797,
  v8798,
  v8799,
  v500,
  v501,
  v502,
  v503,
  v504,
  v505,
  v506,
  v507,
  v508,
  v509,
  v510,
  v511,
  v512,
  v513,
  v514,
  v515,
  v516,
  v517,
  v518,
  v519,
  v520,
  v521,
  v522,
  v523,
  v524,
  v525,
  v526,
  v527,
  v528,
  v529,
  v530,
  v531,
  v532,
  v533,
  v534,
  v535,
  v536,
  v537,
  v538,
  v539,
  v8800,
  v8801,
  v8802,
  v8803,
  v8804,
  v8805,
  v8806,
  v540,
  v8807,
  v541,
  v8808,
  v542,
  v8809,
  v543,
  v544,
  v545,
  v546,
  v547,
  v548,
  v549,
  v8810,
  v8811,
  v8812,
  v8813,
  v8814,
  v8815,
  v8816,
  v550,
  v8817,
  v551,
  v8818,
  v552,
  v8819,
  v553,
  v554,
  v555,
  v556,
  v557,
  v558,
  v559,
  v8820,
  v8821,
  v8822,
  v8823,
  v8824,
  v8825,
  v8826,
  v560,
  v8827,
  v561,
  v8828,
  v562,
  v8829,
  v563,
  v564,
  v565,
  v566,
  v567,
  v568,
  v569,
  v8830,
  v8831,
  v8832,
  v8833,
  v8834,
  v8835,
  v8836,
  v570,
  v8837,
  v571,
  v8838,
  v572,
  v8839,
  v573,
  v574,
  v575,
  v576,
  v577,
  v578,
  v579,
  v8840,
  v8841,
  v8842,
  v8843,
  v8844,
  v8845,
  v8846,
  v580,
  v8847,
  v581,
  v8848,
  v582,
  v8849,
  v583,
  v584,
  v585,
  v586,
  v587,
  v588,
  v589,
  v8850,
  v8851,
  v8852,
  v8853,
  v8854,
  v8855,
  v8856,
  v590,
  v8857,
  v591,
  v8858,
  v592,
  v8859,
  v593,
  v594,
  v595,
  v596,
  v597,
  v598,
  v599,
  v8860,
  v8861,
  v8862,
  v8863,
  v8864,
  v8865,
  v8866,
  v8867,
  v8868,
  v8869,
  v8870,
  v8871,
  v8872,
  v8873,
  v8874,
  v8875,
  v8876,
  v8877,
  v8878,
  v8879,
  v8880,
  v8881,
  v8882,
  v8883,
  v8884,
  v8885,
  v8886,
  v8887,
  v8888,
  v8889,
  v8890,
  v8891,
  v8892,
  v8893,
  v8894,
  v8895,
  v8896,
  v8897,
  v8898,
  v8899,
  v600,
  v601,
  v602,
  v603,
  v604,
  v605,
  v606,
  v607,
  v608,
  v609,
  v610,
  v611,
  v612,
  v613,
  v614,
  v615,
  v616,
  v617,
  v618,
  v619,
  v620,
  v621,
  v622,
  v623,
  v624,
  v625,
  v626,
  v627,
  v628,
  v629,
  v630,
  v631,
  v632,
  v633,
  v634,
  v635,
  v636,
  v637,
  v638,
  v639,
  v8900,
  v8901,
  v8902,
  v8903,
  v8904,
  v8905,
  v8906,
  v640,
  v8907,
  v641,
  v8908,
  v642,
  v8909,
  v643,
  v644,
  v645,
  v646,
  v647,
  v648,
  v649,
  v8910,
  v8911,
  v8912,
  v8913,
  v8914,
  v8915,
  v8916,
  v650,
  v8917,
  v651,
  v8918,
  v652,
  v8919,
  v653,
  v654,
  v655,
  v656,
  v657,
  v658,
  v659,
  v8920,
  v8921,
  v8922,
  v8923,
  v8924,
  v8925,
  v8926,
  v660,
  v8927,
  v661,
  v8928,
  v662,
  v8929,
  v663,
  v664,
  v665,
  v666,
  v667,
  v668,
  v669,
  v8930,
  v8931,
  v8932,
  v8933,
  v8934,
  v8935,
  v8936,
  v670,
  v8937,
  v671,
  v8938,
  v672,
  v8939,
  v673,
  v674,
  v675,
  v676,
  v677,
  v678,
  v679,
  v8940,
  v8941,
  v8942,
  v8943,
  v8944,
  v8945,
  v8946,
  v680,
  v8947,
  v681,
  v8948,
  v682,
  v8949,
  v683,
  v684,
  v685,
  v686,
  v687,
  v688,
  v689,
  v8950,
  v8951,
  v8952,
  v8953,
  v8954,
  v8955,
  v8956,
  v690,
  v8957,
  v691,
  v8958,
  v692,
  v8959,
  v693,
  v694,
  v695,
  v696,
  v697,
  v698,
  v699,
  v8960,
  v8961,
  v8962,
  v8963,
  v8964,
  v8965,
  v8966,
  v8967,
  v8968,
  v8969,
  v8970,
  v8971,
  v8972,
  v8973,
  v8974,
  v8975,
  v8976,
  v8977,
  v8978,
  v8979,
  v8980,
  v8981,
  v8982,
  v8983,
  v8984,
  v8985,
  v8986,
  v8987,
  v8988,
  v8989,
  v8990,
  v8991,
  v8992,
  v8993,
  v8994,
  v8995,
  v8996,
  v8997,
  v8998,
  v8999,
  v700,
  v701,
  v702,
  v703,
  v704,
  v705,
  v706,
  v707,
  v708,
  v709,
  v710,
  v711,
  v712,
  v713,
  v714,
  v715,
  v716,
  v717,
  v718,
  v719,
  v720,
  v721,
  v722,
  v723,
  v724,
  v725,
  v726,
  v727,
  v728,
  v729,
  v730,
  v731,
  v732,
  v733,
  v734,
  v735,
  v736,
  v737,
  v738,
  v739,
  v740,
  v741,
  v742,
  v743,
  v744,
  v745,
  v746,
  v747,
  v748,
  v749,
  v750,
  v751,
  v752,
  v753,
  v754,
  v755,
  v756,
  v757,
  v758,
  v759,
  v760,
  v761,
  v762,
  v763,
  v764,
  v765,
  v766,
  v767,
  v768,
  v769,
  v770,
  v771,
  v772,
  v773,
  v774,
  v775,
  v776,
  v777,
  v778,
  v779,
  v780,
  v781,
  v782,
  v783,
  v784,
  v785,
  v786,
  v787,
  v788,
  v789,
  v790,
  v791,
  v792,
  v793,
  v794,
  v795,
  v796,
  v797,
  v798,
  v799,
  v800,
  v801,
  v802,
  v803,
  v804,
  v805,
  v806,
  v807,
  v808,
  v809,
  v810,
  v811,
  v812,
  v813,
  v814,
  v815,
  v816,
  v817,
  v818,
  v819,
  v820,
  v821,
  v822,
  v823,
  v824,
  v825,
  v826,
  v827,
  v828,
  v829,
  v830,
  v831,
  v832,
  v833,
  v834,
  v835,
  v836,
  v837,
  v838,
  v839,
  v840,
  v841,
  v842,
  v843,
  v844,
  v845,
  v846,
  v847,
  v848,
  v849,
  v850,
  v851,
  v852,
  v853,
  v854,
  v855,
  v856,
  v857,
  v858,
  v859,
  v860,
  v861,
  v862,
  v863,
  v864,
  v865,
  v866,
  v867,
  v868,
  v869,
  v870,
  v871,
  v872,
  v873,
  v874,
  v875,
  v876,
  v877,
  v878,
  v879,
  v880,
  v881,
  v882,
  v883,
  v884,
  v885,
  v886,
  v887,
  v888,
  v889,
  v890,
  v891,
  v892,
  v893,
  v894,
  v895,
  v896,
  v897,
  v898,
  v899,
  v900,
  v901,
  v902,
  v903,
  v904,
  v905,
  v906,
  v907,
  v908,
  v909,
  v910,
  v911,
  v912,
  v913,
  v914,
  v915,
  v916,
  v917,
  v918,
  v919,
  v920,
  v921,
  v922,
  v923,
  v924,
  v925,
  v926,
  v927,
  v928,
  v929,
  v930,
  v931,
  v932,
  v933,
  v934,
  v935,
  v936,
  v937,
  v938,
  v939,
  v940,
  v941,
  v942,
  v943,
  v944,
  v945,
  v946,
  v947,
  v948,
  v949,
  v950,
  v951,
  v952,
  v953,
  v954,
  v955,
  v956,
  v957,
  v958,
  v959,
  v960,
  v961,
  v962,
  v963,
  v964,
  v965,
  v966,
  v967,
  v968,
  v969,
  v970,
  v971,
  v972,
  v973,
  v974,
  v975,
  v976,
  v977,
  v978,
  v979,
  v980,
  v981,
  v982,
  v983,
  v984,
  v985,
  v986,
  v987,
  v988,
  v989,
  v990,
  v991,
  v992,
  v993,
  v994,
  v995,
  v996,
  v997,
  v998,
  v999,
  v9000,
  v9001,
  v9002,
  v9003,
  v9004,
  v9005,
  v9006,
  v9007,
  v9008,
  v9009,
  v9010,
  v9011,
  v9012,
  v9013,
  v9014,
  v9015,
  v9016,
  v9017,
  v9018,
  v9019,
  v9020,
  v9021,
  v9022,
  v9023,
  v9024,
  v9025,
  v9026,
  v9027,
  v9028,
  v9029,
  v9030,
  v9031,
  v9032,
  v9033,
  v9034,
  v9035,
  v9036,
  v9037,
  v9038,
  v9039,
  v9040,
  v9041,
  v9042,
  v9043,
  v9044,
  v9045,
  v9046,
  v9047,
  v9048,
  v9049,
  v9050,
  v9051,
  v9052,
  v9053,
  v9054,
  v9055,
  v9056,
  v9057,
  v9058,
  v9059,
  v9060,
  v9061,
  v9062,
  v9063,
  v9064,
  v9065,
  v9066,
  v9067,
  v9068,
  v9069,
  v9070,
  v9071,
  v9072,
  v9073,
  v9074,
  v9075,
  v9076,
  v9077,
  v9078,
  v9079,
  v9080,
  v9081,
  v9082,
  v9083,
  v9084,
  v9085,
  v9086,
  v9087,
  v9088,
  v9089,
  v9090,
  v9091,
  v9092,
  v9093,
  v9094,
  v9095,
  v9096,
  v9097,
  v9098,
  v9099,
  v9100,
  v9101,
  v9102,
  v9103,
  v9104,
  v9105,
  v9106,
  v9107,
  v9108,
  v9109,
  v9110,
  v9111,
  v9112,
  v9113,
  v9114,
  v9115,
  v9116,
  v9117,
  v9118,
  v9119,
  v9120,
  v9121,
  v9122,
  v9123,
  v9124,
  v9125,
  v9126,
  v9127,
  v9128,
  v9129,
  v9130,
  v9131,
  v9132,
  v9133,
  v9134,
  v9135,
  v9136,
  v9137,
  v9138,
  v9139,
  v9140,
  v9141,
  v9142,
  v9143,
  v9144,
  v9145,
  v9146,
  v9147,
  v9148,
  v9149,
  v9150,
  v9151,
  v9152,
  v9153,
  v9154,
  v9155,
  v9156,
  v9157,
  v9158,
  v9159,
  v9160,
  v9161,
  v9162,
  v9163,
  v9164,
  v9165,
  v9166,
  v9167,
  v9168,
  v9169,
  v9170,
  v9171,
  v9172,
  v9173,
  v9174,
  v9175,
  v9176,
  v9177,
  v9178,
  v9179,
  v9180,
  v9181,
  v9182,
  v9183,
  v9184,
  v9185,
  v9186,
  v9187,
  v9188,
  v9189,
  v9190,
  v9191,
  v9192,
  v9193,
  v9194,
  v9195,
  v9196,
  v9197,
  v9198,
  v9199,
  v9200,
  v9201,
  v9202,
  v9203,
  v9204,
  v9205,
  v9206,
  v9207,
  v9208,
  v9209,
  v9210,
  v9211,
  v9212,
  v9213,
  v9214,
  v9215,
  v9216,
  v9217,
  v9218,
  v9219,
  v9220,
  v9221,
  v9222,
  v9223,
  v9224,
  v9225,
  v9226,
  v9227,
  v9228,
  v9229,
  v9230,
  v9231,
  v9232,
  v9233,
  v9234,
  v9235,
  v9236,
  v9237,
  v9238,
  v9239,
  v9240,
  v9241,
  v9242,
  v9243,
  v9244,
  v9245,
  v9246,
  v9247,
  v9248,
  v9249,
  v9250,
  v9251,
  v9252,
  v9253,
  v9254,
  v9255,
  v9256,
  v9257,
  v9258,
  v9259,
  v9260,
  v9261,
  v9262,
  v9263,
  v9264,
  v9265,
  v9266,
  v9267,
  v9268,
  v9269,
  v9270,
  v9271,
  v9272,
  v9273,
  v9274,
  v9275,
  v9276,
  v9277,
  v9278,
  v9279,
  v9280,
  v9281,
  v9282,
  v9283,
  v9284,
  v9285,
  v9286,
  v9287,
  v9288,
  v9289,
  v9290,
  v9291,
  v9292,
  v9293,
  v9294,
  v9295,
  v9296,
  v9297,
  v9298,
  v9299,
  v9300,
  v9301,
  v9302,
  v9303,
  v9304,
  v9305,
  v9306,
  v9307,
  v9308,
  v9309,
  v9310,
  v9311,
  v9312,
  v9313,
  v9314,
  v9315,
  v9316,
  v9317,
  v9318,
  v9319,
  v9320,
  v9321,
  v9322,
  v9323,
  v9324,
  v9325,
  v9326,
  v9327,
  v9328,
  v9329,
  v9330,
  v9331,
  v9332,
  v9333,
  v9334,
  v9335,
  v9336,
  v9337,
  v9338,
  v9339,
  v9340,
  v9341,
  v9342,
  v9343,
  v9344,
  v9345,
  v9346,
  v9347,
  v9348,
  v9349,
  v9350,
  v9351,
  v9352,
  v9353,
  v9354,
  v9355,
  v9356,
  v9357,
  v9358,
  v9359,
  v9360,
  v9361,
  v9362,
  v9363,
  v9364,
  v9365,
  v9366,
  v9367,
  v9368,
  v9369,
  v9370,
  v9371,
  v9372,
  v9373,
  v9374,
  v9375,
  v9376,
  v9377,
  v9378,
  v9379,
  v9380,
  v9381,
  v9382,
  v9383,
  v9384,
  v9385,
  v9386,
  v9387,
  v9388,
  v9389,
  v9390,
  v9391,
  v9392,
  v9393,
  v9394,
  v9395,
  v9396,
  v9397,
  v9398,
  v9399,
  v9400,
  v9401,
  v9402,
  v9403,
  v9404,
  v9405,
  v9406,
  v9407,
  v9408,
  v9409,
  v9410,
  v9411,
  v9412,
  v9413,
  v9414,
  v9415,
  v9416,
  v9417,
  v9418,
  v9419,
  v9420,
  v9421,
  v9422,
  v9423,
  v9424,
  v9425,
  v9426,
  v9427,
  v9428,
  v9429,
  v9430,
  v9431,
  v9432,
  v9433,
  v9434,
  v9435,
  v9436,
  v9437,
  v9438,
  v9439,
  v9440,
  v9441,
  v9442,
  v9443,
  v9444,
  v9445,
  v9446,
  v9447,
  v9448,
  v9449,
  v9450,
  v9451,
  v9452,
  v9453,
  v9454,
  v9455,
  v9456,
  v9457,
  v9458,
  v9459,
  v9460,
  v9461,
  v9462,
  v9463,
  v9464,
  v9465,
  v9466,
  v9467,
  v9468,
  v9469,
  v9470,
  v9471,
  v9472,
  v9473,
  v9474,
  v9475,
  v9476,
  v9477,
  v9478,
  v9479,
  v9480,
  v9481,
  v9482,
  v9483,
  v9484,
  v9485,
  v9486,
  v9487,
  v9488,
  v9489,
  v9490,
  v9491,
  v9492,
  v9493,
  v9494,
  v9495,
  v9496,
  v9497,
  v9498,
  v9499,
  v9500,
  v9501,
  v9502,
  v9503,
  v9504,
  v9505,
  v9506,
  v9507,
  v9508,
  v9509,
  v9510,
  v9511,
  v9512,
  v9513,
  v9514,
  v9515,
  v9516,
  v9517,
  v9518,
  v9519,
  v9520,
  v9521,
  v9522,
  v9523,
  v9524,
  v9525,
  v9526,
  v9527,
  v9528,
  v9529,
  v9530,
  v9531,
  v9532,
  v9533,
  v9534,
  v9535,
  v9536,
  v9537,
  v9538,
  v9539,
  v9540,
  v9541,
  v9542,
  v9543,
  v9544,
  v9545,
  v9546,
  v9547,
  v9548,
  v9549,
  v9550,
  v9551,
  v9552,
  v9553,
  v9554,
  v9555,
  v9556,
  v9557,
  v9558,
  v9559,
  v9560,
  v9561,
  v9562,
  v9563,
  v9564,
  v9565,
  v9566,
  v9567,
  v9568,
  v9569,
  v9570,
  v9571,
  v9572,
  v9573,
  v9574,
  v9575,
  v9576,
  v9577,
  v9578,
  v9579,
  v9580,
  v9581,
  v9582,
  v9583,
  v9584,
  v9585,
  v9586,
  v9587,
  v9588,
  v9589,
  v9590,
  v9591,
  v9592,
  v9593,
  v9594,
  v9595,
  v9596,
  v9597,
  v9598,
  v9599,
  v9600,
  v9601,
  v9602,
  v9603,
  v9604,
  v9605,
  v9606,
  v9607,
  v9608,
  v9609,
  v9610,
  v9611,
  v9612,
  v9613,
  v9614,
  v9615,
  v9616,
  v9617,
  v9618,
  v9619,
  v9620,
  v9621,
  v9622,
  v9623,
  v9624,
  v9625,
  v9626,
  v9627,
  v9628,
  v9629,
  v9630,
  v9631,
  v9632,
  v9633,
  v9634,
  v9635,
  v9636,
  v9637,
  v9638,
  v9639,
  v9640,
  v9641,
  v9642,
  v9643,
  v9644,
  v9645,
  v9646,
  v9647,
  v9648,
  v9649,
  v9650,
  v9651,
  v9652,
  v9653,
  v9654,
  v9655,
  v9656,
  v9657,
  v9658,
  v9659,
  v9660,
  v9661,
  v9662,
  v9663,
  v9664,
  v9665,
  v9666,
  v9667,
  v9668,
  v9669,
  v9670,
  v9671,
  v9672,
  v9673,
  v9674,
  v9675,
  v9676,
  v9677,
  v9678,
  v9679,
  v9680,
  v9681,
  v9682,
  v9683,
  v9684,
  v9685,
  v9686,
  v9687,
  v9688,
  v9689,
  v9690,
  v9691,
  v9692,
  v9693,
  v9694,
  v9695,
  v9696,
  v9697,
  v9698,
  v9699,
  v9700,
  v9701,
  v9702,
  v9703,
  v9704,
  v9705,
  v9706,
  v9707,
  v9708,
  v9709,
  v9710,
  v9711,
  v9712,
  v9713,
  v9714,
  v9715,
  v9716,
  v9717,
  v9718,
  v9719,
  v9720,
  v9721,
  v9722,
  v9723,
  v9724,
  v9725,
  v9726,
  v9727,
  v9728,
  v9729,
  v9730,
  v9731,
  v9732,
  v9733,
  v9734,
  v9735,
  v9736,
  v9737,
  v9738,
  v9739,
  v9740,
  v9741,
  v9742,
  v9743,
  v9744,
  v9745,
  v9746,
  v9747,
  v9748,
  v9749,
  v9750,
  v9751,
  v9752,
  v9753,
  v9754,
  v9755,
  v9756,
  v9757,
  v9758,
  v9759,
  v9760,
  v9761,
  v9762,
  v9763,
  v9764,
  v9765,
  v9766,
  v9767,
  v9768,
  v9769,
  v9770,
  v9771,
  v9772,
  v9773,
  v9774,
  v9775,
  v9776,
  v9777,
  v9778,
  v9779,
  v9780,
  v9781,
  v9782,
  v9783,
  v9784,
  v9785,
  v9786,
  v9787,
  v9788,
  v9789,
  v9790,
  v9791,
  v9792,
  v9793,
  v9794,
  v9795,
  v9796,
  v9797,
  v9798,
  v9799,
  v9800,
  v9801,
  v9802,
  v9803,
  v9804,
  v9805,
  v9806,
  v9807,
  v9808,
  v9809,
  v9810,
  v9811,
  v9812,
  v9813,
  v9814,
  v9815,
  v9816,
  v9817,
  v9818,
  v9819,
  v9820,
  v9821,
  v9822,
  v9823,
  v9824,
  v9825,
  v9826,
  v9827,
  v9828,
  v9829,
  v9830,
  v9831,
  v9832,
  v9833,
  v9834,
  v9835,
  v9836,
  v9837,
  v9838,
  v9839,
  v9840,
  v9841,
  v9842,
  v9843,
  v9844,
  v9845,
  v9846,
  v9847,
  v9848,
  v9849,
  v9850,
  v9851,
  v9852,
  v9853,
  v9854,
  v9855,
  v9856,
  v9857,
  v9858,
  v9859,
  v9860,
  v9861,
  v9862,
  v9863,
  v9864,
  v9865,
  v9866,
  v9867,
  v9868,
  v9869,
  v9870,
  v9871,
  v9872,
  v9873,
  v9874,
  v9875,
  v9876,
  v9877,
  v9878,
  v9879,
  v9880,
  v9881,
  v9882,
  v9883,
  v9884,
  v9885,
  v9886,
  v9887,
  v9888,
  v9889,
  v9890,
  v9891,
  v9892,
  v9893,
  v9894,
  v9895,
  v9896,
  v9897,
  v9898,
  v9899,
  v9900,
  v9901,
  v9902,
  v9903,
  v9904,
  v9905,
  v9906,
  v9907,
  v9908,
  v9909,
  v9910,
  v9911,
  v9912,
  v9913,
  v9914,
  v9915,
  v9916,
  v9917,
  v9918,
  v9919,
  v9920,
  v9921,
  v9922,
  v9923,
  v9924,
  v9925,
  v9926,
  v9927,
  v9928,
  v9929,
  v9930,
  v9931,
  v9932,
  v9933,
  v9934,
  v9935,
  v9936,
  v9937,
  v9938,
  v9939,
  v9940,
  v9941,
  v9942,
  v9943,
  v9944,
  v9945,
  v9946,
  v9947,
  v9948,
  v9949,
  v9950,
  v9951,
  v9952,
  v9953,
  v9954,
  v9955,
  v9956,
  v9957,
  v9958,
  v9959,
  v9960,
  v9961,
  v9962,
  v9963,
  v9964,
  v9965,
  v9966,
  v9967,
  v9968,
  v9969,
  v9970,
  v9971,
  v9972,
  v9973,
  v9974,
  v9975,
  v9976,
  v9977,
  v9978,
  v9979,
  v9980,
  v9981,
  v9982,
  v9983,
  v9984,
  v9985,
  v9986,
  v9987,
  v9988,
  v9989,
  v9990,
  v9991,
  v9992,
  v9993,
  v9994,
  v9995,
  v9996,
  v9997,
  v9998,
  v9999,
  v10,
  v11,
  v12,
  v13,
  v14,
  v15,
  v16,
  v17,
  v18,
  v19,
  v20,
  v21,
  v22,
  v23,
  v24,
  v25,
  v26,
  v27,
  v28,
  v29,
  v30,
  v31,
  v32,
  v33,
  v34,
  v35,
  v36,
  v37,
  v38,
  v39,
  v40,
  v41,
  v42,
  v43,
  v44,
  v45,
  v46,
  v47,
  v48,
  v49,
  v50,
  v51,
  v52,
  v53,
  v54,
  v55,
  v56,
  v57,
  v58,
  v59,
  v60,
  v61,
  v62,
  v63,
  v64,
  v65,
  v66,
  v67,
  v68,
  v69,
  v70,
  v71,
  v72,
  v73,
  v74,
  v75,
  v76,
  v77,
  v78,
  v79,
  v80,
  v81,
  v82,
  v83,
  v84,
  v85,
  v86,
  v87,
  v88,
  v89,
  v90,
  v91,
  v92,
  v93,
  v94,
  v95,
  v96,
  v97,
  v98,
  v99,
  v1000,
  v1001,
  v1002,
  v1003,
  v1004,
  v1005,
  v1006,
  v1007,
  v1008,
  v1009,
  v1010,
  v1011,
  v1012,
  v1013,
  v1014,
  v1015,
  v1016,
  v1017,
  v1018,
  v1019,
  v1020,
  v1021,
  v1022,
  v1023,
  v1024,
  v1025,
  v1026,
  v1027,
  v1028,
  v1029,
  v1030,
  v1031,
  v1032,
  v1033,
  v1034,
  v1035,
  v1036,
  v1037,
  v1038,
  v1039,
  v1040,
  v1041,
  v1042,
  v1043,
  v1044,
  v1045,
  v1046,
  v1047,
  v1048,
  v1049,
  v1050,
  v1051,
  v1052,
  v1053,
  v1054,
  v1055,
  v1056,
  v1057,
  v1058,
  v1059,
  v1060,
  v1061,
  v1062,
  v1063,
  v1064,
  v1065,
  v1066,
  v1067,
  v1068,
  v1069,
  v1070,
  v1071,
  v1072,
  v1073,
  v1074,
  v1075,
  v1076,
  v1077,
  v1078,
  v1079,
  v1080,
  v1081,
  v1082,
  v1083,
  v1084,
  v1085,
  v1086,
  v1087,
  v1088,
  v1089,
  v1090,
  v1091,
  v1092,
  v1093,
  v1094,
  v1095,
  v1096,
  v1097,
  v1098,
  v1099,
  v1100,
  v1101,
  v1102,
  v1103,
  v1104,
  v1105,
  v1106,
  v1107,
  v1108,
  v1109,
  v1110,
  v1111,
  v1112,
  v1113,
  v1114,
  v1115,
  v1116,
  v1117,
  v1118,
  v1119,
  v1120,
  v1121,
  v1122,
  v1123,
  v1124,
  v1125,
  v1126,
  v1127,
  v1128,
  v1129,
  v1130,
  v1131,
  v1132,
  v1133,
  v1134,
  v1135,
  v1136,
  v1137,
  v1138,
  v1139,
  v1140,
  v1141,
  v1142,
  v1143,
  v1144,
  v1145,
  v1146,
  v1147,
  v1148,
  v1149,
  v1150,
  v1151,
  v1152,
  v1153,
  v1154,
  v1155,
  v1156,
  v1157,
  v1158,
  v1159,
  v1160,
  v1161,
  v1162,
  v1163,
  v1164,
  v1165,
  v1166,
  v1167,
  v1168,
  v1169,
  v1170,
  v1171,
  v1172,
  v1173,
  v1174,
  v1175,
  v1176,
  v1177,
  v1178,
  v1179,
  v1180,
  v1181,
  v1182,
  v1183,
  v1184,
  v1185,
  v1186,
  v1187,
  v1188,
  v1189,
  v1190,
  v1191,
  v1192,
  v1193,
  v1194,
  v1195,
  v1196,
  v1197,
  v1198,
  v1199,
  v1200,
  v1201,
  v1202,
  v1203,
  v1204,
  v1205,
  v1206,
  v1207,
  v1208,
  v1209,
  v1210,
  v1211,
  v1212,
  v1213,
  v1214,
  v1215,
  v1216,
  v1217,
  v1218,
  v1219,
  v1220,
  v1221,
  v1222,
  v1223,
  v1224,
  v1225,
  v1226,
  v1227,
  v1228,
  v1229,
  v1230,
  v1231,
  v1232,
  v1233,
  v1234,
  v1235,
  v1236,
  v1237,
  v1238,
  v1239,
  v1240,
  v1241,
  v1242,
  v1243,
  v1244,
  v1245,
  v1246,
  v1247,
  v1248,
  v1249,
  v1250,
  v1251,
  v1252,
  v1253,
  v1254,
  v1255,
  v1256,
  v1257,
  v1258,
  v1259,
  v1260,
  v1261,
  v1262,
  v1263,
  v1264,
  v1265,
  v1266,
  v1267,
  v1268,
  v1269,
  v1270,
  v1271,
  v1272,
  v1273,
  v1274,
  v1275,
  v1276,
  v1277,
  v1278,
  v1279,
  v1280,
  v1281,
  v1282,
  v1283,
  v1284,
  v1285,
  v1286,
  v1287,
  v1288,
  v1289,
  v1290,
  v1291,
  v1292,
  v1293,
  v1294,
  v1295,
  v1296,
  v1297,
  v1298,
  v1299,
  v1300,
  v1301,
  v1302,
  v1303,
  v1304,
  v1305,
  v1306,
  v1307,
  v1308,
  v1309,
  v1310,
  v1311,
  v1312,
  v1313,
  v1314,
  v1315,
  v1316,
  v1317,
  v1318,
  v1319,
  v1320,
  v1321,
  v1322,
  v1323,
  v1324,
  v1325,
  v1326,
  v1327,
  v1328,
  v1329,
  v1330,
  v1331,
  v1332,
  v1333,
  v1334,
  v1335,
  v1336,
  v1337,
  v1338,
  v1339,
  v1340,
  v1341,
  v1342,
  v1343,
  v1344,
  v1345,
  v1346,
  v1347,
  v1348,
  v1349,
  v1350,
  v1351,
  v1352,
  v1353,
  v1354,
  v1355,
  v1356,
  v1357,
  v1358,
  v1359,
  v1360,
  v1361,
  v1362,
  v1363,
  v1364,
  v1365,
  v1366,
  v1367,
  v1368,
  v1369,
  v1370,
  v1371,
  v1372,
  v1373,
  v1374,
  v1375,
  v1376,
  v1377,
  v1378,
  v1379,
  v1380,
  v1381,
  v1382,
  v1383,
  v1384,
  v1385,
  v1386,
  v1387,
  v1388,
  v1389,
  v1390,
  v1391,
  v1392,
  v1393,
  v1394,
  v1395,
  v1396,
  v1397,
  v1398,
  v1399,
  v1400,
  v1401,
  v1402,
  v1403,
  v1404,
  v1405,
  v1406,
  v1407,
  v1408,
  v1409,
  v1410,
  v1411,
  v1412,
  v1413,
  v1414,
  v1415,
  v1416,
  v1417,
  v1418,
  v1419,
  v1420,
  v1421,
  v1422,
  v1423,
  v1424,
  v1425,
  v1426,
  v1427,
  v1428,
  v1429,
  v1430,
  v1431,
  v1432,
  v1433,
  v1434,
  v1435,
  v1436,
  v1437,
  v1438,
  v1439,
  v1440,
  v1441,
  v1442,
  v1443,
  v1444,
  v1445,
  v1446,
  v1447,
  v1448,
  v1449,
  v1450,
  v1451,
  v1452,
  v1453,
  v1454,
  v1455,
  v1456,
  v1457,
  v1458,
  v1459,
  v1460,
  v1461,
  v1462,
  v1463,
  v1464,
  v1465,
  v1466,
  v1467,
  v1468,
  v1469,
  v1470,
  v1471,
  v1472,
  v1473,
  v1474,
  v1475,
  v1476,
  v1477,
  v1478,
  v1479,
  v1480,
  v1481,
  v1482,
  v1483,
  v1484,
  v1485,
  v1486,
  v1487,
  v1488,
  v1489,
  v1490,
  v1491,
  v1492,
  v1493,
  v1494,
  v1495,
  v1496,
  v1497,
  v1498,
  v1499,
  v1500,
  v1501,
  v1502,
  v1503,
  v1504,
  v1505,
  v1506,
  v1507,
  v1508,
  v1509,
  v1510,
  v1511,
  v1512,
  v1513,
  v1514,
  v1515,
  v1516,
  v1517,
  v1518,
  v1519,
  v1520,
  v1521,
  v1522,
  v1523,
  v1524,
  v1525,
  v1526,
  v1527,
  v1528,
  v1529,
  v1530,
  v1531,
  v1532,
  v1533,
  v1534,
  v1535,
  v1536,
  v1537,
  v1538,
  v1539,
  v1540,
  v1541,
  v1542,
  v1543,
  v1544,
  v1545,
  v1546,
  v1547,
  v1548,
  v1549,
  v1550,
  v1551,
  v1552,
  v1553,
  v1554,
  v1555,
  v1556,
  v1557,
  v1558,
  v1559,
  v1560,
  v1561,
  v1562,
  v1563,
  v1564,
  v1565,
  v1566,
  v1567,
  v1568,
  v1569,
  v1570,
  v1571,
  v1572,
  v1573,
  v1574,
  v1575,
  v1576,
  v1577,
  v1578,
  v1579,
  v1580,
  v1581,
  v1582,
  v1583,
  v1584,
  v1585,
  v1586,
  v1587,
  v1588,
  v1589,
  v1590,
  v1591,
  v1592,
  v1593,
  v1594,
  v1595,
  v1596,
  v1597,
  v1598,
  v1599,
  v1600,
  v1601,
  v1602,
  v1603,
  v1604,
  v1605,
  v1606,
  v1607,
  v1608,
  v1609,
  v1610,
  v1611,
  v1612,
  v1613,
  v1614,
  v1615,
  v1616,
  v1617,
  v1618,
  v1619,
  v1620,
  v1621,
  v1622,
  v1623,
  v1624,
  v1625,
  v1626,
  v1627,
  v1628,
  v1629,
  v1630,
  v1631,
  v1632,
  v1633,
  v1634,
  v1635,
  v1636,
  v1637,
  v1638,
  v1639,
  v1640,
  v1641,
  v1642,
  v1643,
  v1644,
  v1645,
  v1646,
  v1647,
  v1648,
  v1649,
  v1650,
  v1651,
  v1652,
  v1653,
  v1654,
  v1655,
  v1656,
  v1657,
  v1658,
  v1659,
  v1660,
  v1661,
  v1662,
  v1663,
  v1664,
  v1665,
  v1666,
  v1667,
  v1668,
  v1669,
  v1670,
  v1671,
  v1672,
  v1673,
  v1674,
  v1675,
  v1676,
  v1677,
  v1678,
  v1679,
  v1680,
  v1681,
  v1682,
  v1683,
  v1684,
  v1685,
  v1686,
  v1687,
  v1688,
  v1689,
  v1690,
  v1691,
  v1692,
  v1693,
  v1694,
  v1695,
  v1696,
  v1697,
  v1698,
  v1699,
  v1700,
  v1701,
  v1702,
  v1703,
  v1704,
  v1705,
  v1706,
  v1707,
  v1708,
  v1709,
  \*clm_file_1_istate0 ,
  \*clm_file_1_istate1 ,
  v1710,
  v1711,
  v1712,
  v1713,
  v1714,
  v1715,
  v1716,
  v1717,
  v1718,
  v1719,
  v1720,
  v1721,
  v1722,
  v1723,
  v1724,
  v1725,
  v1726,
  v1727,
  v1728,
  v1729,
  v1730,
  v1731,
  v1732,
  v1733,
  v1734,
  v1735,
  v1736,
  v1737,
  v1738,
  v1739,
  v1740,
  v1741,
  v1742,
  v1743,
  v1744,
  v1745,
  v1746,
  v1747,
  v1748,
  v1749,
  v1750,
  v1751,
  v1752,
  v1753,
  v1754,
  v1755,
  v1756,
  v1757,
  v1758,
  v1759,
  v1760,
  v1761,
  v1762,
  v1763,
  v1764,
  v1765,
  v1766,
  v1767,
  v1768,
  v1769,
  v1770,
  v1771,
  v1772,
  v1773,
  v1774,
  v1775,
  v1776,
  v1777,
  v1778,
  v1779,
  v1780,
  v1781,
  v1782,
  v1783,
  v1784,
  v1785,
  v1786,
  v1787,
  v1788,
  v1789,
  v1790,
  v1791,
  v1792,
  v1793,
  v1794,
  v1795,
  v1796,
  v1797,
  v1798,
  v1799,
  v1800,
  v1801,
  v1802,
  v1803,
  v1804,
  v1805,
  v1806,
  v1807,
  v1808,
  v1809,
  v1810,
  v1811,
  v1812,
  v1813,
  v1814,
  v1815,
  v1816,
  v1817,
  v1818,
  v1819,
  v1820,
  v1821,
  v1822,
  v1823,
  v1824,
  v1825,
  v1826,
  v1827,
  v1828,
  v1829,
  v1830,
  v1831,
  v1832,
  v1833,
  v1834,
  v1835,
  v1836,
  v1837,
  v1838,
  v1839,
  v1840,
  v1841,
  v1842,
  v1843,
  v1844,
  v1845,
  v1846,
  v1847,
  v1848,
  v1849,
  v1850,
  v1851,
  v1852,
  v1853,
  v1854,
  v1855,
  v1856,
  v1857,
  v1858,
  v1859,
  v1860,
  v1861,
  v1862,
  v1863,
  v1864,
  v1865,
  v1866,
  v1867,
  v1868,
  v1869,
  v1870,
  v1871,
  v1872,
  v1873,
  v1874,
  v1875,
  v1876,
  v1877,
  v1878,
  v1879,
  v1880,
  v1881,
  v1882,
  v1883,
  v1884,
  v1885,
  v1886,
  v1887,
  v1888,
  v1889,
  v1890,
  v1891,
  v1892,
  v1893,
  v1894,
  v1895,
  v1896,
  v1897,
  v1898,
  v1899,
  v1900,
  v1901,
  v1902,
  v1903,
  v1904,
  v1905,
  v1906,
  v1907,
  v1908,
  v1909,
  v1910,
  v1911,
  v1912,
  v1913,
  v1914,
  v1915,
  v1916,
  v1917,
  v1918,
  v1919,
  v1920,
  v1921,
  v1922,
  v1923,
  v1924,
  v1925,
  v1926,
  v1927,
  v1928,
  v1929,
  v1930,
  v1931,
  v1932,
  v1933,
  v1934,
  v1935,
  v1936,
  v1937,
  v1938,
  v1939,
  v1940,
  v1941,
  v1942,
  v1943,
  v1944,
  v1945,
  v1946,
  v1947,
  v1948,
  v1949,
  v1950,
  v1951,
  v1952,
  v1953,
  v1954,
  v1955,
  v1956,
  v1957,
  v1958,
  v1959,
  v1960,
  v1961,
  v1962,
  v1963,
  v1964,
  v1965,
  v1966,
  v1967,
  v1968,
  v1969,
  v1970,
  v1971,
  v1972,
  v1973,
  v1974,
  v1975,
  v1976,
  v1977,
  v1978,
  v1979,
  v1980,
  v1981,
  v1982,
  v1983,
  v1984,
  v1985,
  v1986,
  v1987,
  v1988,
  v1989,
  v1990,
  v1991,
  v1992,
  v1993,
  v1994,
  v1995,
  v1996,
  v1997,
  v1998,
  v1999,
  v2000,
  v2001,
  v2002,
  v2003,
  v2004,
  v2005,
  v2006,
  v2007,
  v2008,
  v2009,
  v2010,
  v2011,
  v2012,
  v2013,
  v2014,
  v2015,
  v2016,
  v2017,
  v2018,
  v2019,
  v2020,
  v2021,
  v2022,
  v2023,
  v2024,
  v2025,
  v2026,
  v2027,
  v2028,
  v2029,
  v2030,
  v2031,
  v2032,
  v2033,
  v2034,
  v2035,
  v2036,
  v2037,
  v2038,
  v2039,
  v2040,
  v2041,
  v2042,
  v2043,
  v2044,
  v2045,
  v2046,
  v2047,
  v2048,
  v2049,
  v2050,
  v2051,
  v2052,
  v2053,
  v2054,
  v2055,
  v2056,
  v2057,
  v2058,
  v2059,
  v2060,
  v2061,
  v2062,
  v2063,
  v2064,
  v2065,
  v2066,
  v2067,
  v2068,
  v2069,
  v2070,
  v2071,
  v2072,
  v2073,
  v2074,
  v2075,
  v2076,
  v2077,
  v2078,
  v2079,
  v2080,
  v2081,
  v2082,
  v2083,
  v2084,
  v2085,
  v2086,
  v2087,
  v2088,
  v2089,
  v2090,
  v2091,
  v2092,
  v2093,
  v2094,
  v2095,
  v2096,
  v2097,
  v2098,
  v2099,
  v2100,
  v2101,
  v2102,
  v2103,
  v2104,
  v2105,
  v2106,
  v2107,
  v2108,
  v2109,
  v2110,
  v2111,
  v2112,
  v2113,
  v2114,
  v2115,
  v2116,
  v2117,
  v2118,
  v2119,
  v2120,
  v2121,
  v2122,
  v2123,
  v2124,
  v2125,
  v2126,
  v2127,
  v2128,
  v2129,
  v2130,
  v2131,
  v2132,
  v2133,
  v2134,
  v2135,
  v2136,
  v2137,
  v2138,
  v2139,
  v2140,
  v2141,
  v2142,
  v2143,
  v2144,
  v2145,
  v2146,
  v2147,
  v2148,
  v2149,
  v2150,
  v2151,
  v2152,
  v2153,
  v2154,
  v2155,
  v2156,
  v2157,
  v2158,
  v2159,
  v2160,
  v2161,
  v2162,
  v2163,
  v2164,
  v2165,
  v2166,
  v2167,
  v2168,
  v2169,
  v2170,
  v2171,
  v2172,
  v2173,
  v2174,
  v2175,
  v2176,
  v2177,
  v2178,
  v2179,
  v2180,
  v2181,
  v2182,
  v2183,
  v2184,
  v2185,
  v2186,
  v2187,
  v2188,
  v2189,
  v2190,
  v2191,
  v2192,
  v2193,
  v2194,
  v2195,
  v2196,
  v2197,
  v2198,
  v2199,
  v2200,
  v2201,
  v2202,
  v2203,
  v2204,
  v2205,
  v2206,
  v2207,
  v2208,
  v2209,
  v2210,
  v2211,
  v2212,
  v2213,
  v2214,
  v2215,
  v2216,
  v2217,
  v2218,
  v2219,
  v2220,
  v2221,
  v2222,
  v2223,
  v2224,
  v2225,
  v2226,
  v2227,
  v2228,
  v2229,
  v2230,
  v2231,
  v2232,
  v2233,
  v2234,
  v2235,
  v2236,
  v2237,
  v2238,
  v2239,
  v2240,
  v2241,
  v2242,
  v2243,
  v2244,
  v2245,
  v2246,
  v2247,
  v2248,
  v2249,
  v2250,
  v2251,
  v2252,
  v2253,
  v2254,
  v2255,
  v2256,
  v2257,
  v2258,
  v2259,
  v2260,
  v2261,
  v2262,
  v2263,
  v2264,
  v2265,
  v2266,
  v2267,
  v2268,
  v2269,
  v2270,
  v2271,
  v2272,
  v2273,
  v2274,
  v2275,
  v2276,
  v2277,
  v2278,
  v2279,
  v2280,
  v2281,
  v2282,
  v2283,
  v2284,
  v2285,
  v2286,
  v2287,
  v2288,
  v2289,
  v2290,
  v2291,
  v2292,
  v2293,
  v2294,
  v2295,
  v2296,
  v2297,
  v2298,
  v2299,
  v2300,
  v2301,
  v2302,
  v2303,
  v2304,
  v2305,
  v2306,
  v2307,
  v2308,
  v2309,
  v2310,
  v2311,
  v2312,
  v2313,
  v2314,
  v2315,
  v2316,
  v2317,
  v2318,
  v2319,
  v2320,
  v2321,
  v2322,
  v2323,
  v2324,
  v2325,
  v2326,
  v2327,
  v2328,
  v2329,
  v2330,
  v2331,
  v2332,
  v2333,
  v2334,
  v2335,
  v2336,
  v2337,
  v2338,
  v2339,
  v2340,
  v2341,
  v2342,
  v2343,
  v2344,
  v2345,
  v2346,
  v2347,
  v2348,
  v2349,
  v2350,
  v2351,
  v2352,
  v2353,
  v2354,
  v2355,
  v2356,
  v2357,
  v2358,
  v2359,
  v2360,
  v2361,
  v2362,
  v2363,
  v2364,
  v2365,
  v2366,
  v2367,
  v2368,
  v2369,
  v2370,
  v2371,
  v2372,
  v2373,
  v2374,
  v2375,
  v2376,
  v2377,
  v2378,
  v2379,
  v2380,
  v2381,
  v2382,
  v2383,
  v2384,
  v2385,
  v2386,
  v2387,
  v2388,
  v2389,
  v2390,
  v2391,
  v2392,
  v2393,
  v2394,
  v2395,
  v2396,
  v2397,
  v2398,
  v2399,
  v2400,
  v2401,
  v2402,
  v2403,
  v2404,
  v2405,
  v2406,
  v2407,
  v2408,
  v2409,
  v2410,
  v2411,
  v2412,
  v2413,
  v2414,
  v2415,
  v2416,
  v2417,
  v2418,
  v2419,
  v2420,
  v2421,
  v2422,
  v2423,
  v2424,
  v2425,
  v2426,
  v2427,
  v2428,
  v2429,
  v2430,
  v2431,
  v2432,
  v2433,
  v2434,
  v2435,
  v2436,
  v2437,
  v2438,
  v2439,
  v2440,
  v2441,
  v2442,
  v2443,
  v2444,
  v2445,
  v2446,
  v2447,
  v2448,
  v2449,
  v2450,
  v2451,
  v2452,
  v2453,
  v2454,
  v2455,
  v2456,
  v2457,
  v2458,
  v2459,
  v2460,
  v2461,
  v2462,
  v2463,
  v2464,
  v2465,
  v2466,
  v2467,
  v2468,
  v2469,
  v2470,
  v2471,
  v2472,
  v2473,
  v2474,
  v2475,
  v2476,
  v2477,
  v2478,
  v2479,
  v2480,
  v2481,
  v2482,
  v2483,
  v2484,
  v2485,
  v2486,
  v2487,
  v2488,
  v2489,
  v2490,
  v2491,
  v2492,
  v2493,
  v2494,
  v2495,
  v2496,
  v2497,
  v2498,
  v2499,
  v2500,
  v2501,
  v2502,
  v2503,
  v2504,
  v2505,
  v2506,
  v2507,
  v2508,
  v2509,
  v2510,
  v2511,
  v2512,
  v2513,
  v2514,
  v2515,
  v2516,
  v2517,
  v2518,
  v2519,
  v2520,
  v2521,
  v2522,
  v2523,
  v2524,
  v2525,
  v2526,
  v2527,
  v2528,
  v2529,
  v2530,
  v2531,
  v2532,
  v2533,
  v2534,
  v2535,
  v2536,
  v2537,
  v2538,
  v2539,
  v2540,
  v2541,
  v2542,
  v2543,
  v2544,
  v2545,
  v2546,
  v2547,
  v2548,
  v2549,
  v2550,
  v2551,
  v2552,
  v2553,
  v2554,
  v2555,
  v2556,
  v2557,
  v2558,
  v2559,
  v2560,
  v2561,
  v2562,
  v2563,
  v2564,
  v2565,
  v2566,
  v2567,
  v2568,
  v2569,
  v2570,
  v2571,
  v2572,
  v2573,
  v2574,
  v2575,
  v2576,
  v2577,
  v2578,
  v2579,
  v2580,
  v2581,
  v2582,
  v2583,
  v2584,
  v2585,
  v2586,
  v2587,
  v2588,
  v2589,
  v2590,
  v2591,
  v2592,
  v2593,
  v2594,
  v2595,
  v2596,
  v2597,
  v2598,
  v2599,
  v2600,
  v2601,
  v2602,
  v2603,
  v2604,
  v2605,
  v2606,
  v2607,
  v2608,
  v2609,
  v2610,
  v2611,
  v2612,
  v2613,
  v2614,
  v2615,
  v2616,
  v2617,
  v2618,
  v2619,
  v2620,
  v2621,
  v2622,
  v2623,
  v2624,
  v2625,
  v2626,
  v2627,
  v2628,
  v2629,
  v2630,
  v2631,
  v2632,
  v2633,
  v2634,
  v2635,
  v2636,
  v2637,
  v2638,
  v2639,
  v2640,
  v2641,
  v2642,
  v2643,
  v2644,
  v2645,
  v2646,
  v2647,
  v2648,
  v2649,
  v2650,
  v2651,
  v2652,
  v2653,
  v2654,
  v2655,
  v2656,
  v2657,
  v2658,
  v2659,
  v2660,
  v2661,
  v2662,
  v2663,
  v2664,
  v2665,
  v2666,
  v2667,
  v2668,
  v2669,
  v2670,
  v2671,
  v2672,
  v2673,
  v2674,
  v2675,
  v2676,
  v2677,
  v2678,
  v2679,
  v2680,
  v2681,
  v2682,
  v2683,
  v2684,
  v2685,
  v2686,
  v2687,
  v2688,
  v2689,
  v2690,
  v2691,
  v2692,
  v2693,
  v2694,
  v2695,
  v2696,
  v2697,
  v2698,
  v2699,
  v2700,
  v2701,
  v2702,
  v2703,
  v2704,
  v2705,
  v2706,
  v2707,
  v2708,
  v2709,
  v2710,
  v2711,
  v2712,
  v2713,
  v2714,
  v2715,
  v2716,
  v2717,
  v2718,
  v2719,
  v2720,
  v2721,
  v2722,
  v2723,
  v2724,
  v2725,
  v2726,
  v2727,
  v2728,
  v2729,
  v2730,
  v2731,
  v2732,
  v2733,
  v2734,
  v2735,
  v2736,
  v2737,
  v2738,
  v2739,
  v2740,
  v2741,
  v2742,
  v2743,
  v2744,
  v2745,
  v2746,
  v2747,
  v2748,
  v2749,
  v2750,
  v2751,
  v2752,
  v2753,
  v2754,
  v2755,
  v2756,
  v2757,
  v2758,
  v2759,
  v2760,
  v2761,
  v2762,
  v2763,
  v2764,
  v2765,
  v2766,
  v2767,
  v2768,
  v2769,
  v2770,
  v2771,
  v2772,
  v2773,
  v2774,
  v2775,
  v2776,
  v2777,
  v2778,
  v2779,
  v2780,
  v2781,
  v2782,
  v2783,
  v2784,
  v2785,
  v2786,
  v2787,
  v2788,
  v2789,
  v2790,
  v2791,
  v2792,
  v2793,
  v2794,
  v2795,
  v2796,
  v2797,
  v2798,
  v2799,
  v2800,
  v2801,
  v2802,
  v2803,
  v2804,
  v2805,
  v2806,
  v2807,
  v2808,
  v2809,
  v2810,
  v2811,
  v2812,
  v2813,
  v2814,
  v2815,
  v2816,
  v2817,
  v2818,
  v2819,
  v2820,
  v2821,
  v2822,
  v2823,
  v2824,
  v2825,
  v2826,
  v2827,
  v2828,
  v2829,
  v2830,
  v2831,
  v2832,
  v2833,
  v2834,
  v2835,
  v2836,
  v2837,
  v2838,
  v2839,
  v2840,
  v2841,
  v2842,
  v2843,
  v2844,
  v2845,
  v2846,
  v2847,
  v2848,
  v2849,
  v2850,
  v2851,
  v2852,
  v2853,
  v2854,
  v2855,
  v2856,
  v2857,
  v2858,
  v2859,
  v2860,
  v2861,
  v2862,
  v2863,
  v2864,
  v2865,
  v2866,
  v2867,
  v2868,
  v2869,
  v2870,
  v2871,
  v2872,
  v2873,
  v2874,
  v2875,
  v2876,
  v2877,
  v2878,
  v2879,
  v2880,
  v2881,
  v2882,
  v2883,
  v2884,
  v2885,
  v2886,
  v2887,
  v2888,
  v2889,
  v2890,
  v2891,
  v2892,
  v2893,
  v2894,
  v2895,
  v2896,
  v2897,
  v2898,
  v2899,
  v2900,
  v2901,
  v2902,
  v2903,
  v2904,
  v2905,
  v2906,
  v2907,
  v2908,
  v2909,
  v2910,
  v2911,
  v2912,
  v2913,
  v2914,
  v2915,
  v2916,
  v2917,
  v2918,
  v2919,
  v2920,
  v2921,
  v2922,
  v2923,
  v2924,
  v2925,
  v2926,
  v2927,
  v2928,
  v2929,
  v2930,
  v2931,
  v2932,
  v2933,
  v2934,
  v2935,
  v2936,
  v2937,
  v2938,
  v2939,
  v2940,
  v2941,
  v2942,
  v2943,
  v2944,
  v2945,
  v2946,
  v2947,
  v2948,
  v2949,
  v2950,
  v2951,
  v2952,
  v2953,
  v2954,
  v2955,
  v2956,
  v2957,
  v2958,
  v2959,
  v2960,
  v2961,
  v2962,
  v2963,
  v2964,
  v2965,
  v2966,
  v2967,
  v2968,
  v2969,
  v2970,
  v2971,
  v2972,
  v2973,
  v2974,
  v2975,
  v2976,
  v2977,
  v2978,
  v2979,
  v2980,
  v2981,
  v2982,
  v2983,
  v2984,
  v2985,
  v2986,
  v2987,
  v2988,
  v2989,
  v2990,
  v2991,
  v2992,
  v2993,
  v2994,
  v2995,
  v2996,
  v2997,
  v2998,
  v2999,
  v3000,
  v3001,
  v3002,
  v3003,
  v3004,
  v3005,
  v3006,
  v3007,
  v3008,
  v3009,
  v3010,
  v3011,
  v3012,
  v3013,
  v3014,
  v3015,
  v3016,
  v3017,
  v3018,
  v3019,
  v3020,
  v3021,
  v3022,
  v3023,
  v3024,
  v3025,
  v3026,
  v3027,
  v3028,
  v3029,
  v3030,
  v3031,
  v3032,
  v3033,
  v3034,
  v3035,
  v3036,
  v3037,
  v3038,
  v3039,
  v3040,
  v3041,
  v3042,
  v3043,
  v3044,
  v3045,
  v3046,
  v3047,
  v3048,
  v3049,
  v3050,
  v3051,
  v3052,
  v3053,
  v3054,
  v3055,
  v3056,
  v3057,
  v3058,
  v3059,
  v3060,
  v3061,
  v3062,
  v3063,
  v3064,
  v3065,
  v3066,
  v3067,
  v3068,
  v3069,
  v3070,
  v3071,
  v3072,
  v3073,
  v3074,
  v3075,
  v3076,
  v3077,
  v3078,
  v3079,
  v3080,
  v3081,
  v3082,
  v3083,
  v3084,
  v3085,
  v3086,
  v3087,
  v3088,
  v3089,
  v3090,
  v3091,
  v3092,
  v3093,
  v3094,
  v3095,
  v3096,
  v3097,
  v3098,
  v3099,
  v3100,
  v3101,
  v3102,
  v3103,
  v3104,
  v3105,
  v3106,
  v3107,
  v3108,
  v3109,
  v3110,
  v3111,
  v3112,
  v3113,
  v3114,
  v3115,
  v3116,
  v3117,
  v3118,
  v3119,
  v3120,
  v3121,
  v3122,
  v3123,
  v3124,
  v3125,
  v3126,
  v3127,
  v3128,
  v3129,
  v3130,
  v3131,
  v3132,
  v3133,
  v3134,
  v3135,
  v3136,
  v3137,
  v3138,
  v3139,
  v3140,
  v3141,
  v3142,
  v3143,
  v3144,
  v3145,
  v3146,
  v3147,
  v3148,
  v3149,
  v3150,
  v3151,
  v3152,
  v3153,
  v3154,
  v3155,
  v3156,
  v3157,
  v3158,
  v3159,
  v3160,
  v3161,
  v3162,
  v3163,
  v3164,
  v3165,
  v3166,
  v3167,
  v3168,
  v3169,
  v3170,
  v3171,
  v3172,
  v3173,
  v3174,
  v3175,
  v3176,
  v3177,
  v3178,
  v3179,
  v3180,
  v3181,
  v3182,
  v3183,
  v3184,
  v3185,
  v3186,
  v3187,
  v3188,
  v3189,
  v3190,
  v3191,
  v3192,
  v3193,
  v3194,
  v3195,
  v3196,
  v3197,
  v3198,
  v3199,
  v3200,
  v3201,
  v3202,
  v3203,
  v3204,
  v3205,
  v3206,
  v3207,
  v3208,
  v3209,
  v3210,
  v3211,
  v3212,
  v3213,
  v3214,
  v3215,
  v3216,
  v3217,
  v3218,
  v3219,
  v3220,
  v3221,
  v3222,
  v3223,
  v3224,
  v3225,
  v3226,
  v3227,
  v3228,
  v3229,
  v3230,
  v3231,
  v3232,
  v3233,
  v3234,
  v3235,
  v3236,
  v3237,
  v3238,
  v3239,
  v3240,
  v3241,
  v3242,
  v3243,
  v3244,
  v3245,
  v3246,
  v3247,
  v3248,
  v3249,
  v3250,
  v3251,
  v3252,
  v3253,
  v3254,
  v3255,
  v3256,
  v3257,
  v3258,
  v3259,
  v3260,
  v3261,
  v3262,
  v3263,
  v3264,
  v3265,
  v3266,
  v3267,
  v3268,
  v3269,
  v3270,
  v3271,
  v3272,
  v3273,
  v3274,
  v3275,
  v3276,
  v3277,
  v3278,
  v3279,
  v3280,
  v3281,
  v3282,
  v3283,
  v3284,
  v3285,
  v3286,
  v3287,
  v3288,
  v3289,
  v3290,
  v3291,
  v3292,
  v3293,
  v3294,
  v3295,
  v3296,
  v3297,
  v3298,
  v3299,
  v3300,
  v3301,
  v3302,
  v3303,
  v3304,
  v3305,
  v3306,
  v3307,
  v3308,
  v3309,
  v3310,
  v3311,
  v3312,
  v3313,
  v3314,
  v3315,
  v3316,
  v3317,
  v3318,
  v3319,
  v3320,
  v3321,
  v3322,
  v3323,
  v3324,
  v3325,
  v3326,
  v3327,
  v3328,
  v3329,
  v3330,
  v3331,
  v3332,
  v3333,
  v3334,
  v3335,
  v3336,
  v3337,
  v3338,
  v3339,
  v3340,
  v3341,
  v3342,
  v3343,
  v3344,
  v3345,
  v3346,
  v3347,
  v3348,
  v3349,
  v3350,
  v3351,
  v3352,
  v3353,
  v3354,
  v3355,
  v3356,
  v3357,
  v3358,
  v3359,
  v3360,
  v3361,
  v3362,
  v3363,
  v3364,
  v3365,
  v3366,
  v3367,
  v3368,
  v3369,
  v3370,
  v3371,
  v3372,
  v3373,
  v3374,
  v3375,
  v3376,
  v3377,
  v3378,
  v3379,
  v3380,
  v3381,
  v3382,
  v3383,
  v3384,
  v3385,
  v3386,
  v3387,
  v3388,
  v3389,
  v3390,
  v3391,
  v3392,
  v3393,
  v3394,
  v3395,
  v3396,
  v3397,
  v3398,
  v3399,
  v3400,
  v3401,
  v3402,
  v3403,
  v3404,
  v3405,
  v3406,
  v3407,
  v3408,
  v3409,
  v3410,
  v3411,
  v3412,
  v3413,
  v3414,
  v3415,
  v3416,
  v3417,
  v3418,
  v3419,
  v3420,
  v3421,
  v3422,
  v3423,
  v3424,
  v3425,
  v3426,
  v3427,
  v3428,
  v3429,
  v3430,
  v3431,
  v3432,
  v3433,
  v3434,
  v3435,
  v3436,
  v3437,
  v3438,
  v3439,
  v3440,
  v3441,
  v3442,
  v3443,
  v3444,
  v3445,
  v3446,
  v3447,
  v3448,
  v3449,
  v3450,
  v3451,
  v3452,
  v3453,
  v3454,
  v3455,
  v3456,
  v3457,
  v3458,
  v3459,
  v3460,
  v3461,
  v3462,
  v3463,
  v3464,
  v3465,
  v3466,
  v3467,
  v3468,
  v3469,
  v3470,
  v3471,
  v3472,
  v3473,
  v3474,
  v3475,
  v3476,
  v3477,
  v3478,
  v3479,
  v3480,
  v3481,
  v3482,
  v3483,
  v3484,
  v3485,
  v3486,
  v3487,
  v3488,
  v3489,
  v3490,
  v3491,
  v3492,
  v3493,
  v3494,
  v3495,
  v3496,
  v3497,
  v3498,
  v3499,
  v3500,
  v3501,
  v3502,
  v3503,
  v3504,
  v3505,
  v3506,
  v3507,
  v3508,
  v3509,
  v3510,
  v3511,
  v3512,
  v3513,
  v3514,
  v3515,
  v3516,
  v3517,
  v3518,
  v3519,
  v3520,
  v3521,
  v3522,
  v3523,
  v3524,
  v3525,
  v3526,
  v3527,
  v3528,
  v3529,
  v3530,
  v3531,
  v3532,
  v3533,
  v3534,
  v3535,
  v3536,
  v3537,
  v3538,
  v3539,
  v3540,
  v3541,
  v3542,
  v3543,
  v3544,
  v3545,
  v3546,
  v3547,
  v3548,
  v3549,
  v3550,
  v3551,
  v3552,
  v3553,
  v3554,
  v3555,
  v3556,
  v3557,
  v3558,
  v3559,
  v3560,
  v3561,
  v3562,
  v3563,
  v3564,
  v3565,
  v3566,
  v3567,
  v3568,
  v3569,
  v3570,
  v3571,
  v3572,
  v3573,
  v3574,
  v3575,
  v3576,
  v3577,
  v3578,
  v3579,
  v3580,
  v3581,
  v3582,
  v3583,
  v3584,
  v3585,
  v3586,
  v3587,
  v3588,
  v3589,
  v3590,
  v3591,
  v3592,
  v3593,
  v3594,
  v3595,
  v3596,
  v3597,
  v3598,
  v3599,
  v3600,
  v3601,
  v3602,
  v3603,
  v3604,
  v3605,
  v3606,
  v3607,
  v3608,
  v3609,
  v3610,
  v3611,
  v3612,
  v3613,
  v3614,
  v3615,
  v3616,
  v3617,
  v3618,
  v3619,
  v3620,
  v3621,
  v3622,
  v3623,
  v3624,
  v3625,
  v3626,
  v3627,
  v3628,
  v3629,
  v3630,
  v3631,
  v3632,
  v3633,
  v3634,
  v3635,
  v3636,
  v3637,
  v3638,
  v3639,
  v3640,
  v3641,
  v3642,
  v3643,
  v3644,
  v3645,
  v3646,
  v3647,
  v3648,
  v3649,
  v3650,
  v3651,
  v3652,
  v3653,
  v3654,
  v3655,
  v3656,
  v3657,
  v3658,
  v3659,
  v3660,
  v3661,
  v3662,
  v3663,
  v3664,
  v3665,
  v3666,
  v3667,
  v3668,
  v3669,
  v3670,
  v3671,
  v3672,
  v3673,
  v3674,
  v3675,
  v3676,
  v3677,
  v3678,
  v3679,
  v3680,
  v3681,
  v3682,
  v3683,
  v3684,
  v3685,
  v3686,
  v3687,
  v3688,
  v3689,
  v3690,
  v3691,
  v3692,
  v3693,
  v3694,
  v3695,
  v3696,
  v3697,
  v3698,
  v3699,
  v3700,
  v3701,
  v3702,
  v3703,
  v3704,
  v3705,
  v3706,
  v3707,
  v3708,
  v3709,
  v3710,
  v3711,
  v3712,
  v3713,
  v3714,
  v3715,
  v3716,
  v3717,
  v3718,
  v3719,
  v3720,
  v3721,
  v3722,
  v3723,
  v3724,
  v3725,
  v3726,
  v3727,
  v3728,
  v3729,
  v3730,
  v3731,
  v3732,
  v3733,
  v3734,
  v3735,
  v3736,
  v3737,
  v3738,
  v3739,
  v3740,
  v3741,
  v3742,
  v3743,
  v3744,
  v3745,
  v3746,
  v3747,
  v3748,
  v3749,
  v3750,
  v3751,
  v3752,
  v3753,
  v3754,
  v3755,
  v3756,
  v3757,
  v3758,
  v3759,
  v3760,
  v3761,
  v3762,
  v3763,
  v3764,
  v3765,
  v3766,
  v3767,
  v3768,
  v3769,
  v10000,
  v10001,
  v10002,
  v3770,
  v10003,
  v3771,
  v10004,
  v3772,
  v10005,
  v3773,
  v10006,
  v3774,
  v10007,
  v3775,
  v10008,
  v3776,
  v10009,
  v3777,
  v3778,
  v3779,
  v10010,
  v10011,
  v10012,
  v3780,
  v10013,
  v3781,
  v10014,
  v3782,
  v10015,
  v3783,
  v10016,
  v3784,
  v10017,
  v3785,
  v10018,
  v3786,
  v10019,
  v3787,
  v3788,
  v3789,
  v10020,
  v10021,
  v10022,
  v3790,
  v10023,
  v3791,
  v10024,
  v3792,
  v10025,
  v3793,
  v10026,
  v3794,
  v10027,
  v3795,
  v10028,
  v3796,
  v10029,
  v3797,
  v3798,
  v3799,
  v10030,
  v10031,
  v10032,
  v10033,
  v10034,
  v10035,
  v10036,
  v10037,
  v10038,
  v10039,
  v10040,
  v10041,
  v10042,
  v10043,
  v10044,
  v10045,
  v10046,
  v10047,
  v10048,
  v10049,
  v10050,
  v10051,
  v10052,
  v10053,
  v10054,
  v10055,
  v10056,
  v10057,
  v10058,
  v10059,
  v10060,
  v10061,
  v10062,
  v10063,
  v10064,
  v10065,
  v10066,
  v10067,
  v10068,
  v10069,
  v10070,
  v10071,
  v10072,
  v10073,
  v10074,
  v10075,
  v10076,
  v10077,
  v10078,
  v10079,
  v10080,
  v10081,
  v10082,
  v10083,
  v10084,
  v10085,
  v10086,
  v10087,
  v10088,
  v10089,
  v10090,
  v10091,
  v10092,
  v3800,
  v10093,
  v3801,
  v10094,
  v3802,
  v10095,
  v3803,
  v10096,
  v3804,
  v10097,
  v3805,
  v10098,
  v3806,
  v10099,
  v3807,
  v3808,
  v3809,
  v3810,
  v3811,
  v3812,
  v3813,
  v3814,
  v3815,
  v3816,
  v3817,
  v3818,
  v3819,
  v3820,
  v3821,
  v3822,
  v3823,
  v3824,
  v3825,
  v3826,
  v3827,
  v3828,
  v3829,
  v3830,
  v3831,
  v3832,
  v3833,
  v3834,
  v3835,
  v3836,
  v3837,
  v3838,
  v3839,
  v3840,
  v3841,
  v3842,
  v3843,
  v3844,
  v3845,
  v3846,
  v3847,
  v3848,
  v3849,
  v3850,
  v3851,
  v3852,
  v3853,
  v3854,
  v3855,
  v3856,
  v3857,
  v3858,
  v3859,
  v3860,
  v3861,
  v3862,
  v3863,
  v3864,
  v3865,
  v3866,
  v3867,
  v3868,
  v3869,
  v10100,
  v10101,
  v10102,
  v3870,
  v10103,
  v3871,
  v10104,
  v3872,
  v10105,
  v3873,
  v10106,
  v3874,
  v10107,
  v3875,
  v10108,
  v3876,
  v10109,
  v3877,
  v3878,
  v3879,
  v10110,
  v10111,
  v10112,
  v3880,
  v10113,
  v3881,
  v10114,
  v3882,
  v10115,
  v3883,
  v10116,
  v3884,
  v10117,
  v3885,
  v10118,
  v3886,
  v10119,
  v3887,
  v3888,
  v3889,
  v10120,
  v10121,
  v10122,
  v3890,
  v10123,
  v3891,
  v10124,
  v3892,
  v10125,
  v3893,
  v10126,
  v3894,
  v10127,
  v3895,
  v10128,
  v3896,
  v10129,
  v3897,
  v3898,
  v3899,
  v10130,
  v10131,
  v10132,
  v10133,
  v10134,
  v10135,
  v10136,
  v10137,
  v10138,
  v10139,
  v10140,
  v10141,
  v10142,
  v10143,
  v10144,
  v10145,
  v10146,
  v10147,
  v10148,
  v10149,
  v10150,
  v10151,
  v10152,
  v10153,
  v10154,
  v10155,
  v10156,
  v10157,
  v10158,
  v10159,
  v10160,
  v10161,
  v10162,
  v10163,
  v10164,
  v10165,
  v10166,
  v10167,
  v10168,
  v10169,
  v10170,
  v10171,
  v10172,
  v10173,
  v10174,
  v10175,
  v10176,
  v10177,
  v10178,
  v10179,
  v10180,
  v10181,
  v10182,
  v10183,
  v10184,
  v10185,
  v10186,
  v10187,
  v10188,
  v10189,
  v10190,
  v10191,
  v10192,
  v3900,
  v10193,
  v3901,
  v10194,
  v3902,
  v10195,
  v3903,
  v10196,
  v3904,
  v10197,
  v3905,
  v10198,
  v3906,
  v10199,
  v3907,
  v3908,
  v3909,
  v3910,
  v3911,
  v3912,
  v3913,
  v3914,
  v3915,
  v3916,
  v3917,
  v3918,
  v3919,
  v3920,
  v3921,
  v3922,
  v3923,
  v3924,
  v3925,
  v3926,
  v3927,
  v3928,
  v3929,
  v3930,
  v3931,
  v3932,
  v3933,
  v3934,
  v3935,
  v3936,
  v3937,
  v3938,
  v3939,
  v3940,
  v3941,
  v3942,
  v3943,
  v3944,
  v3945,
  v3946,
  v3947,
  v3948,
  v3949,
  v3950,
  v3951,
  v3952,
  v3953,
  v3954,
  v3955,
  v3956,
  v3957,
  v3958,
  v3959,
  v3960,
  v3961,
  v3962,
  v3963,
  v3964,
  v3965,
  v3966,
  v3967,
  v3968,
  v3969,
  v10200,
  v10201,
  v10202,
  v3970,
  v10203,
  v3971,
  v10204,
  v3972,
  v10205,
  v3973,
  v10206,
  v3974,
  v10207,
  v3975,
  v10208,
  v3976,
  v10209,
  v3977,
  v3978,
  v3979,
  v10210,
  v10211,
  v10212,
  v3980,
  v10213,
  v3981,
  v10214,
  v3982,
  v10215,
  v3983,
  v10216,
  v3984,
  v10217,
  v3985,
  v10218,
  v3986,
  v10219,
  v3987,
  v3988,
  v3989,
  v10220,
  v10221,
  v10222,
  v3990,
  v10223,
  v3991,
  v10224,
  v3992,
  v10225,
  v3993,
  v10226,
  v3994,
  v10227,
  v3995,
  v10228,
  v3996,
  v10229,
  v3997,
  v3998,
  v3999,
  v10230,
  v10231,
  v10232,
  v10233,
  v10234,
  v10235,
  v10236,
  v10237,
  v10238,
  v10239,
  v10240,
  v10241,
  v10242,
  v10243,
  v10244,
  v10245,
  v10246,
  v10247,
  v10248,
  v10249,
  v10250,
  v10251,
  v10252,
  v10253,
  v10254,
  v10255,
  v10256,
  v10257,
  v10258,
  v10259,
  v10260,
  v10261,
  v10262,
  v10263,
  v10264,
  v10265,
  v10266,
  v10267,
  v10268,
  v10269,
  v10270,
  v10271,
  v10272,
  v10273,
  v10274,
  v10275,
  v10276,
  v10277,
  v10278,
  v10279,
  v10280,
  v10281,
  v10282,
  v10283,
  v10284,
  v10285,
  v10286,
  v10287,
  v10288,
  v10289,
  v10290,
  v10291,
  v10292,
  v10293,
  v10294,
  v10295,
  v10296,
  v10297,
  v10298,
  v10299,
  v10300,
  v10301,
  v10302,
  v10303,
  v10304,
  v10305,
  v10306,
  v10307,
  v10308,
  v10309,
  v10310,
  v10311,
  v10312,
  v10313,
  v10314,
  v10315,
  v10316,
  v10317,
  v10318,
  v10319,
  v10320,
  v10321,
  v10322,
  v10323,
  v10324,
  v10325,
  v10326,
  v10327,
  v10328,
  v10329,
  v4000,
  v4001,
  v4002,
  v4003,
  v4004,
  v4005,
  v4006,
  v4007,
  v4008,
  v4009,
  v4010,
  v4011,
  v4012,
  v4013,
  v4014,
  v4015,
  v4016,
  v4017,
  v4018,
  v4019,
  v4020,
  v4021,
  v4022,
  v4023,
  v4024,
  v4025,
  v4026,
  v4027,
  v4028,
  v4029,
  v4030,
  v4031,
  v4032,
  v4033,
  v4034,
  v4035,
  v4036,
  v4037,
  v4038,
  v4039,
  v4040,
  v4041,
  v4042,
  v4043,
  v4044,
  v4045,
  v4046,
  v4047,
  v4048,
  v4049,
  v4050,
  v4051,
  v4052,
  v4053,
  v4054,
  v4055,
  v4056,
  v4057,
  \*clm_clk_ctl_time0 ,
  v4058,
  \*clm_clk_ctl_time1 ,
  v4059,
  v4060,
  v4061,
  v4062,
  v4063,
  v4064,
  v4065,
  v4066,
  v4067,
  v4068,
  v4069,
  v4070,
  v4071,
  v4072,
  v4073,
  v4074,
  v4075,
  v4076,
  v4077,
  v4078,
  v4079,
  v4080,
  v4081,
  v4082,
  v4083,
  v4084,
  v4085,
  v4086,
  v4087,
  v4088,
  v4089,
  v4090,
  v4091,
  v4092,
  v4093,
  v4094,
  v4095,
  v4096,
  v4097,
  v4098,
  v4099,
  v4100,
  v4101,
  v4102,
  v4103,
  v4104,
  v4105,
  v4106,
  v4107,
  v4108,
  v4109,
  v4110,
  v4111,
  v4112,
  v4113,
  v4114,
  v4115,
  v4116,
  v4117,
  v4118,
  v4119,
  v4120,
  v4121,
  v4122,
  v4123,
  v4124,
  v4125,
  v4126,
  v4127,
  v4128,
  v4129,
  v4130,
  v4131,
  v4132,
  v4133,
  v4134,
  v4135,
  v4136,
  v4137,
  v4138,
  v4139,
  v4140,
  v4141,
  v4142,
  v4143,
  v4144,
  v4145,
  v4146,
  v4147,
  v4148,
  v4149,
  v4150,
  v4151,
  v4152,
  v4153,
  v4154,
  v4155,
  v4156,
  v4157,
  v4158,
  v4159,
  v4160,
  v4161,
  v4162,
  v4163,
  v4164,
  v4165,
  v4166,
  v4167,
  v4168,
  v4169,
  v4170,
  v4171,
  v4172,
  v4173,
  v4174,
  v4175,
  v4176,
  v4177,
  v4178,
  v4179,
  v4180,
  v4181,
  v4182,
  v4183,
  v4184,
  v4185,
  v4186,
  v4187,
  v4188,
  v4189,
  v4190,
  v4191,
  v4192,
  v4193,
  v4194,
  v4195,
  v4196,
  v4197,
  v4198,
  v4199,
  v4200,
  v4201,
  v4202,
  v4203,
  v4204,
  v4205,
  v4206,
  v4207,
  v4208,
  v4209,
  v4210,
  v4211,
  v4212,
  v4213,
  v4214,
  v4215,
  v4216,
  v4217,
  v4218,
  v4219,
  v4220,
  v4221,
  v4222,
  v4223,
  v4224,
  v4225,
  v4226,
  v4227,
  v4228,
  v4229,
  v4230,
  v4231,
  v4232,
  v4233,
  v4234,
  v4235,
  v4236,
  v4237,
  v4238,
  v4239,
  v4240,
  v4241,
  v4242,
  v4243,
  v4244,
  v4245,
  v4246,
  v4247,
  v4248,
  v4249,
  v4250,
  v4251,
  v4252,
  v4253,
  v4254,
  v4255,
  v4256,
  v4257,
  v4258,
  v4259,
  v4260,
  v4261,
  v4262,
  v4263,
  v4264,
  v4265,
  v4266,
  v4267,
  v4268,
  v4269,
  v4270,
  v4271,
  v4272,
  v4273,
  v4274,
  v4275,
  v4276,
  v4277,
  v4278,
  v4279,
  v4280,
  v4281,
  v4282,
  v4283,
  v4284,
  v4285,
  v4286,
  v4287,
  v4288,
  v4289,
  v4290,
  v4291,
  v4292,
  v4293,
  v4294,
  v4295,
  v4296,
  v4297,
  v4298,
  v4299,
  v4300,
  v4301,
  v4302,
  v4303,
  v4304,
  v4305,
  v4306,
  v4307,
  v4308,
  v4309,
  v4310,
  v4311,
  v4312,
  v4313,
  v4314,
  v4315,
  v4316,
  v4317,
  v4318,
  v4319,
  v4320,
  v4321,
  v4322,
  v4323,
  v4324,
  v4325,
  v4326,
  v4327,
  v4328,
  v4329,
  v4330,
  v4331,
  v4332,
  v4333,
  v4334,
  v4335,
  v4336,
  v4337,
  v4338,
  v4339,
  v4340,
  v4341,
  v4342,
  v4343,
  v4344,
  v4345,
  v4346,
  v4347,
  v4348,
  v4349,
  v4350,
  v4351,
  v4352,
  v4353,
  v4354,
  v4355,
  v4356,
  v4357,
  v4358,
  v4359,
  v4360,
  v4361,
  v4362,
  v4363,
  v4364,
  v4365,
  v4366,
  v4367,
  v4368,
  v4369,
  v4370,
  v4371,
  v4372,
  v4373,
  v4374,
  v4375,
  v4376,
  v4377,
  v4378,
  v4379,
  v4380,
  v4381,
  v4382,
  v4383,
  v4384,
  v4385,
  v4386,
  v4387,
  v4388,
  v4389,
  v4390,
  v4391,
  v4392,
  v4393,
  v4394,
  v4395,
  v4396,
  v4397,
  v4398,
  v4399,
  v4400,
  v4401,
  v4402,
  v4403,
  v4404,
  v4405,
  v4406,
  v4407,
  v4408,
  v4409,
  v4410,
  v4411,
  v4412,
  v4413,
  v4414,
  v4415,
  v4416,
  v4417,
  v4418,
  v4419,
  v4420,
  v4421,
  v4422,
  v4423,
  v4424,
  v4425,
  v4426,
  v4427,
  v4428,
  v4429,
  v4430,
  v4431,
  v4432,
  v4433,
  v4434,
  v4435,
  v4436,
  v4437,
  v4438,
  v4439,
  v4440,
  v4441,
  v4442,
  v4443,
  v4444,
  v4445,
  v4446,
  v4447,
  v4448,
  v4449,
  v4450,
  v4451,
  v4452,
  v4453,
  v4454,
  v4455,
  v4456,
  v4457,
  v4458,
  v4459,
  v4460,
  v4461,
  v4462,
  v4463,
  v4464,
  v4465,
  v4466,
  v4467,
  v4468,
  v4469,
  v4470,
  v4471,
  v4472,
  v4473,
  v4474,
  v4475,
  v4476,
  v4477,
  v4478,
  v4479,
  v4480,
  v4481,
  v4482,
  v4483,
  v4484,
  v4485,
  v4486,
  v4487,
  v4488,
  v4489,
  v4490,
  v4491,
  v4492,
  v4493,
  v4494,
  v4495,
  v4496,
  v4497,
  v4498,
  v4499,
  v4500,
  v4501,
  v4502,
  v4503,
  v4504,
  v4505,
  v4506,
  v4507,
  v4508,
  v4509,
  v4510,
  v4511,
  v4512,
  v4513,
  v4514,
  v4515,
  v4516,
  v4517,
  v4518,
  v4519,
  v4520,
  v4521,
  v4522,
  v4523,
  v4524,
  v4525,
  v4526,
  v4527,
  v4528,
  v4529,
  v4530,
  v4531,
  v4532,
  v4533,
  v4534,
  v4535,
  v4536,
  v4537,
  v4538,
  v4539,
  v4540,
  v4541,
  v4542,
  v4543,
  v4544,
  v4545,
  v4546,
  v4547,
  v4548,
  v4549,
  v4550,
  v4551,
  v4552,
  v4553,
  v4554,
  v4555,
  v4556,
  v4557,
  v4558,
  v4559,
  v4560,
  v4561,
  v4562,
  v4563,
  v4564,
  v4565,
  v4566,
  v4567,
  v4568,
  v4569,
  v4570,
  v4571,
  v4572,
  v4573,
  v4574,
  v4575,
  v4576,
  v4577,
  v4578,
  v4579,
  v4580,
  v4581,
  v4582,
  v4583,
  v4584,
  v4585,
  v4586,
  v4587,
  v4588,
  v4589,
  v4590,
  v4591,
  v4592,
  v4593,
  v4594,
  v4595,
  v4596,
  v4597,
  v4598,
  v4599,
  v4600,
  v4601,
  v4602,
  v4603,
  v4604,
  v4605,
  v4606,
  v4607,
  v4608,
  v4609,
  v4610,
  v4611,
  v4612,
  v4613,
  v4614,
  v4615,
  v4616,
  v4617,
  v4618,
  v4619,
  v4620,
  v4621,
  v4622,
  v4623,
  v4624,
  v4625,
  v4626,
  v4627,
  v4628,
  v4629,
  v4630,
  v4631,
  v4632,
  v4633,
  v4634,
  v4635,
  v4636,
  v4637,
  v4638,
  v4639,
  v4640,
  v4641,
  v4642,
  v4643,
  v4644,
  v4645,
  v4646,
  v4647,
  v4648,
  v4649,
  v4650,
  v4651,
  v4652,
  v4653,
  v4654,
  v4655,
  v4656,
  v4657,
  v4658,
  v4659,
  v4660,
  v4661,
  v4662,
  v4663,
  v4664,
  v4665,
  v4666,
  v4667,
  v4668,
  v4669,
  v4670,
  v4671,
  v4672,
  v4673,
  v4674,
  v4675,
  v4676,
  v4677,
  v4678,
  v4679,
  v4680,
  v4681,
  v4682,
  v4683,
  v4684,
  v4685,
  v4686,
  v4687,
  v4688,
  v4689,
  v4690,
  v4691,
  v4692,
  v4693,
  v4694,
  v4695,
  v4696,
  v4697,
  v4698,
  v4699,
  v4700,
  v4701,
  v4702,
  v4703,
  v4704,
  v4705,
  v4706,
  v4707,
  v4708,
  v4709,
  v4710,
  v4711,
  v4712,
  v4713,
  v4714,
  v4715,
  v4716,
  v4717,
  v4718,
  v4719,
  v4720,
  v4721,
  v4722,
  v4723,
  v4724,
  v4725,
  v4726,
  v4727,
  v4728,
  v4729,
  v4730,
  v4731,
  v4732,
  v4733,
  v4734,
  v4735,
  v4736,
  v4737,
  v4738,
  v4739,
  v4740,
  v4741,
  v4742,
  v4743,
  v4744,
  v4745,
  v4746,
  v4747,
  v4748,
  v4749,
  v4750,
  v4751,
  v4752,
  v4753,
  v4754,
  v4755,
  v4756,
  v4757,
  v4758,
  v4759,
  v4760,
  v4761,
  v4762,
  v4763,
  v4764,
  v4765,
  v4766,
  v4767,
  v4768,
  v4769,
  v4770,
  v4771,
  v4772,
  v4773,
  v4774,
  v4775,
  v4776,
  v4777,
  v4778,
  v4779,
  v4780,
  v4781,
  v4782,
  v4783,
  v4784,
  v4785,
  v4786,
  v4787,
  v4788,
  v4789,
  v4790,
  v4791,
  v4792,
  v4793,
  v4794,
  v4795,
  v4796,
  v4797,
  v4798,
  v4799,
  v4800,
  v4801,
  v4802,
  v4803,
  v4804,
  v4805,
  v4806,
  v4807,
  v4808,
  v4809,
  v4810,
  v4811,
  v4812,
  v4813,
  v4814,
  v4815,
  v4816,
  v4817,
  v4818,
  v4819,
  v4820,
  v4821,
  v4822,
  v4823,
  v4824,
  v4825,
  v4826,
  v4827,
  v4828,
  v4829,
  v4830,
  v4831,
  v4832,
  v4833,
  v4834,
  v4835,
  v4836,
  v4837,
  v4838,
  v4839,
  v4840,
  v4841,
  v4842,
  v4843,
  v4844,
  v4845,
  v4846,
  v4847,
  v4848,
  v4849,
  v4850,
  v4851,
  v4852,
  v4853,
  v4854,
  v4855,
  v4856,
  v4857,
  v4858,
  v4859,
  v4860,
  v4861,
  v4862,
  v4863,
  v4864,
  v4865,
  v4866,
  v4867,
  v4868,
  v4869,
  v4870,
  v4871,
  v4872,
  v4873,
  v4874,
  v4875,
  v4876,
  v4877,
  v4878,
  v4879,
  v4880,
  v4881,
  v4882,
  v4883,
  v4884,
  v4885,
  v4886,
  v4887,
  v4888,
  v4889,
  v4890,
  v4891,
  v4892,
  v4893,
  v4894,
  v4895,
  v4896,
  v4897,
  v4898,
  v4899,
  v4900,
  v4901,
  v4902,
  v4903,
  v4904,
  v4905,
  v4906,
  v4907,
  v4908,
  v4909,
  v4910,
  v4911,
  v4912,
  v4913,
  v4914,
  v4915,
  v4916,
  v4917,
  v4918,
  v4919,
  v4920,
  v4921,
  v4922,
  v4923,
  v4924,
  v4925,
  v4926,
  v4927,
  v4928,
  v4929,
  v4930,
  v4931,
  v4932,
  v4933,
  v4934,
  v4935,
  v4936,
  v4937,
  v4938,
  v4939,
  v4940,
  v4941,
  v4942,
  v4943,
  v4944,
  v4945,
  v4946,
  v4947,
  v4948,
  v4949,
  v4950,
  v4951,
  v4952,
  v4953,
  v4954,
  v4955,
  v4956,
  v4957,
  v4958,
  v4959,
  v4960,
  v4961,
  v4962,
  v4963,
  v4964,
  v4965,
  v4966,
  v4967,
  v4968,
  v4969,
  v4970,
  v4971,
  v4972,
  v4973,
  v4974,
  v4975,
  v4976,
  v4977,
  v4978,
  v4979,
  v4980,
  v4981,
  v4982,
  v4983,
  v4984,
  v4985,
  v4986,
  v4987,
  v4988,
  v4989,
  v4990,
  v4991,
  v4992,
  v4993,
  v4994,
  v4995,
  v4996,
  v4997,
  v4998,
  v4999,
  v5000,
  v5001,
  v5002,
  v5003,
  v5004,
  v5005,
  v5006,
  v5007,
  v5008,
  v5009,
  v5010,
  v5011,
  v5012,
  v5013,
  v5014,
  v5015,
  v5016,
  v5017,
  v5018,
  v5019,
  v5020,
  v5021,
  v5022,
  v5023,
  v5024,
  v5025,
  v5026,
  v5027,
  v5028,
  v5029,
  v5030,
  v5031,
  v5032,
  v5033,
  v5034,
  v5035,
  v5036,
  v5037,
  v5038,
  v5039,
  v5040,
  v5041,
  v5042,
  v5043,
  v5044,
  v5045,
  v5046,
  v5047,
  v5048,
  v5049,
  v5050,
  v5051,
  v5052,
  v5053,
  v5054,
  v5055,
  v5056,
  v5057,
  v5058,
  v5059,
  v5060,
  v5061,
  v5062,
  v5063,
  v5064,
  v5065,
  v5066,
  v5067,
  v5068,
  v5069,
  v5070,
  v5071,
  v5072,
  v5073,
  v5074,
  v5075,
  v5076,
  v5077,
  v5078,
  v5079,
  v5080,
  v5081,
  v5082,
  v5083,
  v5084,
  v5085,
  v5086,
  v5087,
  v5088,
  v5089,
  v5090,
  v5091,
  v5092,
  v5093,
  v5094,
  v5095,
  v5096,
  v5097,
  v5098,
  v5099,
  v5100,
  v5101,
  v5102,
  v5103,
  v5104,
  v5105,
  v5106,
  v5107,
  v5108,
  v5109,
  v5110,
  v5111,
  v5112,
  v5113,
  v5114,
  v5115,
  v5116,
  v5117,
  v5118,
  v5119,
  v5120,
  v5121,
  v5122,
  v5123,
  v5124,
  v5125,
  v5126,
  v5127,
  v5128,
  v5129,
  v5130,
  v5131,
  v5132,
  v5133,
  v5134,
  v5135,
  v5136,
  v5137,
  v5138,
  v5139,
  v5140,
  v5141,
  v5142,
  v5143,
  v5144,
  v5145,
  v5146,
  v5147,
  v5148,
  v5149,
  v5150,
  v5151,
  v5152,
  v5153,
  v5154,
  v5155,
  v5156,
  v5157,
  v5158,
  v5159,
  v5160,
  v5161,
  v5162,
  v5163,
  v5164,
  v5165,
  v5166,
  v5167,
  v5168,
  v5169,
  v5170,
  v5171,
  v5172,
  v5173,
  v5174,
  v5175,
  v5176,
  v5177,
  v5178,
  v5179,
  v5180,
  v5181,
  v5182,
  v5183,
  v5184,
  v5185,
  v5186,
  v5187,
  v5188,
  v5189,
  v5190,
  v5191,
  v5192,
  v5193,
  v5194,
  v5195,
  v5196,
  v5197,
  v5198,
  v5199,
  v5200,
  v5201,
  v5202,
  v5203,
  v5204,
  v5205,
  v5206,
  v5207,
  v5208,
  v5209,
  v5210,
  v5211,
  v5212,
  v5213,
  v5214,
  v5215,
  v5216,
  v5217,
  v5218,
  v5219,
  v5220,
  v5221,
  v5222,
  v5223,
  v5224,
  v5225,
  v5226,
  v5227,
  v5228,
  v5229,
  v5230,
  v5231,
  v5232,
  v5233,
  v5234,
  v5235,
  v5236,
  v5237,
  v5238,
  v5239,
  v5240,
  v5241,
  v5242,
  v5243,
  v5244,
  v5245,
  v5246,
  v5247,
  v5248,
  v5249,
  v5250,
  v5251,
  v5252,
  v5253,
  v5254,
  v5255,
  v5256,
  v5257,
  v5258,
  v5259,
  v5260,
  v5261,
  v5262,
  v5263,
  v5264,
  v5265,
  v5266,
  v5267,
  v5268,
  v5269,
  v5270,
  v5271,
  v5272,
  v5273,
  v5274,
  v5275,
  v5276,
  v5277,
  v5278,
  v5279,
  v5280,
  v5281,
  v5282,
  v5283,
  v5284,
  v5285,
  v5286,
  v5287,
  v5288,
  v5289,
  v5290,
  v5291,
  v5292,
  v5293,
  v5294,
  v5295,
  v5296,
  v5297,
  v5298,
  v5299,
  v5300,
  v5301,
  v5302,
  v5303,
  v5304,
  v5305,
  v5306,
  v5307,
  v5308,
  v5309,
  v5310,
  v5311,
  v5312,
  v5313,
  v5314,
  v5315,
  v5316,
  v5317,
  v5318,
  v5319,
  v5320,
  v5321,
  v5322,
  v5323,
  v5324,
  v5325,
  v5326,
  v5327,
  v5328,
  v5329,
  v5330,
  v5331,
  v5332,
  v5333,
  v5334,
  v5335,
  v5336,
  v5337,
  v5338,
  v5339,
  v5340,
  v5341,
  v5342,
  v5343,
  v5344,
  v5345,
  v5346,
  v5347,
  v5348,
  v5349,
  v5350,
  v5351,
  v5352,
  v5353,
  v5354,
  v5355,
  v5356,
  v5357,
  v5358,
  v5359,
  v5360,
  v5361,
  v5362,
  v5363,
  v5364,
  v5365,
  v5366,
  v5367,
  v5368,
  v5369,
  v5370,
  v5371,
  v5372,
  v5373;
assign
  v5374 = (v5375 & i22) | (v5285 & ~i22),
  v5375 = (v5376 & i25) | (v5287 & ~i25),
  v5376 = (v5070 & i26) | (v4187 & ~i26),
  v5377 = (v5378 & i21) | (v5283 & ~i21),
  v5378 = (v5379 & i22) | (v5285 & ~i22),
  v5379 = (v5380 & i25) | (v5287 & ~i25),
  v5380 = (v5076 & i26) | (v4195 & ~i26),
  v5381 = (v5382 & i21) | (v5283 & ~i21),
  v5382 = (v5383 & i22) | (v5285 & ~i22),
  v5383 = (v5384 & i25) | (v5287 & ~i25),
  v5384 = (v5082 & i26) | (v4203 & ~i26),
  v5385 = (v5405 & i17) | (v5386 & ~i17),
  v5386 = (v5396 & i19) | (v5387 & ~i19),
  v5387 = (v5392 & i20) | (v5388 & ~i20),
  v5388 = (v5389 & i21) | (v5283 & ~i21),
  v5389 = (v5390 & i22) | (v5285 & ~i22),
  v5390 = (v5391 & i25) | (v5287 & ~i25),
  v5391 = (v5091 & i26) | (v4212 & ~i26),
  v5392 = (v5393 & i21) | (v5283 & ~i21),
  v5393 = (v5394 & i22) | (v5285 & ~i22),
  v5394 = (v5395 & i25) | (v5287 & ~i25),
  v5395 = (v5097 & i26) | (v4221 & ~i26),
  v5396 = (v5401 & i20) | (v5397 & ~i20),
  v5397 = (v5398 & i21) | (v5283 & ~i21),
  v5398 = (v5399 & i22) | (v5285 & ~i22),
  v5399 = (v5400 & i25) | (v5287 & ~i25),
  v5400 = (v5104 & i26) | (v4231 & ~i26),
  v5401 = (v5402 & i21) | (v5283 & ~i21),
  v5402 = (v5403 & i22) | (v5285 & ~i22),
  v5403 = (v5404 & i25) | (v5287 & ~i25),
  v5404 = (v5110 & i26) | (v4239 & ~i26),
  v5405 = (v5415 & i19) | (v5406 & ~i19),
  v5406 = (v5411 & i20) | (v5407 & ~i20),
  v5407 = (v5408 & i21) | (v5283 & ~i21),
  v5408 = (v5409 & i22) | (v5285 & ~i22),
  v5409 = (v5410 & i25) | (v5287 & ~i25),
  v5410 = (v5118 & i26) | (v4249 & ~i26),
  v5411 = (v5412 & i21) | (v5283 & ~i21),
  v5412 = (v5413 & i22) | (v5285 & ~i22),
  v5413 = (v5414 & i25) | (v5287 & ~i25),
  v5414 = (v5124 & i26) | (v4257 & ~i26),
  v5415 = (v5416 & i21) | (v5283 & ~i21),
  v5416 = (v5417 & i22) | (v5285 & ~i22),
  v5417 = (v5418 & i25) | (v5287 & ~i25),
  v5418 = (v5130 & i26) | (v4265 & ~i26),
  v5419 = (v5729 & i11) | (v5420 & ~i11),
  v5420 = (v5421 & i12) | (v4521 & ~i12),
  v5421 = (v4523 & i13) | (v5422 & ~i13),
  v5422 = (v5618 & i14) | (v5423 & ~i14),
  v5423 = (v5521 & i15) | (v5424 & ~i15),
  v5424 = (v5473 & i16) | (v5425 & ~i16),
  v5425 = (v5453 & i17) | (v5426 & ~i17),
  v5426 = (v5440 & i19) | (v5427 & ~i19),
  v5427 = (v5434 & i20) | (v5428 & ~i20),
  v5428 = (v5429 & i21) | (v4932 & ~i21),
  v5429 = (v5430 & i22) | (v4938 & ~i22),
  v5430 = (v4530 & i26) | (v5431 & ~i26),
  v5431 = (v4530 & i27) | (v5432 & ~i27),
  v5432 = (v5433 & i29) | (v4947 & ~i29),
  v5433 = (v4935 & i30) | (v4532 & ~i30),
  v5434 = (v5435 & i21) | (v4932 & ~i21),
  v5435 = (v5436 & i22) | (v4938 & ~i22),
  v5436 = (v4537 & i26) | (v5437 & ~i26),
  v5437 = (v4537 & i27) | (v5438 & ~i27),
  v5438 = (v5439 & i29) | (v4953 & ~i29),
  v5439 = (v4935 & i30) | (v4539 & ~i30),
  v5440 = (v5447 & i20) | (v5441 & ~i20),
  v5441 = (v5442 & i21) | (v4932 & ~i21),
  v5442 = (v5443 & i22) | (v4938 & ~i22),
  v5443 = (v4545 & i26) | (v5444 & ~i26),
  v5444 = (v4545 & i27) | (v5445 & ~i27),
  v5445 = (v5446 & i29) | (v4960 & ~i29),
  v5446 = (v4935 & i30) | (v4547 & ~i30),
  v5447 = (v5448 & i21) | (v4932 & ~i21),
  v5448 = (v5449 & i22) | (v4938 & ~i22),
  v5449 = (v4552 & i26) | (v5450 & ~i26),
  v5450 = (v4552 & i27) | (v5451 & ~i27),
  v5451 = (v5452 & i29) | (v4966 & ~i29),
  v5452 = (v4935 & i30) | (v4554 & ~i30),
  v5453 = (v5467 & i19) | (v5454 & ~i19),
  v5454 = (v5461 & i20) | (v5455 & ~i20),
  v5455 = (v5456 & i21) | (v4932 & ~i21),
  v5456 = (v5457 & i22) | (v4938 & ~i22),
  v5457 = (v4561 & i26) | (v5458 & ~i26),
  v5458 = (v4561 & i27) | (v5459 & ~i27),
  v5459 = (v5460 & i29) | (v4974 & ~i29),
  v5460 = (v4935 & i30) | (v4563 & ~i30),
  v5461 = (v5462 & i21) | (v4932 & ~i21),
  v5462 = (v5463 & i22) | (v4938 & ~i22),
  v5463 = (v4568 & i26) | (v5464 & ~i26),
  v5464 = (v4568 & i27) | (v5465 & ~i27),
  v5465 = (v5466 & i29) | (v4980 & ~i29),
  v5466 = (v4935 & i30) | (v4570 & ~i30),
  v5467 = (v5468 & i21) | (v4932 & ~i21),
  v5468 = (v5469 & i22) | (v4938 & ~i22),
  v5469 = (v4575 & i26) | (v5470 & ~i26),
  v5470 = (v4575 & i27) | (v5471 & ~i27),
  v5471 = (v5472 & i29) | (v4986 & ~i29),
  v5472 = (v4935 & i30) | (v4577 & ~i30),
  v5473 = (v5501 & i17) | (v5474 & ~i17),
  v5474 = (v5488 & i19) | (v5475 & ~i19),
  v5475 = (v5482 & i20) | (v5476 & ~i20),
  v5476 = (v5477 & i21) | (v4932 & ~i21),
  v5477 = (v5478 & i22) | (v4938 & ~i22),
  v5478 = (v4585 & i26) | (v5479 & ~i26),
  v5479 = (v4585 & i27) | (v5480 & ~i27),
  v5480 = (v5481 & i29) | (v4995 & ~i29),
  v5481 = (v4935 & i30) | (v4587 & ~i30),
  v5482 = (v5483 & i21) | (v4932 & ~i21),
  v5483 = (v5484 & i22) | (v4938 & ~i22),
  v5484 = (v4592 & i26) | (v5485 & ~i26),
  v5485 = (v4592 & i27) | (v5486 & ~i27),
  v5486 = (v5487 & i29) | (v5001 & ~i29),
  v5487 = (v4935 & i30) | (v4594 & ~i30),
  v5488 = (v5495 & i20) | (v5489 & ~i20),
  v5489 = (v5490 & i21) | (v4932 & ~i21),
  v5490 = (v5491 & i22) | (v4938 & ~i22),
  v5491 = (v4600 & i26) | (v5492 & ~i26),
  v5492 = (v4600 & i27) | (v5493 & ~i27),
  v5493 = (v5494 & i29) | (v5008 & ~i29),
  v5494 = (v4935 & i30) | (v4602 & ~i30),
  v5495 = (v5496 & i21) | (v4932 & ~i21),
  v5496 = (v5497 & i22) | (v4938 & ~i22),
  v5497 = (v4607 & i26) | (v5498 & ~i26),
  v5498 = (v4607 & i27) | (v5499 & ~i27),
  v5499 = (v5500 & i29) | (v5014 & ~i29),
  v5500 = (v4935 & i30) | (v4609 & ~i30),
  v5501 = (v5515 & i19) | (v5502 & ~i19),
  v5502 = (v5509 & i20) | (v5503 & ~i20),
  v5503 = (v5504 & i21) | (v4932 & ~i21),
  v5504 = (v5505 & i22) | (v4938 & ~i22),
  v5505 = (v4616 & i26) | (v5506 & ~i26),
  v5506 = (v4616 & i27) | (v5507 & ~i27),
  v5507 = (v5508 & i29) | (v5022 & ~i29),
  v5508 = (v4935 & i30) | (v4618 & ~i30),
  v5509 = (v5510 & i21) | (v4932 & ~i21),
  v5510 = (v5511 & i22) | (v4938 & ~i22),
  v5511 = (v4623 & i26) | (v5512 & ~i26),
  v5512 = (v4623 & i27) | (v5513 & ~i27),
  v5513 = (v5514 & i29) | (v5028 & ~i29),
  v5514 = (v4935 & i30) | (v4625 & ~i30),
  v5515 = (v5516 & i21) | (v4932 & ~i21),
  v5516 = (v5517 & i22) | (v4938 & ~i22),
  v5517 = (v4630 & i26) | (v5518 & ~i26),
  v5518 = (v4630 & i27) | (v5519 & ~i27),
  v5519 = (v5520 & i29) | (v5034 & ~i29),
  v5520 = (v4935 & i30) | (v4632 & ~i30),
  v5521 = (v5570 & i16) | (v5522 & ~i16),
  v5522 = (v5550 & i17) | (v5523 & ~i17),
  v5523 = (v5537 & i19) | (v5524 & ~i19),
  v5524 = (v5531 & i20) | (v5525 & ~i20),
  v5525 = (v5526 & i21) | (v4932 & ~i21),
  v5526 = (v5527 & i22) | (v4938 & ~i22),
  v5527 = (v4641 & i26) | (v5528 & ~i26),
  v5528 = (v4641 & i27) | (v5529 & ~i27),
  v5529 = (v5530 & i29) | (v5044 & ~i29),
  v5530 = (v4935 & i30) | (v4643 & ~i30),
  v5531 = (v5532 & i21) | (v4932 & ~i21),
  v5532 = (v5533 & i22) | (v4938 & ~i22),
  v5533 = (v4648 & i26) | (v5534 & ~i26),
  v5534 = (v4648 & i27) | (v5535 & ~i27),
  v5535 = (v5536 & i29) | (v5050 & ~i29),
  v5536 = (v4935 & i30) | (v4650 & ~i30),
  v5537 = (v5544 & i20) | (v5538 & ~i20),
  v5538 = (v5539 & i21) | (v4932 & ~i21),
  v5539 = (v5540 & i22) | (v4938 & ~i22),
  v5540 = (v4656 & i26) | (v5541 & ~i26),
  v5541 = (v4656 & i27) | (v5542 & ~i27),
  v5542 = (v5543 & i29) | (v5057 & ~i29),
  v5543 = (v4935 & i30) | (v4658 & ~i30),
  v5544 = (v5545 & i21) | (v4932 & ~i21),
  v5545 = (v5546 & i22) | (v4938 & ~i22),
  v5546 = (v4663 & i26) | (v5547 & ~i26),
  v5547 = (v4663 & i27) | (v5548 & ~i27),
  v5548 = (v5549 & i29) | (v5063 & ~i29),
  v5549 = (v4935 & i30) | (v4665 & ~i30),
  v5550 = (v5564 & i19) | (v5551 & ~i19),
  v5551 = (v5558 & i20) | (v5552 & ~i20),
  v5552 = (v5553 & i21) | (v4932 & ~i21),
  v5553 = (v5554 & i22) | (v4938 & ~i22),
  v5554 = (v4672 & i26) | (v5555 & ~i26),
  v5555 = (v4672 & i27) | (v5556 & ~i27),
  v5556 = (v5557 & i29) | (v5071 & ~i29),
  v5557 = (v4935 & i30) | (v4674 & ~i30),
  v5558 = (v5559 & i21) | (v4932 & ~i21),
  v5559 = (v5560 & i22) | (v4938 & ~i22),
  v5560 = (v4679 & i26) | (v5561 & ~i26),
  v5561 = (v4679 & i27) | (v5562 & ~i27),
  v5562 = (v5563 & i29) | (v5077 & ~i29),
  v5563 = (v4935 & i30) | (v4681 & ~i30),
  v5564 = (v5565 & i21) | (v4932 & ~i21),
  v5565 = (v5566 & i22) | (v4938 & ~i22),
  v5566 = (v4686 & i26) | (v5567 & ~i26),
  v5567 = (v4686 & i27) | (v5568 & ~i27),
  v5568 = (v5569 & i29) | (v5083 & ~i29),
  v5569 = (v4935 & i30) | (v4688 & ~i30),
  v5570 = (v5598 & i17) | (v5571 & ~i17),
  v5571 = (v5585 & i19) | (v5572 & ~i19),
  v5572 = (v5579 & i20) | (v5573 & ~i20),
  v5573 = (v5574 & i21) | (v4932 & ~i21),
  v5574 = (v5575 & i22) | (v4938 & ~i22),
  v5575 = (v4696 & i26) | (v5576 & ~i26),
  v5576 = (v4696 & i27) | (v5577 & ~i27),
  v5577 = (v5578 & i29) | (v5092 & ~i29),
  v5578 = (v4935 & i30) | (v4698 & ~i30),
  v5579 = (v5580 & i21) | (v4932 & ~i21),
  v5580 = (v5581 & i22) | (v4938 & ~i22),
  v5581 = (v4703 & i26) | (v5582 & ~i26),
  v5582 = (v4703 & i27) | (v5583 & ~i27),
  v5583 = (v5584 & i29) | (v5098 & ~i29),
  v5584 = (v4935 & i30) | (v4705 & ~i30),
  v5585 = (v5592 & i20) | (v5586 & ~i20),
  v5586 = (v5587 & i21) | (v4932 & ~i21),
  v5587 = (v5588 & i22) | (v4938 & ~i22),
  v5588 = (v4711 & i26) | (v5589 & ~i26),
  v5589 = (v4711 & i27) | (v5590 & ~i27),
  v5590 = (v5591 & i29) | (v5105 & ~i29),
  v5591 = (v4935 & i30) | (v4713 & ~i30),
  v5592 = (v5593 & i21) | (v4932 & ~i21),
  v5593 = (v5594 & i22) | (v4938 & ~i22),
  v5594 = (v4718 & i26) | (v5595 & ~i26),
  v5595 = (v4718 & i27) | (v5596 & ~i27),
  v5596 = (v5597 & i29) | (v5111 & ~i29),
  v5597 = (v4935 & i30) | (v4720 & ~i30),
  v5598 = (v5612 & i19) | (v5599 & ~i19),
  v5599 = (v5606 & i20) | (v5600 & ~i20),
  v5600 = (v5601 & i21) | (v4932 & ~i21),
  v5601 = (v5602 & i22) | (v4938 & ~i22),
  v5602 = (v4727 & i26) | (v5603 & ~i26),
  v5603 = (v4727 & i27) | (v5604 & ~i27),
  v5604 = (v5605 & i29) | (v5119 & ~i29),
  v5605 = (v4935 & i30) | (v4729 & ~i30),
  v5606 = (v5607 & i21) | (v4932 & ~i21),
  v5607 = (v5608 & i22) | (v4938 & ~i22),
  v5608 = (v4734 & i26) | (v5609 & ~i26),
  v5609 = (v4734 & i27) | (v5610 & ~i27),
  v5610 = (v5611 & i29) | (v5125 & ~i29),
  v5611 = (v4935 & i30) | (v4736 & ~i30),
  v5612 = (v5613 & i21) | (v4932 & ~i21),
  v5613 = (v5614 & i22) | (v4938 & ~i22),
  v5614 = (v4741 & i26) | (v5615 & ~i26),
  v5615 = (v4741 & i27) | (v5616 & ~i27),
  v5616 = (v5617 & i29) | (v5131 & ~i29),
  v5617 = (v4935 & i30) | (v4743 & ~i30),
  v5618 = (v5674 & i15) | (v5619 & ~i15),
  v5619 = (v5647 & i16) | (v5620 & ~i16),
  v5620 = (v5636 & i17) | (v5621 & ~i17),
  v5621 = (v5629 & i19) | (v5622 & ~i19),
  v5622 = (v5626 & i20) | (v5623 & ~i20),
  v5623 = (v5624 & i21) | (v5138 & ~i21),
  v5624 = (v5625 & i22) | (v5140 & ~i22),
  v5625 = (v5432 & i27) | (v4530 & ~i27),
  v5626 = (v5627 & i21) | (v5138 & ~i21),
  v5627 = (v5628 & i22) | (v5140 & ~i22),
  v5628 = (v5438 & i27) | (v4537 & ~i27),
  v5629 = (v5633 & i20) | (v5630 & ~i20),
  v5630 = (v5631 & i21) | (v5138 & ~i21),
  v5631 = (v5632 & i22) | (v5140 & ~i22),
  v5632 = (v5445 & i27) | (v4545 & ~i27),
  v5633 = (v5634 & i21) | (v5138 & ~i21),
  v5634 = (v5635 & i22) | (v5140 & ~i22),
  v5635 = (v5451 & i27) | (v4552 & ~i27),
  v5636 = (v5644 & i19) | (v5637 & ~i19),
  v5637 = (v5641 & i20) | (v5638 & ~i20),
  v5638 = (v5639 & i21) | (v5138 & ~i21),
  v5639 = (v5640 & i22) | (v5140 & ~i22),
  v5640 = (v5459 & i27) | (v4561 & ~i27),
  v5641 = (v5642 & i21) | (v5138 & ~i21),
  v5642 = (v5643 & i22) | (v5140 & ~i22),
  v5643 = (v5465 & i27) | (v4568 & ~i27),
  v5644 = (v5645 & i21) | (v5138 & ~i21),
  v5645 = (v5646 & i22) | (v5140 & ~i22),
  v5646 = (v5471 & i27) | (v4575 & ~i27),
  v5647 = (v5663 & i17) | (v5648 & ~i17),
  v5648 = (v5656 & i19) | (v5649 & ~i19),
  v5649 = (v5653 & i20) | (v5650 & ~i20),
  v5650 = (v5651 & i21) | (v5138 & ~i21),
  v5651 = (v5652 & i22) | (v5140 & ~i22),
  v5652 = (v5480 & i27) | (v4585 & ~i27),
  v5653 = (v5654 & i21) | (v5138 & ~i21),
  v5654 = (v5655 & i22) | (v5140 & ~i22),
  v5655 = (v5486 & i27) | (v4592 & ~i27),
  v5656 = (v5660 & i20) | (v5657 & ~i20),
  v5657 = (v5658 & i21) | (v5138 & ~i21),
  v5658 = (v5659 & i22) | (v5140 & ~i22),
  v5659 = (v5493 & i27) | (v4600 & ~i27),
  v5660 = (v5661 & i21) | (v5138 & ~i21),
  v5661 = (v5662 & i22) | (v5140 & ~i22),
  v5662 = (v5499 & i27) | (v4607 & ~i27),
  v5663 = (v5671 & i19) | (v5664 & ~i19),
  v5664 = (v5668 & i20) | (v5665 & ~i20),
  v5665 = (v5666 & i21) | (v5138 & ~i21),
  v5666 = (v5667 & i22) | (v5140 & ~i22),
  v5667 = (v5507 & i27) | (v4616 & ~i27),
  v5668 = (v5669 & i21) | (v5138 & ~i21),
  v5669 = (v5670 & i22) | (v5140 & ~i22),
  v5670 = (v5513 & i27) | (v4623 & ~i27),
  v5671 = (v5672 & i21) | (v5138 & ~i21),
  v5672 = (v5673 & i22) | (v5140 & ~i22),
  v5673 = (v5519 & i27) | (v4630 & ~i27),
  v5674 = (v5702 & i16) | (v5675 & ~i16),
  v5675 = (v5691 & i17) | (v5676 & ~i17),
  v5676 = (v5684 & i19) | (v5677 & ~i19),
  v5677 = (v5681 & i20) | (v5678 & ~i20),
  v5678 = (v5679 & i21) | (v5138 & ~i21),
  v5679 = (v5680 & i22) | (v5140 & ~i22),
  v5680 = (v5529 & i27) | (v4641 & ~i27),
  v5681 = (v5682 & i21) | (v5138 & ~i21),
  v5682 = (v5683 & i22) | (v5140 & ~i22),
  v5683 = (v5535 & i27) | (v4648 & ~i27),
  v5684 = (v5688 & i20) | (v5685 & ~i20),
  v5685 = (v5686 & i21) | (v5138 & ~i21),
  v5686 = (v5687 & i22) | (v5140 & ~i22),
  v5687 = (v5542 & i27) | (v4656 & ~i27),
  v5688 = (v5689 & i21) | (v5138 & ~i21),
  v5689 = (v5690 & i22) | (v5140 & ~i22),
  v5690 = (v5548 & i27) | (v4663 & ~i27),
  v5691 = (v5699 & i19) | (v5692 & ~i19),
  v5692 = (v5696 & i20) | (v5693 & ~i20),
  v5693 = (v5694 & i21) | (v5138 & ~i21),
  v5694 = (v5695 & i22) | (v5140 & ~i22),
  v5695 = (v5556 & i27) | (v4672 & ~i27),
  v5696 = (v5697 & i21) | (v5138 & ~i21),
  v5697 = (v5698 & i22) | (v5140 & ~i22),
  v5698 = (v5562 & i27) | (v4679 & ~i27),
  v5699 = (v5700 & i21) | (v5138 & ~i21),
  v5700 = (v5701 & i22) | (v5140 & ~i22),
  v5701 = (v5568 & i27) | (v4686 & ~i27),
  v5702 = (v5718 & i17) | (v5703 & ~i17),
  v5703 = (v5711 & i19) | (v5704 & ~i19),
  v5704 = (v5708 & i20) | (v5705 & ~i20),
  v5705 = (v5706 & i21) | (v5138 & ~i21),
  v5706 = (v5707 & i22) | (v5140 & ~i22),
  v5707 = (v5577 & i27) | (v4696 & ~i27),
  v5708 = (v5709 & i21) | (v5138 & ~i21),
  v5709 = (v5710 & i22) | (v5140 & ~i22),
  v5710 = (v5583 & i27) | (v4703 & ~i27),
  v5711 = (v5715 & i20) | (v5712 & ~i20),
  v5712 = (v5713 & i21) | (v5138 & ~i21),
  v5713 = (v5714 & i22) | (v5140 & ~i22),
  v5714 = (v5590 & i27) | (v4711 & ~i27),
  v5715 = (v5716 & i21) | (v5138 & ~i21),
  v5716 = (v5717 & i22) | (v5140 & ~i22),
  v5717 = (v5596 & i27) | (v4718 & ~i27),
  v5718 = (v5726 & i19) | (v5719 & ~i19),
  v5719 = (v5723 & i20) | (v5720 & ~i20),
  v5720 = (v5721 & i21) | (v5138 & ~i21),
  v5721 = (v5722 & i22) | (v5140 & ~i22),
  v5722 = (v5604 & i27) | (v4727 & ~i27),
  v5723 = (v5724 & i21) | (v5138 & ~i21),
  v5724 = (v5725 & i22) | (v5140 & ~i22),
  v5725 = (v5610 & i27) | (v4734 & ~i27),
  v5726 = (v5727 & i21) | (v5138 & ~i21),
  v5727 = (v5728 & i22) | (v5140 & ~i22),
  v5728 = (v5616 & i27) | (v4741 & ~i27),
  v5729 = (v4523 & i12) | (v5730 & ~i12),
  v5730 = (v4523 & i13) | (v5731 & ~i13),
  v5731 = (v5732 & i14) | (v4523 & ~i14),
  v5732 = (v5788 & i15) | (v5733 & ~i15),
  v5733 = (v5761 & i16) | (v5734 & ~i16),
  v5734 = (v5750 & i17) | (v5735 & ~i17),
  v5735 = (v5743 & i19) | (v5736 & ~i19),
  v5736 = (v5740 & i20) | (v5737 & ~i20),
  v5737 = (v5738 & i21) | (v5283 & ~i21),
  v5738 = (v5739 & i22) | (v5285 & ~i22),
  v5739 = (v5431 & i26) | (v4530 & ~i26),
  v5740 = (v5741 & i21) | (v5283 & ~i21),
  v5741 = (v5742 & i22) | (v5285 & ~i22),
  v5742 = (v5437 & i26) | (v4537 & ~i26),
  v5743 = (v5747 & i20) | (v5744 & ~i20),
  v5744 = (v5745 & i21) | (v5283 & ~i21),
  v5745 = (v5746 & i22) | (v5285 & ~i22),
  v5746 = (v5444 & i26) | (v4545 & ~i26),
  v5747 = (v5748 & i21) | (v5283 & ~i21),
  v5748 = (v5749 & i22) | (v5285 & ~i22),
  v5749 = (v5450 & i26) | (v4552 & ~i26),
  v5750 = (v5758 & i19) | (v5751 & ~i19),
  v5751 = (v5755 & i20) | (v5752 & ~i20),
  v5752 = (v5753 & i21) | (v5283 & ~i21),
  v5753 = (v5754 & i22) | (v5285 & ~i22),
  v5754 = (v5458 & i26) | (v4561 & ~i26),
  v5755 = (v5756 & i21) | (v5283 & ~i21),
  v5756 = (v5757 & i22) | (v5285 & ~i22),
  v5757 = (v5464 & i26) | (v4568 & ~i26),
  v5758 = (v5759 & i21) | (v5283 & ~i21),
  v5759 = (v5760 & i22) | (v5285 & ~i22),
  v5760 = (v5470 & i26) | (v4575 & ~i26),
  v5761 = (v5777 & i17) | (v5762 & ~i17),
  v5762 = (v5770 & i19) | (v5763 & ~i19),
  v5763 = (v5767 & i20) | (v5764 & ~i20),
  v5764 = (v5765 & i21) | (v5283 & ~i21),
  v5765 = (v5766 & i22) | (v5285 & ~i22),
  v5766 = (v5479 & i26) | (v4585 & ~i26),
  v5767 = (v5768 & i21) | (v5283 & ~i21),
  v5768 = (v5769 & i22) | (v5285 & ~i22),
  v5769 = (v5485 & i26) | (v4592 & ~i26),
  v5770 = (v5774 & i20) | (v5771 & ~i20),
  v5771 = (v5772 & i21) | (v5283 & ~i21),
  v5772 = (v5773 & i22) | (v5285 & ~i22),
  v5773 = (v5492 & i26) | (v4600 & ~i26),
  v5774 = (v5775 & i21) | (v5283 & ~i21),
  v5775 = (v5776 & i22) | (v5285 & ~i22),
  v5776 = (v5498 & i26) | (v4607 & ~i26),
  v5777 = (v5785 & i19) | (v5778 & ~i19),
  v5778 = (v5782 & i20) | (v5779 & ~i20),
  v5779 = (v5780 & i21) | (v5283 & ~i21),
  v5780 = (v5781 & i22) | (v5285 & ~i22),
  v5781 = (v5506 & i26) | (v4616 & ~i26),
  v5782 = (v5783 & i21) | (v5283 & ~i21),
  v5783 = (v5784 & i22) | (v5285 & ~i22),
  v5784 = (v5512 & i26) | (v4623 & ~i26),
  v5785 = (v5786 & i21) | (v5283 & ~i21),
  v5786 = (v5787 & i22) | (v5285 & ~i22),
  v5787 = (v5518 & i26) | (v4630 & ~i26),
  v5788 = (v5816 & i16) | (v5789 & ~i16),
  v5789 = (v5805 & i17) | (v5790 & ~i17),
  v5790 = (v5798 & i19) | (v5791 & ~i19),
  v5791 = (v5795 & i20) | (v5792 & ~i20),
  v5792 = (v5793 & i21) | (v5283 & ~i21),
  v5793 = (v5794 & i22) | (v5285 & ~i22),
  v5794 = (v5528 & i26) | (v4641 & ~i26),
  v5795 = (v5796 & i21) | (v5283 & ~i21),
  v5796 = (v5797 & i22) | (v5285 & ~i22),
  v5797 = (v5534 & i26) | (v4648 & ~i26),
  v5798 = (v5802 & i20) | (v5799 & ~i20),
  v5799 = (v5800 & i21) | (v5283 & ~i21),
  v5800 = (v5801 & i22) | (v5285 & ~i22),
  v5801 = (v5541 & i26) | (v4656 & ~i26),
  v5802 = (v5803 & i21) | (v5283 & ~i21),
  v5803 = (v5804 & i22) | (v5285 & ~i22),
  v5804 = (v5547 & i26) | (v4663 & ~i26),
  v5805 = (v5813 & i19) | (v5806 & ~i19),
  v5806 = (v5810 & i20) | (v5807 & ~i20),
  v5807 = (v5808 & i21) | (v5283 & ~i21),
  v5808 = (v5809 & i22) | (v5285 & ~i22),
  v5809 = (v5555 & i26) | (v4672 & ~i26),
  v5810 = (v5811 & i21) | (v5283 & ~i21),
  v5811 = (v5812 & i22) | (v5285 & ~i22),
  v5812 = (v5561 & i26) | (v4679 & ~i26),
  v5813 = (v5814 & i21) | (v5283 & ~i21),
  v5814 = (v5815 & i22) | (v5285 & ~i22),
  v5815 = (v5567 & i26) | (v4686 & ~i26),
  v5816 = (v5832 & i17) | (v5817 & ~i17),
  v5817 = (v5825 & i19) | (v5818 & ~i19),
  v5818 = (v5822 & i20) | (v5819 & ~i20),
  v5819 = (v5820 & i21) | (v5283 & ~i21),
  v5820 = (v5821 & i22) | (v5285 & ~i22),
  v5821 = (v5576 & i26) | (v4696 & ~i26),
  v5822 = (v5823 & i21) | (v5283 & ~i21),
  v5823 = (v5824 & i22) | (v5285 & ~i22),
  v5824 = (v5582 & i26) | (v4703 & ~i26),
  v5825 = (v5829 & i20) | (v5826 & ~i20),
  v5826 = (v5827 & i21) | (v5283 & ~i21),
  v5827 = (v5828 & i22) | (v5285 & ~i22),
  v5828 = (v5589 & i26) | (v4711 & ~i26),
  v5829 = (v5830 & i21) | (v5283 & ~i21),
  v5830 = (v5831 & i22) | (v5285 & ~i22),
  v5831 = (v5595 & i26) | (v4718 & ~i26),
  v5832 = (v5840 & i19) | (v5833 & ~i19),
  v5833 = (v5837 & i20) | (v5834 & ~i20),
  v5834 = (v5835 & i21) | (v5283 & ~i21),
  v5835 = (v5836 & i22) | (v5285 & ~i22),
  v5836 = (v5603 & i26) | (v4727 & ~i26),
  v5837 = (v5838 & i21) | (v5283 & ~i21),
  v5838 = (v5839 & i22) | (v5285 & ~i22),
  v5839 = (v5609 & i26) | (v4734 & ~i26),
  v5840 = (v5841 & i21) | (v5283 & ~i21),
  v5841 = (v5842 & i22) | (v5285 & ~i22),
  v5842 = (v5615 & i26) | (v4741 & ~i26),
  v5843 = (v5851 & i11) | (v5844 & ~i11),
  v5844 = (v5845 & i12) | (v4831 & ~i12),
  v5845 = (v4833 & i13) | (v5846 & ~i13),
  v5846 = (v5849 & i14) | (v5847 & ~i14),
  v5847 = (v5848 & i21) | (v4932 & ~i21),
  v5848 = (v4942 & i22) | (v4938 & ~i22),
  v5849 = (v5850 & i21) | (v5138 & ~i21),
  v5850 = (v5142 & i22) | (v5140 & ~i22),
  v5851 = (v4833 & i12) | (v5852 & ~i12),
  v5852 = (v4833 & i13) | (v5853 & ~i13),
  v5853 = (v5854 & i14) | (v4833 & ~i14),
  v5854 = (v5855 & i21) | (v5283 & ~i21),
  v5855 = (v5287 & i22) | (v5285 & ~i22),
  v5856 = (v5843 & i9) | (v5857 & ~i9),
  v5857 = (v6142 & i10) | (v5858 & ~i10),
  v5858 = (v6128 & i11) | (v5859 & ~i11),
  v5859 = (v6098 & i12) | (v5860 & ~i12),
  v5860 = (v5862 & i13) | (v5861 & ~i13),
  v5861 = (v5875 & i14) | (v5862 & ~i14),
  v5862 = (v5868 & i21) | (v5863 & ~i21),
  v5863 = (v27 & i23) | (v5864 & ~i23),
  v5864 = (v27 & i24) | (v5865 & ~i24),
  v5865 = (v5866 & i30) | (v27 & ~i30),
  v5866 = (v27 & i31) | (v5867 & ~i31),
  v5867 = v63 & i32,
  v5868 = (v5872 & i22) | (v5869 & ~i22),
  v5869 = (v3908 & i23) | (v5870 & ~i23),
  v5870 = (v3908 & i24) | (v5871 & ~i24),
  v5871 = (v5866 & i30) | (v3909 & ~i30),
  v5872 = (v3912 & i23) | (v5873 & ~i23),
  v5873 = (v3912 & i24) | (v5874 & ~i24),
  v5874 = (v5866 & i30) | (v3913 & ~i30),
  v5875 = (v5987 & i15) | (v5876 & ~i15),
  v5876 = (v5932 & i16) | (v5877 & ~i16),
  v5877 = (v5909 & i17) | (v5878 & ~i17),
  v5878 = (v5894 & i19) | (v5879 & ~i19),
  v5879 = (v5887 & i20) | (v5880 & ~i20),
  v5880 = (v5881 & i21) | (v5863 & ~i21),
  v5881 = (v5882 & i22) | (v5869 & ~i22),
  v5882 = (v4276 & i23) | (v5883 & ~i23),
  v5883 = (v4276 & i24) | (v5884 & ~i24),
  v5884 = (v5886 & i29) | (v5885 & ~i29),
  v5885 = (v5866 & i30) | (v3921 & ~i30),
  v5886 = (v5866 & i30) | (v4278 & ~i30),
  v5887 = (v5888 & i21) | (v5863 & ~i21),
  v5888 = (v5889 & i22) | (v5869 & ~i22),
  v5889 = (v4284 & i23) | (v5890 & ~i23),
  v5890 = (v4284 & i24) | (v5891 & ~i24),
  v5891 = (v5893 & i29) | (v5892 & ~i29),
  v5892 = (v5866 & i30) | (v3937 & ~i30),
  v5893 = (v5866 & i30) | (v4286 & ~i30),
  v5894 = (v5902 & i20) | (v5895 & ~i20),
  v5895 = (v5896 & i21) | (v5863 & ~i21),
  v5896 = (v5897 & i22) | (v5869 & ~i22),
  v5897 = (v4293 & i23) | (v5898 & ~i23),
  v5898 = (v4293 & i24) | (v5899 & ~i24),
  v5899 = (v5901 & i29) | (v5900 & ~i29),
  v5900 = (v5866 & i30) | (v3954 & ~i30),
  v5901 = (v5866 & i30) | (v4295 & ~i30),
  v5902 = (v5903 & i21) | (v5863 & ~i21),
  v5903 = (v5904 & i22) | (v5869 & ~i22),
  v5904 = (v4301 & i23) | (v5905 & ~i23),
  v5905 = (v4301 & i24) | (v5906 & ~i24),
  v5906 = (v5908 & i29) | (v5907 & ~i29),
  v5907 = (v5866 & i30) | (v3972 & ~i30),
  v5908 = (v5866 & i30) | (v4303 & ~i30),
  v5909 = (v5925 & i19) | (v5910 & ~i19),
  v5910 = (v5918 & i20) | (v5911 & ~i20),
  v5911 = (v5912 & i21) | (v5863 & ~i21),
  v5912 = (v5913 & i22) | (v5869 & ~i22),
  v5913 = (v4311 & i23) | (v5914 & ~i23),
  v5914 = (v4311 & i24) | (v5915 & ~i24),
  v5915 = (v5917 & i29) | (v5916 & ~i29),
  v5916 = (v5866 & i30) | (v3991 & ~i30),
  v5917 = (v5866 & i30) | (v4313 & ~i30),
  v5918 = (v5919 & i21) | (v5863 & ~i21),
  v5919 = (v5920 & i22) | (v5869 & ~i22),
  v5920 = (v4319 & i23) | (v5921 & ~i23),
  v5921 = (v4319 & i24) | (v5922 & ~i24),
  \[402]  = v2,
  v5922 = (v5924 & i29) | (v5923 & ~i29),
  v5923 = (v5866 & i30) | (v4008 & ~i30),
  v5924 = (v5866 & i30) | (v4321 & ~i30),
  v5925 = (v5926 & i21) | (v5863 & ~i21),
  v5926 = (v5927 & i22) | (v5869 & ~i22),
  v5927 = (v4327 & i23) | (v5928 & ~i23),
  v5928 = (v4327 & i24) | (v5929 & ~i24),
  v5929 = (v5931 & i29) | (v5930 & ~i29),
  v5930 = (v5866 & i30) | (v4025 & ~i30),
  v5931 = (v5866 & i30) | (v4329 & ~i30),
  \[403]  = v14,
  v5932 = (v5964 & i17) | (v5933 & ~i17),
  v5933 = (v5949 & i19) | (v5934 & ~i19),
  v5934 = (v5942 & i20) | (v5935 & ~i20),
  v5935 = (v5936 & i21) | (v5863 & ~i21),
  v5936 = (v5937 & i22) | (v5869 & ~i22),
  v5937 = (v4338 & i23) | (v5938 & ~i23),
  v5938 = (v4338 & i24) | (v5939 & ~i24),
  v5939 = (v5941 & i29) | (v5940 & ~i29),
  v5940 = (v5866 & i30) | (v4039 & ~i30),
  v5941 = (v5866 & i30) | (v4340 & ~i30),
  \[404]  = v31,
  v5942 = (v5943 & i21) | (v5863 & ~i21),
  v5943 = (v5944 & i22) | (v5869 & ~i22),
  v5944 = (v4346 & i23) | (v5945 & ~i23),
  v5945 = (v4346 & i24) | (v5946 & ~i24),
  v5946 = (v5948 & i29) | (v5947 & ~i29),
  v5947 = (v5866 & i30) | (v4052 & ~i30),
  v5948 = (v5866 & i30) | (v4348 & ~i30),
  v5949 = (v5957 & i20) | (v5950 & ~i20),
  v5950 = (v5951 & i21) | (v5863 & ~i21),
  v5951 = (v5952 & i22) | (v5869 & ~i22),
  \[405]  = v43,
  v5952 = (v4355 & i23) | (v5953 & ~i23),
  v5953 = (v4355 & i24) | (v5954 & ~i24),
  v5954 = (v5956 & i29) | (v5955 & ~i29),
  v5955 = (v5866 & i30) | (v4066 & ~i30),
  v5956 = (v5866 & i30) | (v4357 & ~i30),
  v5957 = (v5958 & i21) | (v5863 & ~i21),
  v5958 = (v5959 & i22) | (v5869 & ~i22),
  v5959 = (v4363 & i23) | (v5960 & ~i23),
  v5960 = (v4363 & i24) | (v5961 & ~i24),
  v5961 = (v5963 & i29) | (v5962 & ~i29),
  \[406]  = v59,
  v5962 = (v5866 & i30) | (v4083 & ~i30),
  v5963 = (v5866 & i30) | (v4365 & ~i30),
  v5964 = (v5980 & i19) | (v5965 & ~i19),
  v5965 = (v5973 & i20) | (v5966 & ~i20),
  v5966 = (v5967 & i21) | (v5863 & ~i21),
  v5967 = (v5968 & i22) | (v5869 & ~i22),
  v5968 = (v4373 & i23) | (v5969 & ~i23),
  v5969 = (v4373 & i24) | (v5970 & ~i24),
  v5970 = (v5972 & i29) | (v5971 & ~i29),
  v5971 = (v5866 & i30) | (v4102 & ~i30),
  \[407]  = \*clm_file_1_istate1 ,
  v5972 = (v5866 & i30) | (v4375 & ~i30),
  v5973 = (v5974 & i21) | (v5863 & ~i21),
  v5974 = (v5975 & i22) | (v5869 & ~i22),
  v5975 = (v4381 & i23) | (v5976 & ~i23),
  v5976 = (v4381 & i24) | (v5977 & ~i24),
  v5977 = (v5979 & i29) | (v5978 & ~i29),
  v5978 = (v5866 & i30) | (v4119 & ~i30),
  v5979 = (v5866 & i30) | (v4383 & ~i30),
  v5980 = (v5981 & i21) | (v5863 & ~i21),
  v5981 = (v5982 & i22) | (v5869 & ~i22),
  \[408]  = \*clm_file_1_istate0 ,
  v5982 = (v4389 & i23) | (v5983 & ~i23),
  v5983 = (v4389 & i24) | (v5984 & ~i24),
  v5984 = (v5986 & i29) | (v5985 & ~i29),
  v5985 = (v5866 & i30) | (v4136 & ~i30),
  v5986 = (v5866 & i30) | (v4391 & ~i30),
  v5987 = (v6043 & i16) | (v5988 & ~i16),
  v5988 = (v6020 & i17) | (v5989 & ~i17),
  v5989 = (v6005 & i19) | (v5990 & ~i19),
  v5990 = (v5998 & i20) | (v5991 & ~i20),
  v5991 = (v5992 & i21) | (v5863 & ~i21),
  \[409]  = v243,
  v5992 = (v5993 & i22) | (v5869 & ~i22),
  v5993 = (v4401 & i23) | (v5994 & ~i23),
  v5994 = (v4401 & i24) | (v5995 & ~i24),
  v5995 = (v5997 & i29) | (v5996 & ~i29),
  v5996 = (v5866 & i30) | (v4151 & ~i30),
  v5997 = (v5866 & i30) | (v4403 & ~i30),
  v5998 = (v5999 & i21) | (v5863 & ~i21),
  v5999 = (v6000 & i22) | (v5869 & ~i22),
  \[410]  = v294,
  \[411]  = v345,
  \[412]  = v349,
  \[413]  = v437,
  \[414]  = v499,
  \[415]  = v550,
  \[416]  = v601,
  \[417]  = v2153,
  \[418]  = v3888,
  \[419]  = v6425,
  \[420]  = v6437,
  v2 = (v9 & i20) | (v3 & ~i20),
  v3 = (v7 & i22) | (v4 & ~i22),
  v4 = (v6 & i30) | (v5 & ~i30),
  v5 = (v8 & i31) | (v6 & ~i31),
  v6 = v7 & i47,
  v7 = i48,
  v8 = (v7 & i32) | (v6 & ~i32),
  v9 = (v7 & i22) | (v10 & ~i22),
  \[421]  = v8909,
  \[422]  = v10056,
  \[423]  = v10068,
  \[424]  = v10082,
  \[425]  = v10091,
  \[426]  = v10099,
  \[427]  = v10112,
  \[428]  = v10126,
  \[429]  = v10135,
  \[430]  = v10143,
  \[431]  = v10247,
  \[432]  = v10316,
  \[433]  = \*clm_clk_ctl_time1 ,
  \[434]  = \*clm_clk_ctl_time0 ,
  v6000 = (v4409 & i23) | (v6001 & ~i23),
  v6001 = (v4409 & i24) | (v6002 & ~i24),
  v6002 = (v6004 & i29) | (v6003 & ~i29),
  v6003 = (v5866 & i30) | (v4160 & ~i30),
  v6004 = (v5866 & i30) | (v4411 & ~i30),
  v6005 = (v6013 & i20) | (v6006 & ~i20),
  v6006 = (v6007 & i21) | (v5863 & ~i21),
  v6007 = (v6008 & i22) | (v5869 & ~i22),
  v6008 = (v4418 & i23) | (v6009 & ~i23),
  v6009 = (v4418 & i24) | (v6010 & ~i24),
  v6010 = (v6012 & i29) | (v6011 & ~i29),
  v6011 = (v5866 & i30) | (v4170 & ~i30),
  v6012 = (v5866 & i30) | (v4420 & ~i30),
  v6013 = (v6014 & i21) | (v5863 & ~i21),
  v6014 = (v6015 & i22) | (v5869 & ~i22),
  v6015 = (v4426 & i23) | (v6016 & ~i23),
  v6016 = (v4426 & i24) | (v6017 & ~i24),
  v6017 = (v6019 & i29) | (v6018 & ~i29),
  v6018 = (v5866 & i30) | (v4178 & ~i30),
  v6019 = (v5866 & i30) | (v4428 & ~i30),
  v6020 = (v6036 & i19) | (v6021 & ~i19),
  v6021 = (v6029 & i20) | (v6022 & ~i20),
  v6022 = (v6023 & i21) | (v5863 & ~i21),
  v6023 = (v6024 & i22) | (v5869 & ~i22),
  v6024 = (v4436 & i23) | (v6025 & ~i23),
  v6025 = (v4436 & i24) | (v6026 & ~i24),
  v6026 = (v6028 & i29) | (v6027 & ~i29),
  v6027 = (v5866 & i30) | (v4188 & ~i30),
  v6028 = (v5866 & i30) | (v4438 & ~i30),
  v6029 = (v6030 & i21) | (v5863 & ~i21),
  v6030 = (v6031 & i22) | (v5869 & ~i22),
  v6031 = (v4444 & i23) | (v6032 & ~i23),
  v6032 = (v4444 & i24) | (v6033 & ~i24),
  v6033 = (v6035 & i29) | (v6034 & ~i29),
  v6034 = (v5866 & i30) | (v4196 & ~i30),
  v6035 = (v5866 & i30) | (v4446 & ~i30),
  v6036 = (v6037 & i21) | (v5863 & ~i21),
  v6037 = (v6038 & i22) | (v5869 & ~i22),
  v6038 = (v4452 & i23) | (v6039 & ~i23),
  v6039 = (v4452 & i24) | (v6040 & ~i24),
  v6040 = (v6042 & i29) | (v6041 & ~i29),
  v6041 = (v5866 & i30) | (v4204 & ~i30),
  v6042 = (v5866 & i30) | (v4454 & ~i30),
  v6043 = (v6075 & i17) | (v6044 & ~i17),
  v6044 = (v6060 & i19) | (v6045 & ~i19),
  v6045 = (v6053 & i20) | (v6046 & ~i20),
  v6046 = (v6047 & i21) | (v5863 & ~i21),
  v6047 = (v6048 & i22) | (v5869 & ~i22),
  v6048 = (v4463 & i23) | (v6049 & ~i23),
  v6049 = (v4463 & i24) | (v6050 & ~i24),
  v6050 = (v6052 & i29) | (v6051 & ~i29),
  v6051 = (v5866 & i30) | (v4213 & ~i30),
  v6052 = (v5866 & i30) | (v4465 & ~i30),
  v6053 = (v6054 & i21) | (v5863 & ~i21),
  v6054 = (v6055 & i22) | (v5869 & ~i22),
  v6055 = (v4471 & i23) | (v6056 & ~i23),
  v6056 = (v4471 & i24) | (v6057 & ~i24),
  v6057 = (v6059 & i29) | (v6058 & ~i29),
  v6058 = (v5866 & i30) | (v4222 & ~i30),
  v6059 = (v5866 & i30) | (v4473 & ~i30),
  v6060 = (v6068 & i20) | (v6061 & ~i20),
  v6061 = (v6062 & i21) | (v5863 & ~i21),
  v6062 = (v6063 & i22) | (v5869 & ~i22),
  v6063 = (v4480 & i23) | (v6064 & ~i23),
  v6064 = (v4480 & i24) | (v6065 & ~i24),
  v6065 = (v6067 & i29) | (v6066 & ~i29),
  v6066 = (v5866 & i30) | (v4232 & ~i30),
  v6067 = (v5866 & i30) | (v4482 & ~i30),
  v6068 = (v6069 & i21) | (v5863 & ~i21),
  v6069 = (v6070 & i22) | (v5869 & ~i22),
  v6070 = (v4488 & i23) | (v6071 & ~i23),
  v6071 = (v4488 & i24) | (v6072 & ~i24),
  v6072 = (v6074 & i29) | (v6073 & ~i29),
  v6073 = (v5866 & i30) | (v4240 & ~i30),
  v6074 = (v5866 & i30) | (v4490 & ~i30),
  v6075 = (v6091 & i19) | (v6076 & ~i19),
  v6076 = (v6084 & i20) | (v6077 & ~i20),
  v6077 = (v6078 & i21) | (v5863 & ~i21),
  v6078 = (v6079 & i22) | (v5869 & ~i22),
  v6079 = (v4498 & i23) | (v6080 & ~i23),
  v6080 = (v4498 & i24) | (v6081 & ~i24),
  v6081 = (v6083 & i29) | (v6082 & ~i29),
  v6082 = (v5866 & i30) | (v4250 & ~i30),
  v6083 = (v5866 & i30) | (v4500 & ~i30),
  v6084 = (v6085 & i21) | (v5863 & ~i21),
  v6085 = (v6086 & i22) | (v5869 & ~i22),
  v6086 = (v4506 & i23) | (v6087 & ~i23),
  v6087 = (v4506 & i24) | (v6088 & ~i24),
  v6088 = (v6090 & i29) | (v6089 & ~i29),
  v6089 = (v5866 & i30) | (v4258 & ~i30),
  v6090 = (v5866 & i30) | (v4508 & ~i30),
  v6091 = (v6092 & i21) | (v5863 & ~i21),
  v6092 = (v6093 & i22) | (v5869 & ~i22),
  v6093 = (v4514 & i23) | (v6094 & ~i23),
  v6094 = (v4514 & i24) | (v6095 & ~i24),
  v6095 = (v6097 & i29) | (v6096 & ~i29),
  v6096 = (v5866 & i30) | (v4266 & ~i30),
  v6097 = (v5866 & i30) | (v4516 & ~i30),
  v6098 = (v5862 & i13) | (v6099 & ~i13),
  v6099 = (v6117 & i14) | (v6100 & ~i14),
  v6100 = (v6106 & i21) | (v6101 & ~i21),
  v6101 = (v4932 & i23) | (v6102 & ~i23),
  v6102 = (v4932 & i24) | (v6103 & ~i24),
  v6103 = (v5865 & i26) | (v6104 & ~i26),
  v6104 = (v5865 & i27) | (v6105 & ~i27),
  v6105 = (v26 & i30) | (v27 & ~i30),
  v6106 = (v6112 & i22) | (v6107 & ~i22),
  v6107 = (v4938 & i23) | (v6108 & ~i23),
  v6108 = (v4938 & i24) | (v6109 & ~i24),
  v6109 = (v5871 & i26) | (v6110 & ~i26),
  v6110 = (v5871 & i27) | (v6111 & ~i27),
  v6111 = (v26 & i30) | (v3909 & ~i30),
  v6112 = (v4942 & i23) | (v6113 & ~i23),
  v6113 = (v4942 & i24) | (v6114 & ~i24),
  v6114 = (v5874 & i26) | (v6115 & ~i26),
  v6115 = (v5874 & i27) | (v6116 & ~i27),
  v6116 = (v26 & i30) | (v3913 & ~i30),
  v6117 = (v6121 & i21) | (v6118 & ~i21),
  v6118 = (v5138 & i23) | (v6119 & ~i23),
  v6119 = (v5138 & i24) | (v6120 & ~i24),
  v6120 = (v6105 & i27) | (v5865 & ~i27),
  v6121 = (v6125 & i22) | (v6122 & ~i22),
  v6122 = (v5140 & i23) | (v6123 & ~i23),
  v6123 = (v5140 & i24) | (v6124 & ~i24),
  v6124 = (v6111 & i27) | (v5871 & ~i27),
  v6125 = (v5142 & i23) | (v6126 & ~i23),
  v6126 = (v5142 & i24) | (v6127 & ~i24),
  v6127 = (v6116 & i27) | (v5874 & ~i27),
  v6128 = (v5862 & i12) | (v6129 & ~i12),
  v6129 = (v5862 & i13) | (v6130 & ~i13),
  v6130 = (v6131 & i14) | (v5862 & ~i14),
  v6131 = (v6135 & i21) | (v6132 & ~i21),
  v6132 = (v5283 & i23) | (v6133 & ~i23),
  v6133 = (v5283 & i24) | (v6134 & ~i24),
  v6134 = (v6104 & i26) | (v5865 & ~i26),
  v6135 = (v6139 & i22) | (v6136 & ~i22),
  v6136 = (v5285 & i23) | (v6137 & ~i23),
  v6137 = (v5285 & i24) | (v6138 & ~i24),
  v6138 = (v6110 & i26) | (v5871 & ~i26),
  v6139 = (v5287 & i23) | (v6140 & ~i23),
  v6140 = (v5287 & i24) | (v6141 & ~i24),
  v6141 = (v6115 & i26) | (v5874 & ~i26),
  v6142 = (v6274 & i11) | (v6143 & ~i11),
  v6143 = (v6262 & i12) | (v6144 & ~i12),
  v6144 = (v6146 & i13) | (v6145 & ~i13),
  v6145 = (v6151 & i14) | (v6146 & ~i14),
  v6146 = (v6148 & i21) | (v6147 & ~i21),
  v6147 = (v5865 & i24) | (v27 & ~i24),
  v6148 = (v6150 & i22) | (v6149 & ~i22),
  v6149 = (v5871 & i24) | (v3908 & ~i24),
  v6150 = (v5874 & i24) | (v3912 & ~i24),
  v6151 = (v6207 & i15) | (v6152 & ~i15),
  v6152 = (v6180 & i16) | (v6153 & ~i16),
  v6153 = (v6169 & i17) | (v6154 & ~i17),
  v6154 = (v6162 & i19) | (v6155 & ~i19),
  v6155 = (v6159 & i20) | (v6156 & ~i20),
  v6156 = (v6157 & i21) | (v6147 & ~i21),
  v6157 = (v6158 & i22) | (v6149 & ~i22),
  v6158 = (v5884 & i24) | (v4276 & ~i24),
  v6159 = (v6160 & i21) | (v6147 & ~i21),
  v6160 = (v6161 & i22) | (v6149 & ~i22),
  v6161 = (v5891 & i24) | (v4284 & ~i24),
  v6162 = (v6166 & i20) | (v6163 & ~i20),
  v6163 = (v6164 & i21) | (v6147 & ~i21),
  v6164 = (v6165 & i22) | (v6149 & ~i22),
  v6165 = (v5899 & i24) | (v4293 & ~i24),
  v6166 = (v6167 & i21) | (v6147 & ~i21),
  v6167 = (v6168 & i22) | (v6149 & ~i22),
  v6168 = (v5906 & i24) | (v4301 & ~i24),
  v6169 = (v6177 & i19) | (v6170 & ~i19),
  v6170 = (v6174 & i20) | (v6171 & ~i20),
  v6171 = (v6172 & i21) | (v6147 & ~i21),
  v6172 = (v6173 & i22) | (v6149 & ~i22),
  v6173 = (v5915 & i24) | (v4311 & ~i24),
  v6174 = (v6175 & i21) | (v6147 & ~i21),
  v6175 = (v6176 & i22) | (v6149 & ~i22),
  v6176 = (v5922 & i24) | (v4319 & ~i24),
  v6177 = (v6178 & i21) | (v6147 & ~i21),
  v6178 = (v6179 & i22) | (v6149 & ~i22),
  v6179 = (v5929 & i24) | (v4327 & ~i24),
  v6180 = (v6196 & i17) | (v6181 & ~i17),
  v6181 = (v6189 & i19) | (v6182 & ~i19),
  v6182 = (v6186 & i20) | (v6183 & ~i20),
  v6183 = (v6184 & i21) | (v6147 & ~i21),
  v6184 = (v6185 & i22) | (v6149 & ~i22),
  v6185 = (v5939 & i24) | (v4338 & ~i24),
  v6186 = (v6187 & i21) | (v6147 & ~i21),
  v6187 = (v6188 & i22) | (v6149 & ~i22),
  v6188 = (v5946 & i24) | (v4346 & ~i24),
  v6189 = (v6193 & i20) | (v6190 & ~i20),
  v6190 = (v6191 & i21) | (v6147 & ~i21),
  v6191 = (v6192 & i22) | (v6149 & ~i22),
  v6192 = (v5954 & i24) | (v4355 & ~i24),
  v6193 = (v6194 & i21) | (v6147 & ~i21),
  v6194 = (v6195 & i22) | (v6149 & ~i22),
  v6195 = (v5961 & i24) | (v4363 & ~i24),
  v6196 = (v6204 & i19) | (v6197 & ~i19),
  v6197 = (v6201 & i20) | (v6198 & ~i20),
  v6198 = (v6199 & i21) | (v6147 & ~i21),
  v6199 = (v6200 & i22) | (v6149 & ~i22),
  v6200 = (v5970 & i24) | (v4373 & ~i24),
  v6201 = (v6202 & i21) | (v6147 & ~i21),
  v6202 = (v6203 & i22) | (v6149 & ~i22),
  v6203 = (v5977 & i24) | (v4381 & ~i24),
  v6204 = (v6205 & i21) | (v6147 & ~i21),
  v6205 = (v6206 & i22) | (v6149 & ~i22),
  v6206 = (v5984 & i24) | (v4389 & ~i24),
  v6207 = (v6235 & i16) | (v6208 & ~i16),
  v6208 = (v6224 & i17) | (v6209 & ~i17),
  v6209 = (v6217 & i19) | (v6210 & ~i19),
  v6210 = (v6214 & i20) | (v6211 & ~i20),
  v6211 = (v6212 & i21) | (v6147 & ~i21),
  v6212 = (v6213 & i22) | (v6149 & ~i22),
  v6213 = (v5995 & i24) | (v4401 & ~i24),
  v6214 = (v6215 & i21) | (v6147 & ~i21),
  v6215 = (v6216 & i22) | (v6149 & ~i22),
  v6216 = (v6002 & i24) | (v4409 & ~i24),
  v6217 = (v6221 & i20) | (v6218 & ~i20),
  v6218 = (v6219 & i21) | (v6147 & ~i21),
  v6219 = (v6220 & i22) | (v6149 & ~i22),
  v6220 = (v6010 & i24) | (v4418 & ~i24),
  v6221 = (v6222 & i21) | (v6147 & ~i21),
  v6222 = (v6223 & i22) | (v6149 & ~i22),
  v6223 = (v6017 & i24) | (v4426 & ~i24),
  v6224 = (v6232 & i19) | (v6225 & ~i19),
  v6225 = (v6229 & i20) | (v6226 & ~i20),
  v6226 = (v6227 & i21) | (v6147 & ~i21),
  v6227 = (v6228 & i22) | (v6149 & ~i22),
  v6228 = (v6026 & i24) | (v4436 & ~i24),
  v6229 = (v6230 & i21) | (v6147 & ~i21),
  v6230 = (v6231 & i22) | (v6149 & ~i22),
  v6231 = (v6033 & i24) | (v4444 & ~i24),
  v6232 = (v6233 & i21) | (v6147 & ~i21),
  v6233 = (v6234 & i22) | (v6149 & ~i22),
  v6234 = (v6040 & i24) | (v4452 & ~i24),
  v6235 = (v6251 & i17) | (v6236 & ~i17),
  v6236 = (v6244 & i19) | (v6237 & ~i19),
  v6237 = (v6241 & i20) | (v6238 & ~i20),
  v6238 = (v6239 & i21) | (v6147 & ~i21),
  v6239 = (v6240 & i22) | (v6149 & ~i22),
  v6240 = (v6050 & i24) | (v4463 & ~i24),
  v6241 = (v6242 & i21) | (v6147 & ~i21),
  v6242 = (v6243 & i22) | (v6149 & ~i22),
  v6243 = (v6057 & i24) | (v4471 & ~i24),
  v6244 = (v6248 & i20) | (v6245 & ~i20),
  v6245 = (v6246 & i21) | (v6147 & ~i21),
  v6246 = (v6247 & i22) | (v6149 & ~i22),
  v6247 = (v6065 & i24) | (v4480 & ~i24),
  v6248 = (v6249 & i21) | (v6147 & ~i21),
  v6249 = (v6250 & i22) | (v6149 & ~i22),
  v6250 = (v6072 & i24) | (v4488 & ~i24),
  v6251 = (v6259 & i19) | (v6252 & ~i19),
  v6252 = (v6256 & i20) | (v6253 & ~i20),
  v6253 = (v6254 & i21) | (v6147 & ~i21),
  v6254 = (v6255 & i22) | (v6149 & ~i22),
  v6255 = (v6081 & i24) | (v4498 & ~i24),
  v6256 = (v6257 & i21) | (v6147 & ~i21),
  v6257 = (v6258 & i22) | (v6149 & ~i22),
  v6258 = (v6088 & i24) | (v4506 & ~i24),
  v6259 = (v6260 & i21) | (v6147 & ~i21),
  v6260 = (v6261 & i22) | (v6149 & ~i22),
  v6261 = (v6095 & i24) | (v4514 & ~i24),
  v6262 = (v6146 & i13) | (v6263 & ~i13),
  v6263 = (v6269 & i14) | (v6264 & ~i14),
  v6264 = (v6266 & i21) | (v6265 & ~i21),
  v6265 = (v6103 & i24) | (v4932 & ~i24),
  v6266 = (v6268 & i22) | (v6267 & ~i22),
  v6267 = (v6109 & i24) | (v4938 & ~i24),
  v6268 = (v6114 & i24) | (v4942 & ~i24),
  v6269 = (v6271 & i21) | (v6270 & ~i21),
  v6270 = (v6120 & i24) | (v5138 & ~i24),
  v6271 = (v6273 & i22) | (v6272 & ~i22),
  v6272 = (v6124 & i24) | (v5140 & ~i24),
  v6273 = (v6127 & i24) | (v5142 & ~i24),
  v6274 = (v6146 & i12) | (v6275 & ~i12),
  v6275 = (v6146 & i13) | (v6276 & ~i13),
  v6276 = (v6277 & i14) | (v6146 & ~i14),
  v6277 = (v6279 & i21) | (v6278 & ~i21),
  v6278 = (v6134 & i24) | (v5283 & ~i24),
  v6279 = (v6281 & i22) | (v6280 & ~i22),
  v6280 = (v6138 & i24) | (v5285 & ~i24),
  v6281 = (v6141 & i24) | (v5287 & ~i24),
  v6282 = (v5843 & i8) | (v6283 & ~i8),
  v6283 = (v5843 & i9) | (v6284 & ~i9),
  v6284 = (v6285 & i10) | (v5843 & ~i10),
  v6285 = (v6417 & i11) | (v6286 & ~i11),
  v6286 = (v6405 & i12) | (v6287 & ~i12),
  v6287 = (v6289 & i13) | (v6288 & ~i13),
  v6288 = (v6294 & i14) | (v6289 & ~i14),
  v6289 = (v6291 & i21) | (v6290 & ~i21),
  v6290 = (v5864 & i23) | (v27 & ~i23),
  v6291 = (v6293 & i22) | (v6292 & ~i22),
  v6292 = (v5870 & i23) | (v3908 & ~i23),
  v6293 = (v5873 & i23) | (v3912 & ~i23),
  v6294 = (v6350 & i15) | (v6295 & ~i15),
  v6295 = (v6323 & i16) | (v6296 & ~i16),
  v6296 = (v6312 & i17) | (v6297 & ~i17),
  v6297 = (v6305 & i19) | (v6298 & ~i19),
  v6298 = (v6302 & i20) | (v6299 & ~i20),
  v6299 = (v6300 & i21) | (v6290 & ~i21),
  v6300 = (v6301 & i22) | (v6292 & ~i22),
  v6301 = (v5883 & i23) | (v4276 & ~i23),
  v6302 = (v6303 & i21) | (v6290 & ~i21),
  v6303 = (v6304 & i22) | (v6292 & ~i22),
  v6304 = (v5890 & i23) | (v4284 & ~i23),
  v6305 = (v6309 & i20) | (v6306 & ~i20),
  v6306 = (v6307 & i21) | (v6290 & ~i21),
  v6307 = (v6308 & i22) | (v6292 & ~i22),
  v6308 = (v5898 & i23) | (v4293 & ~i23),
  v6309 = (v6310 & i21) | (v6290 & ~i21),
  v6310 = (v6311 & i22) | (v6292 & ~i22),
  v6311 = (v5905 & i23) | (v4301 & ~i23),
  v6312 = (v6320 & i19) | (v6313 & ~i19),
  v6313 = (v6317 & i20) | (v6314 & ~i20),
  v6314 = (v6315 & i21) | (v6290 & ~i21),
  v6315 = (v6316 & i22) | (v6292 & ~i22),
  v6316 = (v5914 & i23) | (v4311 & ~i23),
  v6317 = (v6318 & i21) | (v6290 & ~i21),
  v6318 = (v6319 & i22) | (v6292 & ~i22),
  v6319 = (v5921 & i23) | (v4319 & ~i23),
  v6320 = (v6321 & i21) | (v6290 & ~i21),
  v6321 = (v6322 & i22) | (v6292 & ~i22),
  v6322 = (v5928 & i23) | (v4327 & ~i23),
  v6323 = (v6339 & i17) | (v6324 & ~i17),
  v6324 = (v6332 & i19) | (v6325 & ~i19),
  v6325 = (v6329 & i20) | (v6326 & ~i20),
  v6326 = (v6327 & i21) | (v6290 & ~i21),
  v6327 = (v6328 & i22) | (v6292 & ~i22),
  v6328 = (v5938 & i23) | (v4338 & ~i23),
  v6329 = (v6330 & i21) | (v6290 & ~i21),
  v6330 = (v6331 & i22) | (v6292 & ~i22),
  v6331 = (v5945 & i23) | (v4346 & ~i23),
  v6332 = (v6336 & i20) | (v6333 & ~i20),
  v6333 = (v6334 & i21) | (v6290 & ~i21),
  v6334 = (v6335 & i22) | (v6292 & ~i22),
  v6335 = (v5953 & i23) | (v4355 & ~i23),
  v6336 = (v6337 & i21) | (v6290 & ~i21),
  v6337 = (v6338 & i22) | (v6292 & ~i22),
  v6338 = (v5960 & i23) | (v4363 & ~i23),
  v6339 = (v6347 & i19) | (v6340 & ~i19),
  v6340 = (v6344 & i20) | (v6341 & ~i20),
  v6341 = (v6342 & i21) | (v6290 & ~i21),
  v6342 = (v6343 & i22) | (v6292 & ~i22),
  v6343 = (v5969 & i23) | (v4373 & ~i23),
  v6344 = (v6345 & i21) | (v6290 & ~i21),
  v6345 = (v6346 & i22) | (v6292 & ~i22),
  v6346 = (v5976 & i23) | (v4381 & ~i23),
  v6347 = (v6348 & i21) | (v6290 & ~i21),
  v6348 = (v6349 & i22) | (v6292 & ~i22),
  v6349 = (v5983 & i23) | (v4389 & ~i23),
  v6350 = (v6378 & i16) | (v6351 & ~i16),
  v6351 = (v6367 & i17) | (v6352 & ~i17),
  v6352 = (v6360 & i19) | (v6353 & ~i19),
  v6353 = (v6357 & i20) | (v6354 & ~i20),
  v6354 = (v6355 & i21) | (v6290 & ~i21),
  v6355 = (v6356 & i22) | (v6292 & ~i22),
  v6356 = (v5994 & i23) | (v4401 & ~i23),
  v6357 = (v6358 & i21) | (v6290 & ~i21),
  v6358 = (v6359 & i22) | (v6292 & ~i22),
  v6359 = (v6001 & i23) | (v4409 & ~i23),
  v6360 = (v6364 & i20) | (v6361 & ~i20),
  v6361 = (v6362 & i21) | (v6290 & ~i21),
  v6362 = (v6363 & i22) | (v6292 & ~i22),
  v6363 = (v6009 & i23) | (v4418 & ~i23),
  v6364 = (v6365 & i21) | (v6290 & ~i21),
  v6365 = (v6366 & i22) | (v6292 & ~i22),
  v6366 = (v6016 & i23) | (v4426 & ~i23),
  v6367 = (v6375 & i19) | (v6368 & ~i19),
  v6368 = (v6372 & i20) | (v6369 & ~i20),
  v6369 = (v6370 & i21) | (v6290 & ~i21),
  v6370 = (v6371 & i22) | (v6292 & ~i22),
  v6371 = (v6025 & i23) | (v4436 & ~i23),
  v6372 = (v6373 & i21) | (v6290 & ~i21),
  v6373 = (v6374 & i22) | (v6292 & ~i22),
  v6374 = (v6032 & i23) | (v4444 & ~i23),
  v6375 = (v6376 & i21) | (v6290 & ~i21),
  v6376 = (v6377 & i22) | (v6292 & ~i22),
  v6377 = (v6039 & i23) | (v4452 & ~i23),
  v6378 = (v6394 & i17) | (v6379 & ~i17),
  v6379 = (v6387 & i19) | (v6380 & ~i19),
  v6380 = (v6384 & i20) | (v6381 & ~i20),
  v6381 = (v6382 & i21) | (v6290 & ~i21),
  v6382 = (v6383 & i22) | (v6292 & ~i22),
  v6383 = (v6049 & i23) | (v4463 & ~i23),
  v6384 = (v6385 & i21) | (v6290 & ~i21),
  v6385 = (v6386 & i22) | (v6292 & ~i22),
  v6386 = (v6056 & i23) | (v4471 & ~i23),
  v6387 = (v6391 & i20) | (v6388 & ~i20),
  v6388 = (v6389 & i21) | (v6290 & ~i21),
  v6389 = (v6390 & i22) | (v6292 & ~i22),
  v6390 = (v6064 & i23) | (v4480 & ~i23),
  v6391 = (v6392 & i21) | (v6290 & ~i21),
  v6392 = (v6393 & i22) | (v6292 & ~i22),
  v6393 = (v6071 & i23) | (v4488 & ~i23),
  v6394 = (v6402 & i19) | (v6395 & ~i19),
  v6395 = (v6399 & i20) | (v6396 & ~i20),
  v6396 = (v6397 & i21) | (v6290 & ~i21),
  v6397 = (v6398 & i22) | (v6292 & ~i22),
  v6398 = (v6080 & i23) | (v4498 & ~i23),
  v6399 = (v6400 & i21) | (v6290 & ~i21),
  v6400 = (v6401 & i22) | (v6292 & ~i22),
  v6401 = (v6087 & i23) | (v4506 & ~i23),
  v6402 = (v6403 & i21) | (v6290 & ~i21),
  v6403 = (v6404 & i22) | (v6292 & ~i22),
  v6404 = (v6094 & i23) | (v4514 & ~i23),
  v6405 = (v6289 & i13) | (v6406 & ~i13),
  v6406 = (v6412 & i14) | (v6407 & ~i14),
  v6407 = (v6409 & i21) | (v6408 & ~i21),
  v6408 = (v6102 & i23) | (v4932 & ~i23),
  v6409 = (v6411 & i22) | (v6410 & ~i22),
  v6410 = (v6108 & i23) | (v4938 & ~i23),
  v6411 = (v6113 & i23) | (v4942 & ~i23),
  v6412 = (v6414 & i21) | (v6413 & ~i21),
  v6413 = (v6119 & i23) | (v5138 & ~i23),
  v6414 = (v6416 & i22) | (v6415 & ~i22),
  v6415 = (v6123 & i23) | (v5140 & ~i23),
  v6416 = (v6126 & i23) | (v5142 & ~i23),
  v6417 = (v6289 & i12) | (v6418 & ~i12),
  v6418 = (v6289 & i13) | (v6419 & ~i13),
  v6419 = (v6420 & i14) | (v6289 & ~i14),
  v6420 = (v6422 & i21) | (v6421 & ~i21),
  v6421 = (v6133 & i23) | (v5283 & ~i23),
  v6422 = (v6424 & i22) | (v6423 & ~i22),
  v6423 = (v6137 & i23) | (v5285 & ~i23),
  v6424 = (v6140 & i23) | (v5287 & ~i23),
  v6425 = (v6430 & i2) | (v6426 & ~i2),
  v6426 = (v6430 & i3) | (v6427 & ~i3),
  v6427 = (v6431 & i21) | (v6428 & ~i21),
  v6428 = (v6430 & i30) | (v6429 & ~i30),
  v6429 = (~v27 & ~i31) | i31,
  v6430 = i31,
  v6431 = (v6432 & i22) | (v6428 & ~i22),
  v6432 = (v6430 & i30) | (v6433 & ~i30),
  v6433 = (~v6434 & ~i31) | i31,
  v6434 = (~v6435 & ~i32) | i32,
  v6435 = (v6436 & i37) | (v633 & ~i37),
  v6436 = (v633 & i38) | ~i38,
  v6437 = (v6456 & i2) | (v6438 & ~i2),
  v6438 = (v6456 & i3) | (v6439 & ~i3),
  v6439 = (v7431 & i4) | (v6440 & ~i4),
  v6440 = (v7431 & i5) | (v6441 & ~i5),
  v6441 = (v7431 & i6) | (v6442 & ~i6),
  v6442 = (v7342 & i7) | (v6443 & ~i7),
  v6443 = (v7342 & i8) | (v6444 & ~i8),
  v6444 = (v7342 & i9) | (v6445 & ~i9),
  v6445 = (v7032 & i10) | (v6446 & ~i10),
  v6446 = (v6450 & i11) | (v6447 & ~i11),
  v6447 = (v6450 & i12) | (v6448 & ~i12),
  v6448 = (v6450 & i13) | (v6449 & ~i13),
  v6449 = (v6781 & i14) | (v6450 & ~i14),
  v6450 = (v6664 & i15) | (v6451 & ~i15),
  v6451 = (v6563 & i16) | (v6452 & ~i16),
  v6452 = (v6522 & i17) | (v6453 & ~i17),
  v6453 = (v6490 & i19) | (v6454 & ~i19),
  v6454 = (v6476 & i20) | (v6455 & ~i20),
  v6455 = (v6457 & i21) | (v6456 & ~i21),
  v6456 = i30,
  v6457 = (v6458 & i22) | (v6456 & ~i22),
  v6458 = (v6465 & i25) | (v6459 & ~i25),
  v6459 = (~v6460 & ~i30) | i30,
  v6460 = (v6461 & ~i31) | i31,
  v6461 = (v6462 & ~i32) | i32,
  v6462 = (v6464 & i37) | (v6463 & ~i37),
  v6463 = (v669 & i42) | ~i42,
  v6464 = (v6463 & i38) | (v632 & ~i38),
  v6465 = (~v6466 & ~i30) | i30,
  v6466 = (v6467 & ~i31) | i31,
  v6467 = (v6468 & ~i32) | i32,
  v6468 = (v6475 & i36) | (v6469 & ~i36),
  v6469 = (v6474 & i37) | (v6470 & ~i37),
  v6470 = (v6472 & i38) | (v6471 & ~i38),
  v6471 = (v632 & i39) | (v6472 & ~i39),
  v6472 = (v6463 & i41) | (v6473 & ~i41),
  v6473 = (v669 & i42) | (v630 & ~i42),
  v6474 = (v6472 & i38) | (v632 & ~i38),
  v6475 = (v6474 & i37) | (v6472 & ~i37),
  v6476 = (v6477 & i21) | (v6456 & ~i21),
  v6477 = (v6478 & i22) | (v6456 & ~i22),
  v6478 = (v6479 & i25) | (v6459 & ~i25),
  v6479 = (~v6480 & ~i30) | i30,
  v6480 = (v6481 & ~i31) | i31,
  v6481 = (v6482 & ~i32) | i32,
  v6482 = (v6489 & i36) | (v6483 & ~i36),
  v6483 = (v6488 & i37) | (v6484 & ~i37),
  v6484 = (v6486 & i38) | (v6485 & ~i38),
  v6485 = (v6486 & i39) | (v632 & ~i39),
  v6486 = (v6463 & i41) | (v6487 & ~i41),
  v6487 = (v669 & i42) | (v650 & ~i42),
  v6488 = (v6486 & i38) | (v632 & ~i38),
  v6489 = (v6488 & i37) | (v6486 & ~i37),
  v6490 = (v6507 & i20) | (v6491 & ~i20),
  v6491 = (v6492 & i21) | (v6456 & ~i21),
  v6492 = (v6493 & i22) | (v6456 & ~i22),
  v6493 = (v6494 & i25) | (v6459 & ~i25),
  v6494 = (~v6495 & ~i30) | i30,
  v6495 = (v6496 & ~i31) | i31,
  v6496 = (v6497 & ~i32) | i32,
  v6497 = (v6503 & i35) | (v6498 & ~i35),
  v6498 = (v6502 & i36) | (v6499 & ~i36),
  v6499 = (v6500 & i38) | (v632 & ~i38),
  v6500 = (v6472 & i40) | (v6501 & ~i40),
  v6501 = (v6463 & i41) | (v669 & ~i41),
  v6502 = (v6499 & i37) | (v6500 & ~i37),
  v6503 = (v6502 & i36) | (v6504 & ~i36),
  v6504 = (v6499 & i37) | (v6505 & ~i37),
  v6505 = (v6500 & i38) | (v6506 & ~i38),
  v6506 = (v632 & i39) | (v6500 & ~i39),
  v6507 = (v6508 & i21) | (v6456 & ~i21),
  v6508 = (v6509 & i22) | (v6456 & ~i22),
  v6509 = (v6510 & i25) | (v6459 & ~i25),
  v6510 = (~v6511 & ~i30) | i30,
  v6511 = (v6512 & ~i31) | i31,
  v6512 = (v6513 & ~i32) | i32,
  v6513 = (v6518 & i35) | (v6514 & ~i35),
  v6514 = (v6517 & i36) | (v6515 & ~i36),
  v6515 = (v6516 & i38) | (v632 & ~i38),
  v6516 = (v6486 & i40) | (v6501 & ~i40),
  v6517 = (v6515 & i37) | (v6516 & ~i37),
  v6518 = (v6517 & i36) | (v6519 & ~i36),
  v6519 = (v6515 & i37) | (v6520 & ~i37),
  v6520 = (v6516 & i38) | (v6521 & ~i38),
  v6521 = (v6516 & i39) | (v632 & ~i39),
  v6522 = (v6554 & i19) | (v6523 & ~i19),
  v6523 = (v6539 & i20) | (v6524 & ~i20),
  v6524 = (v6525 & i21) | (v6456 & ~i21),
  v6525 = (v6526 & i22) | (v6456 & ~i22),
  v6526 = (v6527 & i25) | (v6459 & ~i25),
  v6527 = (~v6528 & ~i30) | i30,
  v6528 = (v6529 & ~i31) | i31,
  v6529 = (v6530 & ~i32) | i32,
  v6530 = (v6538 & i35) | (v6531 & ~i35),
  v6531 = (v6537 & i36) | (v6532 & ~i36),
  v6532 = (v6536 & i37) | (v6533 & ~i37),
  v6533 = (v6535 & i38) | (v6534 & ~i38),
  v6534 = (v632 & i39) | (v6535 & ~i39),
  v6535 = (v6501 & i40) | (v6472 & ~i40),
  v6536 = (v6535 & i38) | (v632 & ~i38),
  v6537 = (v6536 & i37) | (v6535 & ~i37),
  v6538 = (v6537 & i36) | (v6536 & ~i36),
  v6539 = (v6540 & i21) | (v6456 & ~i21),
  v6540 = (v6541 & i22) | (v6456 & ~i22),
  v6541 = (v6542 & i25) | (v6459 & ~i25),
  v6542 = (~v6543 & ~i30) | i30,
  v6543 = (v6544 & ~i31) | i31,
  v6544 = (v6545 & ~i32) | i32,
  v6545 = (v6553 & i35) | (v6546 & ~i35),
  v6546 = (v6552 & i36) | (v6547 & ~i36),
  v6547 = (v6551 & i37) | (v6548 & ~i37),
  v6548 = (v6550 & i38) | (v6549 & ~i38),
  v6549 = (v6550 & i39) | (v632 & ~i39),
  v6550 = (v6501 & i40) | (v6486 & ~i40),
  v6551 = (v6550 & i38) | (v632 & ~i38),
  v6552 = (v6551 & i37) | (v6550 & ~i37),
  v6553 = (v6552 & i36) | (v6551 & ~i36),
  v6554 = (v6555 & i21) | (v6456 & ~i21),
  v6555 = (v6556 & i22) | (v6456 & ~i22),
  v6556 = (v6557 & i25) | (v6459 & ~i25),
  v6557 = (~v6558 & ~i30) | i30,
  v6558 = (v6559 & ~i31) | i31,
  v6559 = (v6560 & ~i32) | i32,
  v6560 = (v6562 & i36) | (v6561 & ~i36),
  v6561 = (v6501 & i38) | (v632 & ~i38),
  v6562 = (v6561 & i37) | (v6501 & ~i37),
  v6563 = (v6623 & i17) | (v6564 & ~i17),
  v6564 = (v6592 & i19) | (v6565 & ~i19),
  v6565 = (v6579 & i20) | (v6566 & ~i20),
  v6566 = (v6567 & i21) | (v6456 & ~i21),
  v6567 = (v6568 & i22) | (v6456 & ~i22),
  v6568 = (v6569 & i25) | (v6459 & ~i25),
  v6569 = (~v6570 & ~i30) | i30,
  v6570 = (v6571 & ~i31) | i31,
  v6571 = (v6572 & ~i32) | i32,
  v6572 = (v6578 & i36) | (v6573 & ~i36),
  v6573 = (v6577 & i37) | (v6574 & ~i37),
  v6574 = (v6576 & i38) | (v6575 & ~i38),
  v6575 = (v632 & i39) | (v6576 & ~i39),
  v6576 = (v669 & i41) | (v6473 & ~i41),
  v6577 = (v6576 & i38) | (v632 & ~i38),
  v6578 = (v6577 & i37) | (v6576 & ~i37),
  v6579 = (v6580 & i21) | (v6456 & ~i21),
  v6580 = (v6581 & i22) | (v6456 & ~i22),
  v6581 = (v6582 & i25) | (v6459 & ~i25),
  v6582 = (~v6583 & ~i30) | i30,
  v6583 = (v6584 & ~i31) | i31,
  v6584 = (v6585 & ~i32) | i32,
  v6585 = (v6591 & i36) | (v6586 & ~i36),
  v6586 = (v6590 & i37) | (v6587 & ~i37),
  v6587 = (v6589 & i38) | (v6588 & ~i38),
  v6588 = (v6589 & i39) | (v632 & ~i39),
  v6589 = (v669 & i41) | (v6487 & ~i41),
  v6590 = (v6589 & i38) | (v632 & ~i38),
  v6591 = (v6590 & i37) | (v6589 & ~i37),
  v6592 = (v6608 & i20) | (v6593 & ~i20),
  v6593 = (v6594 & i21) | (v6456 & ~i21),
  v6594 = (v6595 & i22) | (v6456 & ~i22),
  v6595 = (v6596 & i25) | (v6459 & ~i25),
  v6596 = (~v6597 & ~i30) | i30,
  v6597 = (v6598 & ~i31) | i31,
  v6598 = (v6599 & ~i32) | i32,
  v6599 = (v6604 & i35) | (v6600 & ~i35),
  v6600 = (v6603 & i36) | (v6601 & ~i36),
  v6601 = (v6602 & i38) | (v632 & ~i38),
  v6602 = (v6576 & i40) | (v669 & ~i40),
  v6603 = (v6601 & i37) | (v6602 & ~i37),
  v6604 = (v6603 & i36) | (v6605 & ~i36),
  v6605 = (v6601 & i37) | (v6606 & ~i37),
  v6606 = (v6602 & i38) | (v6607 & ~i38),
  v6607 = (v632 & i39) | (v6602 & ~i39),
  v6608 = (v6609 & i21) | (v6456 & ~i21),
  v6609 = (v6610 & i22) | (v6456 & ~i22),
  v6610 = (v6611 & i25) | (v6459 & ~i25),
  v6611 = (~v6612 & ~i30) | i30,
  v6612 = (v6613 & ~i31) | i31,
  v6613 = (v6614 & ~i32) | i32,
  v6614 = (v6619 & i35) | (v6615 & ~i35),
  v6615 = (v6618 & i36) | (v6616 & ~i36),
  v6616 = (v6617 & i38) | (v632 & ~i38),
  v6617 = (v6589 & i40) | (v669 & ~i40),
  v6618 = (v6616 & i37) | (v6617 & ~i37),
  v6619 = (v6618 & i36) | (v6620 & ~i36),
  v6620 = (v6616 & i37) | (v6621 & ~i37),
  v6621 = (v6617 & i38) | (v6622 & ~i38),
  v6622 = (v6617 & i39) | (v632 & ~i39),
  v6623 = (v6655 & i19) | (v6624 & ~i19),
  v6624 = (v6640 & i20) | (v6625 & ~i20),
  v6625 = (v6626 & i21) | (v6456 & ~i21),
  v6626 = (v6627 & i22) | (v6456 & ~i22),
  v6627 = (v6628 & i25) | (v6459 & ~i25),
  v6628 = (~v6629 & ~i30) | i30,
  v6629 = (v6630 & ~i31) | i31,
  v6630 = (v6631 & ~i32) | i32,
  v6631 = (v6639 & i35) | (v6632 & ~i35),
  v6632 = (v6638 & i36) | (v6633 & ~i36),
  v6633 = (v6637 & i37) | (v6634 & ~i37),
  v6634 = (v6636 & i38) | (v6635 & ~i38),
  v6635 = (v632 & i39) | (v6636 & ~i39),
  v6636 = (v669 & i40) | (v6576 & ~i40),
  v6637 = (v6636 & i38) | (v632 & ~i38),
  v6638 = (v6637 & i37) | (v6636 & ~i37),
  v6639 = (v6638 & i36) | (v6637 & ~i36),
  v6640 = (v6641 & i21) | (v6456 & ~i21),
  v6641 = (v6642 & i22) | (v6456 & ~i22),
  v6642 = (v6643 & i25) | (v6459 & ~i25),
  v6643 = (~v6644 & ~i30) | i30,
  v6644 = (v6645 & ~i31) | i31,
  v6645 = (v6646 & ~i32) | i32,
  v6646 = (v6654 & i35) | (v6647 & ~i35),
  v6647 = (v6653 & i36) | (v6648 & ~i36),
  v6648 = (v6652 & i37) | (v6649 & ~i37),
  v6649 = (v6651 & i38) | (v6650 & ~i38),
  v6650 = (v6651 & i39) | (v632 & ~i39),
  v6651 = (v669 & i40) | (v6589 & ~i40),
  v6652 = (v6651 & i38) | (v632 & ~i38),
  v6653 = (v6652 & i37) | (v6651 & ~i37),
  v6654 = (v6653 & i36) | (v6652 & ~i36),
  v6655 = (v6656 & i21) | (v6456 & ~i21),
  v6656 = (v6657 & i22) | (v6456 & ~i22),
  v6657 = (v6658 & i25) | (v6459 & ~i25),
  v6658 = (~v6659 & ~i30) | i30,
  v6659 = (v6660 & ~i31) | i31,
  v6660 = (v6661 & ~i32) | i32,
  v6661 = (v6663 & i36) | (v6662 & ~i36),
  v6662 = (v669 & i38) | (v632 & ~i38),
  v6663 = (v6662 & i37) | (v669 & ~i37),
  v6664 = (v6723 & i16) | (v6665 & ~i16),
  v6665 = (v6699 & i17) | (v6666 & ~i17),
  v6666 = (v6682 & i19) | (v6667 & ~i19),
  v6667 = (v6675 & i20) | (v6668 & ~i20),
  v6668 = (v6669 & i21) | (v6456 & ~i21),
  v6669 = (v6670 & i22) | (v6456 & ~i22),
  v6670 = (v6671 & i25) | (v6459 & ~i25),
  v6671 = (~v6672 & ~i30) | i30,
  v6672 = (v6673 & ~i31) | i31,
  v6673 = (v6674 & ~i32) | i32,
  v6674 = (v6474 & i36) | (v6469 & ~i36),
  v6675 = (v6676 & i21) | (v6456 & ~i21),
  v6676 = (v6677 & i22) | (v6456 & ~i22),
  v6677 = (v6678 & i25) | (v6459 & ~i25),
  v6678 = (~v6679 & ~i30) | i30,
  v6679 = (v6680 & ~i31) | i31,
  v6680 = (v6681 & ~i32) | i32,
  v6681 = (v6488 & i36) | (v6483 & ~i36),
  v6682 = (v6691 & i20) | (v6683 & ~i20),
  v6683 = (v6684 & i21) | (v6456 & ~i21),
  v6684 = (v6685 & i22) | (v6456 & ~i22),
  v6685 = (v6686 & i25) | (v6459 & ~i25),
  v6686 = (~v6687 & ~i30) | i30,
  v6687 = (v6688 & ~i31) | i31,
  v6688 = (v6689 & ~i32) | i32,
  v6689 = (v6690 & i35) | (v6499 & ~i35),
  v6690 = (v6499 & i36) | (v6504 & ~i36),
  v6691 = (v6692 & i21) | (v6456 & ~i21),
  v6692 = (v6693 & i22) | (v6456 & ~i22),
  v6693 = (v6694 & i25) | (v6459 & ~i25),
  v6694 = (~v6695 & ~i30) | i30,
  v6695 = (v6696 & ~i31) | i31,
  v6696 = (v6697 & ~i32) | i32,
  v6697 = (v6698 & i35) | (v6515 & ~i35),
  v6698 = (v6515 & i36) | (v6519 & ~i36),
  v6699 = (v6717 & i19) | (v6700 & ~i19),
  v6700 = (v6709 & i20) | (v6701 & ~i20),
  v6701 = (v6702 & i21) | (v6456 & ~i21),
  v6702 = (v6703 & i22) | (v6456 & ~i22),
  v6703 = (v6704 & i25) | (v6459 & ~i25),
  v6704 = (~v6705 & ~i30) | i30,
  v6705 = (v6706 & ~i31) | i31,
  v6706 = (v6707 & ~i32) | i32,
  v6707 = (v6536 & i35) | (v6708 & ~i35),
  v6708 = (v6536 & i36) | (v6532 & ~i36),
  v6709 = (v6710 & i21) | (v6456 & ~i21),
  v6710 = (v6711 & i22) | (v6456 & ~i22),
  v6711 = (v6712 & i25) | (v6459 & ~i25),
  v6712 = (~v6713 & ~i30) | i30,
  v6713 = (v6714 & ~i31) | i31,
  v6714 = (v6715 & ~i32) | i32,
  v6715 = (v6551 & i35) | (v6716 & ~i35),
  v6716 = (v6551 & i36) | (v6547 & ~i36),
  v6717 = (v6718 & i21) | (v6456 & ~i21),
  v6718 = (v6719 & i22) | (v6456 & ~i22),
  v6719 = (v6720 & i25) | (v6459 & ~i25),
  v6720 = (~v6721 & ~i30) | i30,
  v6721 = (v6722 & ~i31) | i31,
  v6722 = (v6561 & ~i32) | i32,
  v6723 = (v6757 & i17) | (v6724 & ~i17),
  v6724 = (v6740 & i19) | (v6725 & ~i19),
  v6725 = (v6733 & i20) | (v6726 & ~i20),
  v6726 = (v6727 & i21) | (v6456 & ~i21),
  v6727 = (v6728 & i22) | (v6456 & ~i22),
  v6728 = (v6729 & i25) | (v6459 & ~i25),
  v6729 = (~v6730 & ~i30) | i30,
  v6730 = (v6731 & ~i31) | i31,
  v6731 = (v6732 & ~i32) | i32,
  v6732 = (v6577 & i36) | (v6573 & ~i36),
  v6733 = (v6734 & i21) | (v6456 & ~i21),
  v6734 = (v6735 & i22) | (v6456 & ~i22),
  v6735 = (v6736 & i25) | (v6459 & ~i25),
  v6736 = (~v6737 & ~i30) | i30,
  v6737 = (v6738 & ~i31) | i31,
  v6738 = (v6739 & ~i32) | i32,
  v6739 = (v6590 & i36) | (v6586 & ~i36),
  v6740 = (v6749 & i20) | (v6741 & ~i20),
  v6741 = (v6742 & i21) | (v6456 & ~i21),
  v6742 = (v6743 & i22) | (v6456 & ~i22),
  v6743 = (v6744 & i25) | (v6459 & ~i25),
  v6744 = (~v6745 & ~i30) | i30,
  v6745 = (v6746 & ~i31) | i31,
  v6746 = (v6747 & ~i32) | i32,
  v6747 = (v6748 & i35) | (v6601 & ~i35),
  v6748 = (v6601 & i36) | (v6605 & ~i36),
  v6749 = (v6750 & i21) | (v6456 & ~i21),
  v6750 = (v6751 & i22) | (v6456 & ~i22),
  v6751 = (v6752 & i25) | (v6459 & ~i25),
  v6752 = (~v6753 & ~i30) | i30,
  v6753 = (v6754 & ~i31) | i31,
  v6754 = (v6755 & ~i32) | i32,
  v6755 = (v6756 & i35) | (v6616 & ~i35),
  v6756 = (v6616 & i36) | (v6620 & ~i36),
  v6757 = (v6775 & i19) | (v6758 & ~i19),
  v6758 = (v6767 & i20) | (v6759 & ~i20),
  v6759 = (v6760 & i21) | (v6456 & ~i21),
  v6760 = (v6761 & i22) | (v6456 & ~i22),
  v6761 = (v6762 & i25) | (v6459 & ~i25),
  v6762 = (~v6763 & ~i30) | i30,
  v6763 = (v6764 & ~i31) | i31,
  v6764 = (v6765 & ~i32) | i32,
  v6765 = (v6637 & i35) | (v6766 & ~i35),
  v6766 = (v6637 & i36) | (v6633 & ~i36),
  v6767 = (v6768 & i21) | (v6456 & ~i21),
  v6768 = (v6769 & i22) | (v6456 & ~i22),
  v6769 = (v6770 & i25) | (v6459 & ~i25),
  v6770 = (~v6771 & ~i30) | i30,
  v6771 = (v6772 & ~i31) | i31,
  v6772 = (v6773 & ~i32) | i32,
  v6773 = (v6652 & i35) | (v6774 & ~i35),
  v6774 = (v6652 & i36) | (v6648 & ~i36),
  v6775 = (v6776 & i21) | (v6456 & ~i21),
  v6776 = (v6777 & i22) | (v6456 & ~i22),
  v6777 = (v6778 & i25) | (v6459 & ~i25),
  v6778 = (~v6779 & ~i30) | i30,
  v6779 = (v6780 & ~i31) | i31,
  v6780 = (v6662 & ~i32) | i32,
  v6781 = (v6907 & i15) | (v6782 & ~i15),
  v6782 = (v6845 & i16) | (v6783 & ~i16),
  v6783 = (v6819 & i17) | (v6784 & ~i17),
  v6784 = (v6802 & i19) | (v6785 & ~i19),
  v6785 = (v6794 & i20) | (v6786 & ~i20),
  v6786 = (v6787 & i21) | (v6456 & ~i21),
  v6787 = (v6788 & i22) | (v6456 & ~i22),
  v6788 = (v6465 & i25) | (v6789 & ~i25),
  v6789 = (v6790 & i29) | (v6465 & ~i29),
  v6790 = (~v6791 & ~i30) | i30,
  v6791 = (v6792 & ~i31) | i31,
  v6792 = (v6793 & ~i32) | i32,
  v6793 = (v6462 & i33) | (v6468 & ~i33),
  v6794 = (v6795 & i21) | (v6456 & ~i21),
  v6795 = (v6796 & i22) | (v6456 & ~i22),
  v6796 = (v6479 & i25) | (v6797 & ~i25),
  v6797 = (v6798 & i29) | (v6479 & ~i29),
  v6798 = (~v6799 & ~i30) | i30,
  v6799 = (v6800 & ~i31) | i31,
  v6800 = (v6801 & ~i32) | i32,
  v6801 = (v6462 & i33) | (v6482 & ~i33),
  v6802 = (v6811 & i20) | (v6803 & ~i20),
  v6803 = (v6804 & i21) | (v6456 & ~i21),
  v6804 = (v6805 & i22) | (v6456 & ~i22),
  v6805 = (v6494 & i25) | (v6806 & ~i25),
  v6806 = (v6807 & i29) | (v6494 & ~i29),
  v6807 = (~v6808 & ~i30) | i30,
  v6808 = (v6809 & ~i31) | i31,
  v6809 = (v6810 & ~i32) | i32,
  v6810 = (v6462 & i33) | (v6497 & ~i33),
  v6811 = (v6812 & i21) | (v6456 & ~i21),
  v6812 = (v6813 & i22) | (v6456 & ~i22),
  v6813 = (v6510 & i25) | (v6814 & ~i25),
  v6814 = (v6815 & i29) | (v6510 & ~i29),
  v6815 = (~v6816 & ~i30) | i30,
  v6816 = (v6817 & ~i31) | i31,
  v6817 = (v6818 & ~i32) | i32,
  v6818 = (v6462 & i33) | (v6513 & ~i33),
  v6819 = (v6837 & i19) | (v6820 & ~i19),
  v6820 = (v6829 & i20) | (v6821 & ~i20),
  v6821 = (v6822 & i21) | (v6456 & ~i21),
  v6822 = (v6823 & i22) | (v6456 & ~i22),
  v6823 = (v6527 & i25) | (v6824 & ~i25),
  v6824 = (v6825 & i29) | (v6527 & ~i29),
  v6825 = (~v6826 & ~i30) | i30,
  v6826 = (v6827 & ~i31) | i31,
  v6827 = (v6828 & ~i32) | i32,
  v6828 = (v6462 & i33) | (v6530 & ~i33),
  v6829 = (v6830 & i21) | (v6456 & ~i21),
  v6830 = (v6831 & i22) | (v6456 & ~i22),
  v6831 = (v6542 & i25) | (v6832 & ~i25),
  v6832 = (v6833 & i29) | (v6542 & ~i29),
  v6833 = (~v6834 & ~i30) | i30,
  v6834 = (v6835 & ~i31) | i31,
  v6835 = (v6836 & ~i32) | i32,
  v6836 = (v6462 & i33) | (v6545 & ~i33),
  v6837 = (v6838 & i21) | (v6456 & ~i21),
  v6838 = (v6839 & i22) | (v6456 & ~i22),
  v6839 = (v6557 & i25) | (v6840 & ~i25),
  v6840 = (v6841 & i29) | (v6557 & ~i29),
  v6841 = (~v6842 & ~i30) | i30,
  v6842 = (v6843 & ~i31) | i31,
  v6843 = (v6844 & ~i32) | i32,
  v6844 = (v6462 & i33) | (v6560 & ~i33),
  v6845 = (v6881 & i17) | (v6846 & ~i17),
  v6846 = (v6864 & i19) | (v6847 & ~i19),
  v6847 = (v6856 & i20) | (v6848 & ~i20),
  v6848 = (v6849 & i21) | (v6456 & ~i21),
  v6849 = (v6850 & i22) | (v6456 & ~i22),
  v6850 = (v6569 & i25) | (v6851 & ~i25),
  v6851 = (v6852 & i29) | (v6569 & ~i29),
  v6852 = (~v6853 & ~i30) | i30,
  v6853 = (v6854 & ~i31) | i31,
  v6854 = (v6855 & ~i32) | i32,
  v6855 = (v6462 & i33) | (v6572 & ~i33),
  v6856 = (v6857 & i21) | (v6456 & ~i21),
  v6857 = (v6858 & i22) | (v6456 & ~i22),
  v6858 = (v6582 & i25) | (v6859 & ~i25),
  v6859 = (v6860 & i29) | (v6582 & ~i29),
  v6860 = (~v6861 & ~i30) | i30,
  v6861 = (v6862 & ~i31) | i31,
  v6862 = (v6863 & ~i32) | i32,
  v6863 = (v6462 & i33) | (v6585 & ~i33),
  v6864 = (v6873 & i20) | (v6865 & ~i20),
  v6865 = (v6866 & i21) | (v6456 & ~i21),
  v6866 = (v6867 & i22) | (v6456 & ~i22),
  v6867 = (v6596 & i25) | (v6868 & ~i25),
  v6868 = (v6869 & i29) | (v6596 & ~i29),
  v6869 = (~v6870 & ~i30) | i30,
  v6870 = (v6871 & ~i31) | i31,
  v6871 = (v6872 & ~i32) | i32,
  v6872 = (v6462 & i33) | (v6599 & ~i33),
  v6873 = (v6874 & i21) | (v6456 & ~i21),
  v6874 = (v6875 & i22) | (v6456 & ~i22),
  v6875 = (v6611 & i25) | (v6876 & ~i25),
  v6876 = (v6877 & i29) | (v6611 & ~i29),
  v6877 = (~v6878 & ~i30) | i30,
  v6878 = (v6879 & ~i31) | i31,
  v6879 = (v6880 & ~i32) | i32,
  v6880 = (v6462 & i33) | (v6614 & ~i33),
  v6881 = (v6899 & i19) | (v6882 & ~i19),
  v6882 = (v6891 & i20) | (v6883 & ~i20),
  v6883 = (v6884 & i21) | (v6456 & ~i21),
  v6884 = (v6885 & i22) | (v6456 & ~i22),
  v6885 = (v6628 & i25) | (v6886 & ~i25),
  v6886 = (v6887 & i29) | (v6628 & ~i29),
  v6887 = (~v6888 & ~i30) | i30,
  v6888 = (v6889 & ~i31) | i31,
  v6889 = (v6890 & ~i32) | i32,
  v6890 = (v6462 & i33) | (v6631 & ~i33),
  v6891 = (v6892 & i21) | (v6456 & ~i21),
  v6892 = (v6893 & i22) | (v6456 & ~i22),
  v6893 = (v6643 & i25) | (v6894 & ~i25),
  v6894 = (v6895 & i29) | (v6643 & ~i29),
  v6895 = (~v6896 & ~i30) | i30,
  v6896 = (v6897 & ~i31) | i31,
  v6897 = (v6898 & ~i32) | i32,
  v6898 = (v6462 & i33) | (v6646 & ~i33),
  v6899 = (v6900 & i21) | (v6456 & ~i21),
  v6900 = (v6901 & i22) | (v6456 & ~i22),
  v6901 = (v6658 & i25) | (v6902 & ~i25),
  v6902 = (v6903 & i29) | (v6658 & ~i29),
  v6903 = (~v6904 & ~i30) | i30,
  v6904 = (v6905 & ~i31) | i31,
  v6905 = (v6906 & ~i32) | i32,
  v6906 = (v6462 & i33) | (v6661 & ~i33),
  v6907 = (v6970 & i16) | (v6908 & ~i16),
  v6908 = (v6944 & i17) | (v6909 & ~i17),
  v6909 = (v6927 & i19) | (v6910 & ~i19),
  v6910 = (v6919 & i20) | (v6911 & ~i20),
  v6911 = (v6912 & i21) | (v6456 & ~i21),
  v6912 = (v6913 & i22) | (v6456 & ~i22),
  v6913 = (v6671 & i25) | (v6914 & ~i25),
  v6914 = (v6915 & i29) | (v6671 & ~i29),
  v6915 = (~v6916 & ~i30) | i30,
  v6916 = (v6917 & ~i31) | i31,
  v6917 = (v6918 & ~i32) | i32,
  v6918 = (v6462 & i33) | (v6674 & ~i33),
  v6919 = (v6920 & i21) | (v6456 & ~i21),
  v6920 = (v6921 & i22) | (v6456 & ~i22),
  v6921 = (v6678 & i25) | (v6922 & ~i25),
  v6922 = (v6923 & i29) | (v6678 & ~i29),
  v6923 = (~v6924 & ~i30) | i30,
  v6924 = (v6925 & ~i31) | i31,
  v6925 = (v6926 & ~i32) | i32,
  v6926 = (v6462 & i33) | (v6681 & ~i33),
  v6927 = (v6936 & i20) | (v6928 & ~i20),
  v6928 = (v6929 & i21) | (v6456 & ~i21),
  v6929 = (v6930 & i22) | (v6456 & ~i22),
  v6930 = (v6686 & i25) | (v6931 & ~i25),
  v6931 = (v6932 & i29) | (v6686 & ~i29),
  v6932 = (~v6933 & ~i30) | i30,
  v6933 = (v6934 & ~i31) | i31,
  v6934 = (v6935 & ~i32) | i32,
  v6935 = (v6462 & i33) | (v6689 & ~i33),
  v6936 = (v6937 & i21) | (v6456 & ~i21),
  v6937 = (v6938 & i22) | (v6456 & ~i22),
  v6938 = (v6694 & i25) | (v6939 & ~i25),
  v6939 = (v6940 & i29) | (v6694 & ~i29),
  v6940 = (~v6941 & ~i30) | i30,
  v6941 = (v6942 & ~i31) | i31,
  v6942 = (v6943 & ~i32) | i32,
  v6943 = (v6462 & i33) | (v6697 & ~i33),
  v6944 = (v6962 & i19) | (v6945 & ~i19),
  v6945 = (v6954 & i20) | (v6946 & ~i20),
  v6946 = (v6947 & i21) | (v6456 & ~i21),
  v6947 = (v6948 & i22) | (v6456 & ~i22),
  v6948 = (v6704 & i25) | (v6949 & ~i25),
  v6949 = (v6950 & i29) | (v6704 & ~i29),
  v6950 = (~v6951 & ~i30) | i30,
  v6951 = (v6952 & ~i31) | i31,
  v6952 = (v6953 & ~i32) | i32,
  v6953 = (v6462 & i33) | (v6707 & ~i33),
  v6954 = (v6955 & i21) | (v6456 & ~i21),
  v6955 = (v6956 & i22) | (v6456 & ~i22),
  v6956 = (v6712 & i25) | (v6957 & ~i25),
  v6957 = (v6958 & i29) | (v6712 & ~i29),
  v6958 = (~v6959 & ~i30) | i30,
  v6959 = (v6960 & ~i31) | i31,
  v6960 = (v6961 & ~i32) | i32,
  v6961 = (v6462 & i33) | (v6715 & ~i33),
  v6962 = (v6963 & i21) | (v6456 & ~i21),
  v6963 = (v6964 & i22) | (v6456 & ~i22),
  v6964 = (v6720 & i25) | (v6965 & ~i25),
  v6965 = (v6966 & i29) | (v6720 & ~i29),
  v6966 = (~v6967 & ~i30) | i30,
  v6967 = (v6968 & ~i31) | i31,
  v6968 = (v6969 & ~i32) | i32,
  v6969 = (v6462 & i33) | (v6561 & ~i33),
  v6970 = (v7006 & i17) | (v6971 & ~i17),
  v6971 = (v6989 & i19) | (v6972 & ~i19),
  v6972 = (v6981 & i20) | (v6973 & ~i20),
  v6973 = (v6974 & i21) | (v6456 & ~i21),
  v6974 = (v6975 & i22) | (v6456 & ~i22),
  v6975 = (v6729 & i25) | (v6976 & ~i25),
  v6976 = (v6977 & i29) | (v6729 & ~i29),
  v6977 = (~v6978 & ~i30) | i30,
  v6978 = (v6979 & ~i31) | i31,
  v6979 = (v6980 & ~i32) | i32,
  v6980 = (v6462 & i33) | (v6732 & ~i33),
  v6981 = (v6982 & i21) | (v6456 & ~i21),
  v6982 = (v6983 & i22) | (v6456 & ~i22),
  v6983 = (v6736 & i25) | (v6984 & ~i25),
  v6984 = (v6985 & i29) | (v6736 & ~i29),
  v6985 = (~v6986 & ~i30) | i30,
  v6986 = (v6987 & ~i31) | i31,
  v6987 = (v6988 & ~i32) | i32,
  v6988 = (v6462 & i33) | (v6739 & ~i33),
  v6989 = (v6998 & i20) | (v6990 & ~i20),
  v6990 = (v6991 & i21) | (v6456 & ~i21),
  v6991 = (v6992 & i22) | (v6456 & ~i22),
  v6992 = (v6744 & i25) | (v6993 & ~i25),
  v6993 = (v6994 & i29) | (v6744 & ~i29),
  v6994 = (~v6995 & ~i30) | i30,
  v6995 = (v6996 & ~i31) | i31,
  v6996 = (v6997 & ~i32) | i32,
  v6997 = (v6462 & i33) | (v6747 & ~i33),
  v6998 = (v6999 & i21) | (v6456 & ~i21),
  v6999 = (v7000 & i22) | (v6456 & ~i22),
  v7000 = (v6752 & i25) | (v7001 & ~i25),
  v7001 = (v7002 & i29) | (v6752 & ~i29),
  v7002 = (~v7003 & ~i30) | i30,
  v7003 = (v7004 & ~i31) | i31,
  v7004 = (v7005 & ~i32) | i32,
  v7005 = (v6462 & i33) | (v6755 & ~i33),
  v7006 = (v7024 & i19) | (v7007 & ~i19),
  v7007 = (v7016 & i20) | (v7008 & ~i20),
  v7008 = (v7009 & i21) | (v6456 & ~i21),
  v7009 = (v7010 & i22) | (v6456 & ~i22),
  v7010 = (v6762 & i25) | (v7011 & ~i25),
  v7011 = (v7012 & i29) | (v6762 & ~i29),
  v7012 = (~v7013 & ~i30) | i30,
  v7013 = (v7014 & ~i31) | i31,
  v7014 = (v7015 & ~i32) | i32,
  v7015 = (v6462 & i33) | (v6765 & ~i33),
  v7016 = (v7017 & i21) | (v6456 & ~i21),
  v7017 = (v7018 & i22) | (v6456 & ~i22),
  v7018 = (v6770 & i25) | (v7019 & ~i25),
  v7019 = (v7020 & i29) | (v6770 & ~i29),
  v7020 = (~v7021 & ~i30) | i30,
  v7021 = (v7022 & ~i31) | i31,
  v7022 = (v7023 & ~i32) | i32,
  v7023 = (v6462 & i33) | (v6773 & ~i33),
  v7024 = (v7025 & i21) | (v6456 & ~i21),
  v7025 = (v7026 & i22) | (v6456 & ~i22),
  v7026 = (v6778 & i25) | (v7027 & ~i25),
  v7027 = (v7028 & i29) | (v6778 & ~i29),
  v7028 = (~v7029 & ~i30) | i30,
  v7029 = (v7030 & ~i31) | i31,
  v7030 = (v7031 & ~i32) | i32,
  v7031 = (v6462 & i33) | (v6662 & ~i33),
  v7032 = (v7036 & i11) | (v7033 & ~i11),
  v7033 = (v7036 & i12) | (v7034 & ~i12),
  v7034 = (v7036 & i13) | (v7035 & ~i13),
  v7035 = (v7259 & i14) | (v7036 & ~i14),
  v7036 = (v7148 & i15) | (v7037 & ~i15),
  v7037 = (v7093 & i16) | (v7038 & ~i16),
  v7038 = (v7070 & i17) | (v7039 & ~i17),
  v7039 = (v7055 & i19) | (v7040 & ~i19),
  v7040 = (v7048 & i20) | (v7041 & ~i20),
  v7041 = (v7042 & i21) | (v6456 & ~i21),
  v7042 = (v7043 & i22) | (v6456 & ~i22),
  v7043 = (v7044 & i29) | (v6465 & ~i29),
  v7044 = (~v7045 & ~i30) | i30,
  v7045 = (v7046 & ~i31) | i31,
  v7046 = (v7047 & ~i32) | i32,
  v7047 = (v6468 & i33) | (v6462 & ~i33),
  v7048 = (v7049 & i21) | (v6456 & ~i21),
  v7049 = (v7050 & i22) | (v6456 & ~i22),
  v7050 = (v7051 & i29) | (v6479 & ~i29),
  v7051 = (~v7052 & ~i30) | i30,
  v7052 = (v7053 & ~i31) | i31,
  v7053 = (v7054 & ~i32) | i32,
  v7054 = (v6482 & i33) | (v6462 & ~i33),
  v7055 = (v7063 & i20) | (v7056 & ~i20),
  v7056 = (v7057 & i21) | (v6456 & ~i21),
  v7057 = (v7058 & i22) | (v6456 & ~i22),
  v7058 = (v7059 & i29) | (v6494 & ~i29),
  v7059 = (~v7060 & ~i30) | i30,
  v7060 = (v7061 & ~i31) | i31,
  v7061 = (v7062 & ~i32) | i32,
  v7062 = (v6497 & i33) | (v6462 & ~i33),
  v7063 = (v7064 & i21) | (v6456 & ~i21),
  v7064 = (v7065 & i22) | (v6456 & ~i22),
  v7065 = (v7066 & i29) | (v6510 & ~i29),
  v7066 = (~v7067 & ~i30) | i30,
  v7067 = (v7068 & ~i31) | i31,
  v7068 = (v7069 & ~i32) | i32,
  v7069 = (v6513 & i33) | (v6462 & ~i33),
  v7070 = (v7086 & i19) | (v7071 & ~i19),
  v7071 = (v7079 & i20) | (v7072 & ~i20),
  v7072 = (v7073 & i21) | (v6456 & ~i21),
  v7073 = (v7074 & i22) | (v6456 & ~i22),
  v7074 = (v7075 & i29) | (v6527 & ~i29),
  v7075 = (~v7076 & ~i30) | i30,
  v7076 = (v7077 & ~i31) | i31,
  v7077 = (v7078 & ~i32) | i32,
  v7078 = (v6530 & i33) | (v6462 & ~i33),
  v7079 = (v7080 & i21) | (v6456 & ~i21),
  v7080 = (v7081 & i22) | (v6456 & ~i22),
  v7081 = (v7082 & i29) | (v6542 & ~i29),
  v7082 = (~v7083 & ~i30) | i30,
  v7083 = (v7084 & ~i31) | i31,
  v7084 = (v7085 & ~i32) | i32,
  v7085 = (v6545 & i33) | (v6462 & ~i33),
  v7086 = (v7087 & i21) | (v6456 & ~i21),
  v7087 = (v7088 & i22) | (v6456 & ~i22),
  v7088 = (v7089 & i29) | (v6557 & ~i29),
  v7089 = (~v7090 & ~i30) | i30,
  v7090 = (v7091 & ~i31) | i31,
  v7091 = (v7092 & ~i32) | i32,
  v7092 = (v6560 & i33) | (v6462 & ~i33),
  v7093 = (v7125 & i17) | (v7094 & ~i17),
  v7094 = (v7110 & i19) | (v7095 & ~i19),
  v7095 = (v7103 & i20) | (v7096 & ~i20),
  v7096 = (v7097 & i21) | (v6456 & ~i21),
  v7097 = (v7098 & i22) | (v6456 & ~i22),
  v7098 = (v7099 & i29) | (v6569 & ~i29),
  v7099 = (~v7100 & ~i30) | i30,
  v7100 = (v7101 & ~i31) | i31,
  v7101 = (v7102 & ~i32) | i32,
  v7102 = (v6572 & i33) | (v6462 & ~i33),
  v7103 = (v7104 & i21) | (v6456 & ~i21),
  v7104 = (v7105 & i22) | (v6456 & ~i22),
  v7105 = (v7106 & i29) | (v6582 & ~i29),
  v7106 = (~v7107 & ~i30) | i30,
  v7107 = (v7108 & ~i31) | i31,
  v7108 = (v7109 & ~i32) | i32,
  v7109 = (v6585 & i33) | (v6462 & ~i33),
  v7110 = (v7118 & i20) | (v7111 & ~i20),
  v7111 = (v7112 & i21) | (v6456 & ~i21),
  v7112 = (v7113 & i22) | (v6456 & ~i22),
  v7113 = (v7114 & i29) | (v6596 & ~i29),
  v7114 = (~v7115 & ~i30) | i30,
  v7115 = (v7116 & ~i31) | i31,
  v7116 = (v7117 & ~i32) | i32,
  v7117 = (v6599 & i33) | (v6462 & ~i33),
  v7118 = (v7119 & i21) | (v6456 & ~i21),
  v7119 = (v7120 & i22) | (v6456 & ~i22),
  v7120 = (v7121 & i29) | (v6611 & ~i29),
  v7121 = (~v7122 & ~i30) | i30,
  v7122 = (v7123 & ~i31) | i31,
  v7123 = (v7124 & ~i32) | i32,
  v7124 = (v6614 & i33) | (v6462 & ~i33),
  v7125 = (v7141 & i19) | (v7126 & ~i19),
  v7126 = (v7134 & i20) | (v7127 & ~i20),
  v7127 = (v7128 & i21) | (v6456 & ~i21),
  v7128 = (v7129 & i22) | (v6456 & ~i22),
  v7129 = (v7130 & i29) | (v6628 & ~i29),
  v7130 = (~v7131 & ~i30) | i30,
  v7131 = (v7132 & ~i31) | i31,
  v7132 = (v7133 & ~i32) | i32,
  v7133 = (v6631 & i33) | (v6462 & ~i33),
  v7134 = (v7135 & i21) | (v6456 & ~i21),
  v7135 = (v7136 & i22) | (v6456 & ~i22),
  v7136 = (v7137 & i29) | (v6643 & ~i29),
  v7137 = (~v7138 & ~i30) | i30,
  v7138 = (v7139 & ~i31) | i31,
  v7139 = (v7140 & ~i32) | i32,
  v7140 = (v6646 & i33) | (v6462 & ~i33),
  v7141 = (v7142 & i21) | (v6456 & ~i21),
  v7142 = (v7143 & i22) | (v6456 & ~i22),
  v7143 = (v7144 & i29) | (v6658 & ~i29),
  v7144 = (~v7145 & ~i30) | i30,
  v7145 = (v7146 & ~i31) | i31,
  v7146 = (v7147 & ~i32) | i32,
  v7147 = (v6661 & i33) | (v6462 & ~i33),
  v7148 = (v7204 & i16) | (v7149 & ~i16),
  v7149 = (v7181 & i17) | (v7150 & ~i17),
  v7150 = (v7166 & i19) | (v7151 & ~i19),
  v7151 = (v7159 & i20) | (v7152 & ~i20),
  v7152 = (v7153 & i21) | (v6456 & ~i21),
  v7153 = (v7154 & i22) | (v6456 & ~i22),
  v7154 = (v7155 & i29) | (v6671 & ~i29),
  v7155 = (~v7156 & ~i30) | i30,
  v7156 = (v7157 & ~i31) | i31,
  v7157 = (v7158 & ~i32) | i32,
  v7158 = (v6674 & i33) | (v6462 & ~i33),
  v7159 = (v7160 & i21) | (v6456 & ~i21),
  v7160 = (v7161 & i22) | (v6456 & ~i22),
  v7161 = (v7162 & i29) | (v6678 & ~i29),
  v7162 = (~v7163 & ~i30) | i30,
  v7163 = (v7164 & ~i31) | i31,
  v7164 = (v7165 & ~i32) | i32,
  v7165 = (v6681 & i33) | (v6462 & ~i33),
  v7166 = (v7174 & i20) | (v7167 & ~i20),
  v7167 = (v7168 & i21) | (v6456 & ~i21),
  v7168 = (v7169 & i22) | (v6456 & ~i22),
  v7169 = (v7170 & i29) | (v6686 & ~i29),
  v7170 = (~v7171 & ~i30) | i30,
  v7171 = (v7172 & ~i31) | i31,
  v7172 = (v7173 & ~i32) | i32,
  v7173 = (v6689 & i33) | (v6462 & ~i33),
  v7174 = (v7175 & i21) | (v6456 & ~i21),
  v7175 = (v7176 & i22) | (v6456 & ~i22),
  v7176 = (v7177 & i29) | (v6694 & ~i29),
  v7177 = (~v7178 & ~i30) | i30,
  v7178 = (v7179 & ~i31) | i31,
  v7179 = (v7180 & ~i32) | i32,
  v7180 = (v6697 & i33) | (v6462 & ~i33),
  v7181 = (v7197 & i19) | (v7182 & ~i19),
  v7182 = (v7190 & i20) | (v7183 & ~i20),
  v7183 = (v7184 & i21) | (v6456 & ~i21),
  v7184 = (v7185 & i22) | (v6456 & ~i22),
  v7185 = (v7186 & i29) | (v6704 & ~i29),
  v7186 = (~v7187 & ~i30) | i30,
  v7187 = (v7188 & ~i31) | i31,
  v7188 = (v7189 & ~i32) | i32,
  v7189 = (v6707 & i33) | (v6462 & ~i33),
  v7190 = (v7191 & i21) | (v6456 & ~i21),
  v7191 = (v7192 & i22) | (v6456 & ~i22),
  v7192 = (v7193 & i29) | (v6712 & ~i29),
  v7193 = (~v7194 & ~i30) | i30,
  v7194 = (v7195 & ~i31) | i31,
  v7195 = (v7196 & ~i32) | i32,
  v7196 = (v6715 & i33) | (v6462 & ~i33),
  v7197 = (v7198 & i21) | (v6456 & ~i21),
  v7198 = (v7199 & i22) | (v6456 & ~i22),
  v7199 = (v7200 & i29) | (v6720 & ~i29),
  v7200 = (~v7201 & ~i30) | i30,
  v7201 = (v7202 & ~i31) | i31,
  v7202 = (v7203 & ~i32) | i32,
  v7203 = (v6561 & i33) | (v6462 & ~i33),
  v7204 = (v7236 & i17) | (v7205 & ~i17),
  v7205 = (v7221 & i19) | (v7206 & ~i19),
  v7206 = (v7214 & i20) | (v7207 & ~i20),
  v7207 = (v7208 & i21) | (v6456 & ~i21),
  v7208 = (v7209 & i22) | (v6456 & ~i22),
  v7209 = (v7210 & i29) | (v6729 & ~i29),
  v7210 = (~v7211 & ~i30) | i30,
  v7211 = (v7212 & ~i31) | i31,
  v7212 = (v7213 & ~i32) | i32,
  v7213 = (v6732 & i33) | (v6462 & ~i33),
  v7214 = (v7215 & i21) | (v6456 & ~i21),
  v7215 = (v7216 & i22) | (v6456 & ~i22),
  v7216 = (v7217 & i29) | (v6736 & ~i29),
  v7217 = (~v7218 & ~i30) | i30,
  v7218 = (v7219 & ~i31) | i31,
  v7219 = (v7220 & ~i32) | i32,
  v7220 = (v6739 & i33) | (v6462 & ~i33),
  v7221 = (v7229 & i20) | (v7222 & ~i20),
  v7222 = (v7223 & i21) | (v6456 & ~i21),
  v7223 = (v7224 & i22) | (v6456 & ~i22),
  v7224 = (v7225 & i29) | (v6744 & ~i29),
  v7225 = (~v7226 & ~i30) | i30,
  v7226 = (v7227 & ~i31) | i31,
  v7227 = (v7228 & ~i32) | i32,
  v7228 = (v6747 & i33) | (v6462 & ~i33),
  v7229 = (v7230 & i21) | (v6456 & ~i21),
  v7230 = (v7231 & i22) | (v6456 & ~i22),
  v7231 = (v7232 & i29) | (v6752 & ~i29),
  v7232 = (~v7233 & ~i30) | i30,
  v7233 = (v7234 & ~i31) | i31,
  v7234 = (v7235 & ~i32) | i32,
  v7235 = (v6755 & i33) | (v6462 & ~i33),
  v7236 = (v7252 & i19) | (v7237 & ~i19),
  v7237 = (v7245 & i20) | (v7238 & ~i20),
  v7238 = (v7239 & i21) | (v6456 & ~i21),
  v7239 = (v7240 & i22) | (v6456 & ~i22),
  v7240 = (v7241 & i29) | (v6762 & ~i29),
  v7241 = (~v7242 & ~i30) | i30,
  v7242 = (v7243 & ~i31) | i31,
  v7243 = (v7244 & ~i32) | i32,
  v7244 = (v6765 & i33) | (v6462 & ~i33),
  v7245 = (v7246 & i21) | (v6456 & ~i21),
  v7246 = (v7247 & i22) | (v6456 & ~i22),
  v7247 = (v7248 & i29) | (v6770 & ~i29),
  v7248 = (~v7249 & ~i30) | i30,
  v7249 = (v7250 & ~i31) | i31,
  v7250 = (v7251 & ~i32) | i32,
  v7251 = (v6773 & i33) | (v6462 & ~i33),
  v7252 = (v7253 & i21) | (v6456 & ~i21),
  v7253 = (v7254 & i22) | (v6456 & ~i22),
  v7254 = (v7255 & i29) | (v6778 & ~i29),
  v7255 = (~v7256 & ~i30) | i30,
  v7256 = (v7257 & ~i31) | i31,
  v7257 = (v7258 & ~i32) | i32,
  v7258 = (v6662 & i33) | (v6462 & ~i33),
  v7259 = (v7301 & i15) | (v7260 & ~i15),
  v7260 = (v7281 & i16) | (v7261 & ~i16),
  v7261 = (v7273 & i17) | (v7262 & ~i17),
  v7262 = (v7268 & i19) | (v7263 & ~i19),
  v7263 = (v7266 & i20) | (v7264 & ~i20),
  v7264 = (v7265 & i21) | (v6456 & ~i21),
  v7265 = (v6465 & i22) | (v6456 & ~i22),
  v7266 = (v7267 & i21) | (v6456 & ~i21),
  v7267 = (v6479 & i22) | (v6456 & ~i22),
  v7268 = (v7271 & i20) | (v7269 & ~i20),
  v7269 = (v7270 & i21) | (v6456 & ~i21),
  v7270 = (v6494 & i22) | (v6456 & ~i22),
  v7271 = (v7272 & i21) | (v6456 & ~i21),
  v7272 = (v6510 & i22) | (v6456 & ~i22),
  v7273 = (v7279 & i19) | (v7274 & ~i19),
  v7274 = (v7277 & i20) | (v7275 & ~i20),
  v7275 = (v7276 & i21) | (v6456 & ~i21),
  v7276 = (v6527 & i22) | (v6456 & ~i22),
  v7277 = (v7278 & i21) | (v6456 & ~i21),
  v7278 = (v6542 & i22) | (v6456 & ~i22),
  v7279 = (v7280 & i21) | (v6456 & ~i21),
  v7280 = (v6557 & i22) | (v6456 & ~i22),
  v7281 = (v7293 & i17) | (v7282 & ~i17),
  v7282 = (v7288 & i19) | (v7283 & ~i19),
  v7283 = (v7286 & i20) | (v7284 & ~i20),
  v7284 = (v7285 & i21) | (v6456 & ~i21),
  v7285 = (v6569 & i22) | (v6456 & ~i22),
  v7286 = (v7287 & i21) | (v6456 & ~i21),
  v7287 = (v6582 & i22) | (v6456 & ~i22),
  v7288 = (v7291 & i20) | (v7289 & ~i20),
  v7289 = (v7290 & i21) | (v6456 & ~i21),
  v7290 = (v6596 & i22) | (v6456 & ~i22),
  v7291 = (v7292 & i21) | (v6456 & ~i21),
  v7292 = (v6611 & i22) | (v6456 & ~i22),
  v7293 = (v7299 & i19) | (v7294 & ~i19),
  v7294 = (v7297 & i20) | (v7295 & ~i20),
  v7295 = (v7296 & i21) | (v6456 & ~i21),
  v7296 = (v6628 & i22) | (v6456 & ~i22),
  v7297 = (v7298 & i21) | (v6456 & ~i21),
  v7298 = (v6643 & i22) | (v6456 & ~i22),
  v7299 = (v7300 & i21) | (v6456 & ~i21),
  v7300 = (v6658 & i22) | (v6456 & ~i22),
  v7301 = (v7322 & i16) | (v7302 & ~i16),
  v7302 = (v7314 & i17) | (v7303 & ~i17),
  v7303 = (v7309 & i19) | (v7304 & ~i19),
  v7304 = (v7307 & i20) | (v7305 & ~i20),
  v7305 = (v7306 & i21) | (v6456 & ~i21),
  v7306 = (v6671 & i22) | (v6456 & ~i22),
  v7307 = (v7308 & i21) | (v6456 & ~i21),
  v7308 = (v6678 & i22) | (v6456 & ~i22),
  v7309 = (v7312 & i20) | (v7310 & ~i20),
  v7310 = (v7311 & i21) | (v6456 & ~i21),
  v7311 = (v6686 & i22) | (v6456 & ~i22),
  v7312 = (v7313 & i21) | (v6456 & ~i21),
  v7313 = (v6694 & i22) | (v6456 & ~i22),
  v7314 = (v7320 & i19) | (v7315 & ~i19),
  v7315 = (v7318 & i20) | (v7316 & ~i20),
  v7316 = (v7317 & i21) | (v6456 & ~i21),
  v7317 = (v6704 & i22) | (v6456 & ~i22),
  v7318 = (v7319 & i21) | (v6456 & ~i21),
  v7319 = (v6712 & i22) | (v6456 & ~i22),
  v7320 = (v7321 & i21) | (v6456 & ~i21),
  v7321 = (v6720 & i22) | (v6456 & ~i22),
  v7322 = (v7334 & i17) | (v7323 & ~i17),
  v7323 = (v7329 & i19) | (v7324 & ~i19),
  v7324 = (v7327 & i20) | (v7325 & ~i20),
  v7325 = (v7326 & i21) | (v6456 & ~i21),
  v7326 = (v6729 & i22) | (v6456 & ~i22),
  v7327 = (v7328 & i21) | (v6456 & ~i21),
  v7328 = (v6736 & i22) | (v6456 & ~i22),
  v7329 = (v7332 & i20) | (v7330 & ~i20),
  v7330 = (v7331 & i21) | (v6456 & ~i21),
  v7331 = (v6744 & i22) | (v6456 & ~i22),
  v7332 = (v7333 & i21) | (v6456 & ~i21),
  v7333 = (v6752 & i22) | (v6456 & ~i22),
  v7334 = (v7340 & i19) | (v7335 & ~i19),
  v7335 = (v7338 & i20) | (v7336 & ~i20),
  v7336 = (v7337 & i21) | (v6456 & ~i21),
  v7337 = (v6762 & i22) | (v6456 & ~i22),
  v7338 = (v7339 & i21) | (v6456 & ~i21),
  v7339 = (v6770 & i22) | (v6456 & ~i22),
  v7340 = (v7341 & i21) | (v6456 & ~i21),
  v7341 = (v6778 & i22) | (v6456 & ~i22),
  v7342 = (v7346 & i11) | (v7343 & ~i11),
  v7343 = (v7346 & i12) | (v7344 & ~i12),
  v7344 = (v7346 & i13) | (v7345 & ~i13),
  v7345 = (v7348 & i14) | (v7346 & ~i14),
  v7346 = (v7347 & i21) | (v6456 & ~i21),
  v7347 = (v6459 & i22) | (v6456 & ~i22),
  v7348 = (v7390 & i15) | (v7349 & ~i15),
  v7349 = (v7370 & i16) | (v7350 & ~i16),
  v7350 = (v7362 & i17) | (v7351 & ~i17),
  v7351 = (v7357 & i19) | (v7352 & ~i19),
  v7352 = (v7355 & i20) | (v7353 & ~i20),
  v7353 = (v7354 & i21) | (v6456 & ~i21),
  v7354 = (v6789 & i22) | (v6456 & ~i22),
  v7355 = (v7356 & i21) | (v6456 & ~i21),
  v7356 = (v6797 & i22) | (v6456 & ~i22),
  v7357 = (v7360 & i20) | (v7358 & ~i20),
  v7358 = (v7359 & i21) | (v6456 & ~i21),
  v7359 = (v6806 & i22) | (v6456 & ~i22),
  v7360 = (v7361 & i21) | (v6456 & ~i21),
  v7361 = (v6814 & i22) | (v6456 & ~i22),
  v7362 = (v7368 & i19) | (v7363 & ~i19),
  v7363 = (v7366 & i20) | (v7364 & ~i20),
  v7364 = (v7365 & i21) | (v6456 & ~i21),
  v7365 = (v6824 & i22) | (v6456 & ~i22),
  v7366 = (v7367 & i21) | (v6456 & ~i21),
  v7367 = (v6832 & i22) | (v6456 & ~i22),
  v7368 = (v7369 & i21) | (v6456 & ~i21),
  v7369 = (v6840 & i22) | (v6456 & ~i22),
  v7370 = (v7382 & i17) | (v7371 & ~i17),
  v7371 = (v7377 & i19) | (v7372 & ~i19),
  v7372 = (v7375 & i20) | (v7373 & ~i20),
  v7373 = (v7374 & i21) | (v6456 & ~i21),
  v7374 = (v6851 & i22) | (v6456 & ~i22),
  v7375 = (v7376 & i21) | (v6456 & ~i21),
  v7376 = (v6859 & i22) | (v6456 & ~i22),
  v7377 = (v7380 & i20) | (v7378 & ~i20),
  v7378 = (v7379 & i21) | (v6456 & ~i21),
  v7379 = (v6868 & i22) | (v6456 & ~i22),
  v7380 = (v7381 & i21) | (v6456 & ~i21),
  v7381 = (v6876 & i22) | (v6456 & ~i22),
  v7382 = (v7388 & i19) | (v7383 & ~i19),
  v7383 = (v7386 & i20) | (v7384 & ~i20),
  v7384 = (v7385 & i21) | (v6456 & ~i21),
  v7385 = (v6886 & i22) | (v6456 & ~i22),
  v7386 = (v7387 & i21) | (v6456 & ~i21),
  v7387 = (v6894 & i22) | (v6456 & ~i22),
  v7388 = (v7389 & i21) | (v6456 & ~i21),
  v7389 = (v6902 & i22) | (v6456 & ~i22),
  v7390 = (v7411 & i16) | (v7391 & ~i16),
  v7391 = (v7403 & i17) | (v7392 & ~i17),
  v7392 = (v7398 & i19) | (v7393 & ~i19),
  v7393 = (v7396 & i20) | (v7394 & ~i20),
  v7394 = (v7395 & i21) | (v6456 & ~i21),
  v7395 = (v6914 & i22) | (v6456 & ~i22),
  v7396 = (v7397 & i21) | (v6456 & ~i21),
  v7397 = (v6922 & i22) | (v6456 & ~i22),
  v7398 = (v7401 & i20) | (v7399 & ~i20),
  v7399 = (v7400 & i21) | (v6456 & ~i21),
  v7400 = (v6931 & i22) | (v6456 & ~i22),
  v7401 = (v7402 & i21) | (v6456 & ~i21),
  v7402 = (v6939 & i22) | (v6456 & ~i22),
  v7403 = (v7409 & i19) | (v7404 & ~i19),
  v7404 = (v7407 & i20) | (v7405 & ~i20),
  v7405 = (v7406 & i21) | (v6456 & ~i21),
  v7406 = (v6949 & i22) | (v6456 & ~i22),
  v7407 = (v7408 & i21) | (v6456 & ~i21),
  v7408 = (v6957 & i22) | (v6456 & ~i22),
  v7409 = (v7410 & i21) | (v6456 & ~i21),
  v7410 = (v6965 & i22) | (v6456 & ~i22),
  v7411 = (v7423 & i17) | (v7412 & ~i17),
  v7412 = (v7418 & i19) | (v7413 & ~i19),
  v7413 = (v7416 & i20) | (v7414 & ~i20),
  v7414 = (v7415 & i21) | (v6456 & ~i21),
  v7415 = (v6976 & i22) | (v6456 & ~i22),
  v7416 = (v7417 & i21) | (v6456 & ~i21),
  v7417 = (v6984 & i22) | (v6456 & ~i22),
  v7418 = (v7421 & i20) | (v7419 & ~i20),
  v7419 = (v7420 & i21) | (v6456 & ~i21),
  v7420 = (v6993 & i22) | (v6456 & ~i22),
  v7421 = (v7422 & i21) | (v6456 & ~i21),
  v7422 = (v7001 & i22) | (v6456 & ~i22),
  v7423 = (v7429 & i19) | (v7424 & ~i19),
  v7424 = (v7427 & i20) | (v7425 & ~i20),
  v7425 = (v7426 & i21) | (v6456 & ~i21),
  v7426 = (v7011 & i22) | (v6456 & ~i22),
  v7427 = (v7428 & i21) | (v6456 & ~i21),
  v7428 = (v7019 & i22) | (v6456 & ~i22),
  v7429 = (v7430 & i21) | (v6456 & ~i21),
  v7430 = (v7027 & i22) | (v6456 & ~i22),
  v7431 = (v8770 & i7) | (v7432 & ~i7),
  v7432 = (v8363 & i8) | (v7433 & ~i8),
  v7433 = (v8350 & i9) | (v7434 & ~i9),
  v7434 = (v7926 & i10) | (v7435 & ~i10),
  v7435 = (v7782 & i11) | (v7436 & ~i11),
  v7436 = (v7437 & i12) | (v6448 & ~i12),
  v7437 = (v6450 & i13) | (v7438 & ~i13),
  v7438 = (v7641 & i14) | (v7439 & ~i14),
  v7439 = (v7544 & i15) | (v7440 & ~i15),
  v7440 = (v7496 & i16) | (v7441 & ~i16),
  v7441 = (v7476 & i17) | (v7442 & ~i17),
  v7442 = (v7463 & i19) | (v7443 & ~i19),
  v7443 = (v7457 & i20) | (v7444 & ~i20),
  v7444 = (v7449 & i21) | (v7445 & ~i21),
  v7445 = (v6456 & i26) | (v7446 & ~i26),
  v7446 = (v6456 & i27) | (v7447 & ~i27),
  v7447 = v7448 & i30,
  v7448 = (~v63 & ~i31) | i31,
  v7449 = (v7450 & i22) | (v7445 & ~i22),
  v7450 = (v7454 & i25) | (v7451 & ~i25),
  v7451 = (v6459 & i26) | (v7452 & ~i26),
  v7452 = (v6459 & i27) | (v7453 & ~i27),
  v7453 = (v7448 & i30) | (~v6460 & ~i30),
  v7454 = (v6465 & i26) | (v7455 & ~i26),
  v7455 = (v6465 & i27) | (v7456 & ~i27),
  v7456 = (v7448 & i30) | (~v6466 & ~i30),
  v7457 = (v7458 & i21) | (v7445 & ~i21),
  v7458 = (v7459 & i22) | (v7445 & ~i22),
  v7459 = (v7460 & i25) | (v7451 & ~i25),
  v7460 = (v6479 & i26) | (v7461 & ~i26),
  v7461 = (v6479 & i27) | (v7462 & ~i27),
  v7462 = (v7448 & i30) | (~v6480 & ~i30),
  v7463 = (v7470 & i20) | (v7464 & ~i20),
  v7464 = (v7465 & i21) | (v7445 & ~i21),
  v7465 = (v7466 & i22) | (v7445 & ~i22),
  v7466 = (v7467 & i25) | (v7451 & ~i25),
  v7467 = (v6494 & i26) | (v7468 & ~i26),
  v7468 = (v6494 & i27) | (v7469 & ~i27),
  v7469 = (v7448 & i30) | (~v6495 & ~i30),
  v7470 = (v7471 & i21) | (v7445 & ~i21),
  v7471 = (v7472 & i22) | (v7445 & ~i22),
  v7472 = (v7473 & i25) | (v7451 & ~i25),
  v7473 = (v6510 & i26) | (v7474 & ~i26),
  v7474 = (v6510 & i27) | (v7475 & ~i27),
  v7475 = (v7448 & i30) | (~v6511 & ~i30),
  v7476 = (v7490 & i19) | (v7477 & ~i19),
  v7477 = (v7484 & i20) | (v7478 & ~i20),
  v7478 = (v7479 & i21) | (v7445 & ~i21),
  v7479 = (v7480 & i22) | (v7445 & ~i22),
  v7480 = (v7481 & i25) | (v7451 & ~i25),
  v7481 = (v6527 & i26) | (v7482 & ~i26),
  v7482 = (v6527 & i27) | (v7483 & ~i27),
  v7483 = (v7448 & i30) | (~v6528 & ~i30),
  v7484 = (v7485 & i21) | (v7445 & ~i21),
  v7485 = (v7486 & i22) | (v7445 & ~i22),
  v7486 = (v7487 & i25) | (v7451 & ~i25),
  v7487 = (v6542 & i26) | (v7488 & ~i26),
  v7488 = (v6542 & i27) | (v7489 & ~i27),
  v7489 = (v7448 & i30) | (~v6543 & ~i30),
  v7490 = (v7491 & i21) | (v7445 & ~i21),
  v7491 = (v7492 & i22) | (v7445 & ~i22),
  v7492 = (v7493 & i25) | (v7451 & ~i25),
  v7493 = (v6557 & i26) | (v7494 & ~i26),
  v7494 = (v6557 & i27) | (v7495 & ~i27),
  v7495 = (v7448 & i30) | (~v6558 & ~i30),
  v7496 = (v7524 & i17) | (v7497 & ~i17),
  v7497 = (v7511 & i19) | (v7498 & ~i19),
  v7498 = (v7505 & i20) | (v7499 & ~i20),
  v7499 = (v7500 & i21) | (v7445 & ~i21),
  v7500 = (v7501 & i22) | (v7445 & ~i22),
  v7501 = (v7502 & i25) | (v7451 & ~i25),
  v7502 = (v6569 & i26) | (v7503 & ~i26),
  v7503 = (v6569 & i27) | (v7504 & ~i27),
  v7504 = (v7448 & i30) | (~v6570 & ~i30),
  v7505 = (v7506 & i21) | (v7445 & ~i21),
  v7506 = (v7507 & i22) | (v7445 & ~i22),
  v7507 = (v7508 & i25) | (v7451 & ~i25),
  v7508 = (v6582 & i26) | (v7509 & ~i26),
  v7509 = (v6582 & i27) | (v7510 & ~i27),
  v7510 = (v7448 & i30) | (~v6583 & ~i30),
  v7511 = (v7518 & i20) | (v7512 & ~i20),
  v7512 = (v7513 & i21) | (v7445 & ~i21),
  v7513 = (v7514 & i22) | (v7445 & ~i22),
  v7514 = (v7515 & i25) | (v7451 & ~i25),
  v7515 = (v6596 & i26) | (v7516 & ~i26),
  v7516 = (v6596 & i27) | (v7517 & ~i27),
  v7517 = (v7448 & i30) | (~v6597 & ~i30),
  v7518 = (v7519 & i21) | (v7445 & ~i21),
  v7519 = (v7520 & i22) | (v7445 & ~i22),
  v7520 = (v7521 & i25) | (v7451 & ~i25),
  v7521 = (v6611 & i26) | (v7522 & ~i26),
  v7522 = (v6611 & i27) | (v7523 & ~i27),
  v7523 = (v7448 & i30) | (~v6612 & ~i30),
  v7524 = (v7538 & i19) | (v7525 & ~i19),
  v7525 = (v7532 & i20) | (v7526 & ~i20),
  v7526 = (v7527 & i21) | (v7445 & ~i21),
  v7527 = (v7528 & i22) | (v7445 & ~i22),
  v7528 = (v7529 & i25) | (v7451 & ~i25),
  v7529 = (v6628 & i26) | (v7530 & ~i26),
  v7530 = (v6628 & i27) | (v7531 & ~i27),
  v7531 = (v7448 & i30) | (~v6629 & ~i30),
  v7532 = (v7533 & i21) | (v7445 & ~i21),
  v7533 = (v7534 & i22) | (v7445 & ~i22),
  v7534 = (v7535 & i25) | (v7451 & ~i25),
  v7535 = (v6643 & i26) | (v7536 & ~i26),
  v7536 = (v6643 & i27) | (v7537 & ~i27),
  v7537 = (v7448 & i30) | (~v6644 & ~i30),
  v7538 = (v7539 & i21) | (v7445 & ~i21),
  v7539 = (v7540 & i22) | (v7445 & ~i22),
  v7540 = (v7541 & i25) | (v7451 & ~i25),
  v7541 = (v6658 & i26) | (v7542 & ~i26),
  v7542 = (v6658 & i27) | (v7543 & ~i27),
  v7543 = (v7448 & i30) | (~v6659 & ~i30),
  v7544 = (v7593 & i16) | (v7545 & ~i16),
  v7545 = (v7573 & i17) | (v7546 & ~i17),
  v7546 = (v7560 & i19) | (v7547 & ~i19),
  v7547 = (v7554 & i20) | (v7548 & ~i20),
  v7548 = (v7549 & i21) | (v7445 & ~i21),
  v7549 = (v7550 & i22) | (v7445 & ~i22),
  v7550 = (v7551 & i25) | (v7451 & ~i25),
  v7551 = (v6671 & i26) | (v7552 & ~i26),
  v7552 = (v6671 & i27) | (v7553 & ~i27),
  v7553 = (v7448 & i30) | (~v6672 & ~i30),
  v7554 = (v7555 & i21) | (v7445 & ~i21),
  v7555 = (v7556 & i22) | (v7445 & ~i22),
  v7556 = (v7557 & i25) | (v7451 & ~i25),
  v7557 = (v6678 & i26) | (v7558 & ~i26),
  v7558 = (v6678 & i27) | (v7559 & ~i27),
  v7559 = (v7448 & i30) | (~v6679 & ~i30),
  v7560 = (v7567 & i20) | (v7561 & ~i20),
  v7561 = (v7562 & i21) | (v7445 & ~i21),
  v7562 = (v7563 & i22) | (v7445 & ~i22),
  v7563 = (v7564 & i25) | (v7451 & ~i25),
  v7564 = (v6686 & i26) | (v7565 & ~i26),
  v7565 = (v6686 & i27) | (v7566 & ~i27),
  v7566 = (v7448 & i30) | (~v6687 & ~i30),
  v7567 = (v7568 & i21) | (v7445 & ~i21),
  v7568 = (v7569 & i22) | (v7445 & ~i22),
  v7569 = (v7570 & i25) | (v7451 & ~i25),
  v7570 = (v6694 & i26) | (v7571 & ~i26),
  v7571 = (v6694 & i27) | (v7572 & ~i27),
  v7572 = (v7448 & i30) | (~v6695 & ~i30),
  v7573 = (v7587 & i19) | (v7574 & ~i19),
  v7574 = (v7581 & i20) | (v7575 & ~i20),
  v7575 = (v7576 & i21) | (v7445 & ~i21),
  v7576 = (v7577 & i22) | (v7445 & ~i22),
  v7577 = (v7578 & i25) | (v7451 & ~i25),
  v7578 = (v6704 & i26) | (v7579 & ~i26),
  v7579 = (v6704 & i27) | (v7580 & ~i27),
  v7580 = (v7448 & i30) | (~v6705 & ~i30),
  v7581 = (v7582 & i21) | (v7445 & ~i21),
  v7582 = (v7583 & i22) | (v7445 & ~i22),
  v7583 = (v7584 & i25) | (v7451 & ~i25),
  v7584 = (v6712 & i26) | (v7585 & ~i26),
  v7585 = (v6712 & i27) | (v7586 & ~i27),
  v7586 = (v7448 & i30) | (~v6713 & ~i30),
  v7587 = (v7588 & i21) | (v7445 & ~i21),
  v7588 = (v7589 & i22) | (v7445 & ~i22),
  v7589 = (v7590 & i25) | (v7451 & ~i25),
  v7590 = (v6720 & i26) | (v7591 & ~i26),
  v7591 = (v6720 & i27) | (v7592 & ~i27),
  v7592 = (v7448 & i30) | (~v6721 & ~i30),
  v7593 = (v7621 & i17) | (v7594 & ~i17),
  v7594 = (v7608 & i19) | (v7595 & ~i19),
  v7595 = (v7602 & i20) | (v7596 & ~i20),
  v7596 = (v7597 & i21) | (v7445 & ~i21),
  v7597 = (v7598 & i22) | (v7445 & ~i22),
  v7598 = (v7599 & i25) | (v7451 & ~i25),
  v7599 = (v6729 & i26) | (v7600 & ~i26),
  v7600 = (v6729 & i27) | (v7601 & ~i27),
  v7601 = (v7448 & i30) | (~v6730 & ~i30),
  v7602 = (v7603 & i21) | (v7445 & ~i21),
  v7603 = (v7604 & i22) | (v7445 & ~i22),
  v7604 = (v7605 & i25) | (v7451 & ~i25),
  v7605 = (v6736 & i26) | (v7606 & ~i26),
  v7606 = (v6736 & i27) | (v7607 & ~i27),
  v7607 = (v7448 & i30) | (~v6737 & ~i30),
  v7608 = (v7615 & i20) | (v7609 & ~i20),
  v7609 = (v7610 & i21) | (v7445 & ~i21),
  v7610 = (v7611 & i22) | (v7445 & ~i22),
  v7611 = (v7612 & i25) | (v7451 & ~i25),
  v7612 = (v6744 & i26) | (v7613 & ~i26),
  v7613 = (v6744 & i27) | (v7614 & ~i27),
  v7614 = (v7448 & i30) | (~v6745 & ~i30),
  v7615 = (v7616 & i21) | (v7445 & ~i21),
  v7616 = (v7617 & i22) | (v7445 & ~i22),
  v7617 = (v7618 & i25) | (v7451 & ~i25),
  v7618 = (v6752 & i26) | (v7619 & ~i26),
  v7619 = (v6752 & i27) | (v7620 & ~i27),
  v7620 = (v7448 & i30) | (~v6753 & ~i30),
  v7621 = (v7635 & i19) | (v7622 & ~i19),
  v7622 = (v7629 & i20) | (v7623 & ~i20),
  v7623 = (v7624 & i21) | (v7445 & ~i21),
  v7624 = (v7625 & i22) | (v7445 & ~i22),
  v7625 = (v7626 & i25) | (v7451 & ~i25),
  v7626 = (v6762 & i26) | (v7627 & ~i26),
  v7627 = (v6762 & i27) | (v7628 & ~i27),
  v7628 = (v7448 & i30) | (~v6763 & ~i30),
  v7629 = (v7630 & i21) | (v7445 & ~i21),
  v7630 = (v7631 & i22) | (v7445 & ~i22),
  v7631 = (v7632 & i25) | (v7451 & ~i25),
  v7632 = (v6770 & i26) | (v7633 & ~i26),
  v7633 = (v6770 & i27) | (v7634 & ~i27),
  v7634 = (v7448 & i30) | (~v6771 & ~i30),
  v7635 = (v7636 & i21) | (v7445 & ~i21),
  v7636 = (v7637 & i22) | (v7445 & ~i22),
  v7637 = (v7638 & i25) | (v7451 & ~i25),
  v7638 = (v6778 & i26) | (v7639 & ~i26),
  v7639 = (v6778 & i27) | (v7640 & ~i27),
  v7640 = (v7448 & i30) | (~v6779 & ~i30),
  v7641 = (v7713 & i15) | (v7642 & ~i15),
  v7642 = (v7679 & i16) | (v7643 & ~i16),
  v7643 = (v7665 & i17) | (v7644 & ~i17),
  v7644 = (v7656 & i19) | (v7645 & ~i19),
  v7645 = (v7652 & i20) | (v7646 & ~i20),
  v7646 = (v7648 & i21) | (v7647 & ~i21),
  v7647 = (v7447 & i27) | (v6456 & ~i27),
  v7648 = (v7649 & i22) | (v7647 & ~i22),
  v7649 = (v7651 & i25) | (v7650 & ~i25),
  v7650 = (v7453 & i27) | (v6459 & ~i27),
  v7651 = (v7456 & i27) | (v6465 & ~i27),
  v7652 = (v7653 & i21) | (v7647 & ~i21),
  v7653 = (v7654 & i22) | (v7647 & ~i22),
  v7654 = (v7655 & i25) | (v7650 & ~i25),
  v7655 = (v7462 & i27) | (v6479 & ~i27),
  v7656 = (v7661 & i20) | (v7657 & ~i20),
  v7657 = (v7658 & i21) | (v7647 & ~i21),
  v7658 = (v7659 & i22) | (v7647 & ~i22),
  v7659 = (v7660 & i25) | (v7650 & ~i25),
  v7660 = (v7469 & i27) | (v6494 & ~i27),
  v7661 = (v7662 & i21) | (v7647 & ~i21),
  v7662 = (v7663 & i22) | (v7647 & ~i22),
  v7663 = (v7664 & i25) | (v7650 & ~i25),
  v7664 = (v7475 & i27) | (v6510 & ~i27),
  v7665 = (v7675 & i19) | (v7666 & ~i19),
  v7666 = (v7671 & i20) | (v7667 & ~i20),
  v7667 = (v7668 & i21) | (v7647 & ~i21),
  v7668 = (v7669 & i22) | (v7647 & ~i22),
  v7669 = (v7670 & i25) | (v7650 & ~i25),
  v7670 = (v7483 & i27) | (v6527 & ~i27),
  v7671 = (v7672 & i21) | (v7647 & ~i21),
  v7672 = (v7673 & i22) | (v7647 & ~i22),
  v7673 = (v7674 & i25) | (v7650 & ~i25),
  v7674 = (v7489 & i27) | (v6542 & ~i27),
  v7675 = (v7676 & i21) | (v7647 & ~i21),
  v7676 = (v7677 & i22) | (v7647 & ~i22),
  v7677 = (v7678 & i25) | (v7650 & ~i25),
  v7678 = (v7495 & i27) | (v6557 & ~i27),
  v7679 = (v7699 & i17) | (v7680 & ~i17),
  v7680 = (v7690 & i19) | (v7681 & ~i19),
  v7681 = (v7686 & i20) | (v7682 & ~i20),
  v7682 = (v7683 & i21) | (v7647 & ~i21),
  v7683 = (v7684 & i22) | (v7647 & ~i22),
  v7684 = (v7685 & i25) | (v7650 & ~i25),
  v7685 = (v7504 & i27) | (v6569 & ~i27),
  v7686 = (v7687 & i21) | (v7647 & ~i21),
  v7687 = (v7688 & i22) | (v7647 & ~i22),
  v7688 = (v7689 & i25) | (v7650 & ~i25),
  v7689 = (v7510 & i27) | (v6582 & ~i27),
  v7690 = (v7695 & i20) | (v7691 & ~i20),
  v7691 = (v7692 & i21) | (v7647 & ~i21),
  v7692 = (v7693 & i22) | (v7647 & ~i22),
  v7693 = (v7694 & i25) | (v7650 & ~i25),
  v7694 = (v7517 & i27) | (v6596 & ~i27),
  v7695 = (v7696 & i21) | (v7647 & ~i21),
  v7696 = (v7697 & i22) | (v7647 & ~i22),
  v7697 = (v7698 & i25) | (v7650 & ~i25),
  v7698 = (v7523 & i27) | (v6611 & ~i27),
  v7699 = (v7709 & i19) | (v7700 & ~i19),
  v7700 = (v7705 & i20) | (v7701 & ~i20),
  v7701 = (v7702 & i21) | (v7647 & ~i21),
  v7702 = (v7703 & i22) | (v7647 & ~i22),
  v7703 = (v7704 & i25) | (v7650 & ~i25),
  v7704 = (v7531 & i27) | (v6628 & ~i27),
  v7705 = (v7706 & i21) | (v7647 & ~i21),
  v7706 = (v7707 & i22) | (v7647 & ~i22),
  v7707 = (v7708 & i25) | (v7650 & ~i25),
  v7708 = (v7537 & i27) | (v6643 & ~i27),
  v7709 = (v7710 & i21) | (v7647 & ~i21),
  v7710 = (v7711 & i22) | (v7647 & ~i22),
  v7711 = (v7712 & i25) | (v7650 & ~i25),
  v7712 = (v7543 & i27) | (v6658 & ~i27),
  v7713 = (v7748 & i16) | (v7714 & ~i16),
  v7714 = (v7734 & i17) | (v7715 & ~i17),
  v7715 = (v7725 & i19) | (v7716 & ~i19),
  v7716 = (v7721 & i20) | (v7717 & ~i20),
  v7717 = (v7718 & i21) | (v7647 & ~i21),
  v7718 = (v7719 & i22) | (v7647 & ~i22),
  v7719 = (v7720 & i25) | (v7650 & ~i25),
  v7720 = (v7553 & i27) | (v6671 & ~i27),
  v7721 = (v7722 & i21) | (v7647 & ~i21),
  v7722 = (v7723 & i22) | (v7647 & ~i22),
  v7723 = (v7724 & i25) | (v7650 & ~i25),
  v7724 = (v7559 & i27) | (v6678 & ~i27),
  v7725 = (v7730 & i20) | (v7726 & ~i20),
  v7726 = (v7727 & i21) | (v7647 & ~i21),
  v7727 = (v7728 & i22) | (v7647 & ~i22),
  v7728 = (v7729 & i25) | (v7650 & ~i25),
  v7729 = (v7566 & i27) | (v6686 & ~i27),
  v7730 = (v7731 & i21) | (v7647 & ~i21),
  v7731 = (v7732 & i22) | (v7647 & ~i22),
  v7732 = (v7733 & i25) | (v7650 & ~i25),
  v7733 = (v7572 & i27) | (v6694 & ~i27),
  v7734 = (v7744 & i19) | (v7735 & ~i19),
  v7735 = (v7740 & i20) | (v7736 & ~i20),
  v7736 = (v7737 & i21) | (v7647 & ~i21),
  v7737 = (v7738 & i22) | (v7647 & ~i22),
  v7738 = (v7739 & i25) | (v7650 & ~i25),
  v7739 = (v7580 & i27) | (v6704 & ~i27),
  v7740 = (v7741 & i21) | (v7647 & ~i21),
  v7741 = (v7742 & i22) | (v7647 & ~i22),
  v7742 = (v7743 & i25) | (v7650 & ~i25),
  v7743 = (v7586 & i27) | (v6712 & ~i27),
  v7744 = (v7745 & i21) | (v7647 & ~i21),
  v7745 = (v7746 & i22) | (v7647 & ~i22),
  v7746 = (v7747 & i25) | (v7650 & ~i25),
  v7747 = (v7592 & i27) | (v6720 & ~i27),
  v7748 = (v7768 & i17) | (v7749 & ~i17),
  v7749 = (v7759 & i19) | (v7750 & ~i19),
  v7750 = (v7755 & i20) | (v7751 & ~i20),
  v7751 = (v7752 & i21) | (v7647 & ~i21),
  v7752 = (v7753 & i22) | (v7647 & ~i22),
  v7753 = (v7754 & i25) | (v7650 & ~i25),
  v7754 = (v7601 & i27) | (v6729 & ~i27),
  v7755 = (v7756 & i21) | (v7647 & ~i21),
  v7756 = (v7757 & i22) | (v7647 & ~i22),
  v7757 = (v7758 & i25) | (v7650 & ~i25),
  v7758 = (v7607 & i27) | (v6736 & ~i27),
  v7759 = (v7764 & i20) | (v7760 & ~i20),
  v7760 = (v7761 & i21) | (v7647 & ~i21),
  v7761 = (v7762 & i22) | (v7647 & ~i22),
  v7762 = (v7763 & i25) | (v7650 & ~i25),
  v7763 = (v7614 & i27) | (v6744 & ~i27),
  v7764 = (v7765 & i21) | (v7647 & ~i21),
  v7765 = (v7766 & i22) | (v7647 & ~i22),
  v7766 = (v7767 & i25) | (v7650 & ~i25),
  v7767 = (v7620 & i27) | (v6752 & ~i27),
  v7768 = (v7778 & i19) | (v7769 & ~i19),
  v7769 = (v7774 & i20) | (v7770 & ~i20),
  v7770 = (v7771 & i21) | (v7647 & ~i21),
  v7771 = (v7772 & i22) | (v7647 & ~i22),
  v7772 = (v7773 & i25) | (v7650 & ~i25),
  v7773 = (v7628 & i27) | (v6762 & ~i27),
  v7774 = (v7775 & i21) | (v7647 & ~i21),
  v7775 = (v7776 & i22) | (v7647 & ~i22),
  v7776 = (v7777 & i25) | (v7650 & ~i25),
  v7777 = (v7634 & i27) | (v6770 & ~i27),
  v7778 = (v7779 & i21) | (v7647 & ~i21),
  v7779 = (v7780 & i22) | (v7647 & ~i22),
  v7780 = (v7781 & i25) | (v7650 & ~i25),
  v7781 = (v7640 & i27) | (v6778 & ~i27),
  v7782 = (v6450 & i12) | (v7783 & ~i12),
  v7783 = (v6450 & i13) | (v7784 & ~i13),
  v7784 = (v7785 & i14) | (v6450 & ~i14),
  v7785 = (v7857 & i15) | (v7786 & ~i15),
  v7786 = (v7823 & i16) | (v7787 & ~i16),
  v7787 = (v7809 & i17) | (v7788 & ~i17),
  v7788 = (v7800 & i19) | (v7789 & ~i19),
  v7789 = (v7796 & i20) | (v7790 & ~i20),
  v7790 = (v7792 & i21) | (v7791 & ~i21),
  v7791 = (v7446 & i26) | (v6456 & ~i26),
  v7792 = (v7793 & i22) | (v7791 & ~i22),
  v7793 = (v7795 & i25) | (v7794 & ~i25),
  v7794 = (v7452 & i26) | (v6459 & ~i26),
  v7795 = (v7455 & i26) | (v6465 & ~i26),
  v7796 = (v7797 & i21) | (v7791 & ~i21),
  v7797 = (v7798 & i22) | (v7791 & ~i22),
  v7798 = (v7799 & i25) | (v7794 & ~i25),
  v7799 = (v7461 & i26) | (v6479 & ~i26),
  v7800 = (v7805 & i20) | (v7801 & ~i20),
  v7801 = (v7802 & i21) | (v7791 & ~i21),
  v7802 = (v7803 & i22) | (v7791 & ~i22),
  v7803 = (v7804 & i25) | (v7794 & ~i25),
  v7804 = (v7468 & i26) | (v6494 & ~i26),
  v7805 = (v7806 & i21) | (v7791 & ~i21),
  v7806 = (v7807 & i22) | (v7791 & ~i22),
  v7807 = (v7808 & i25) | (v7794 & ~i25),
  v7808 = (v7474 & i26) | (v6510 & ~i26),
  v7809 = (v7819 & i19) | (v7810 & ~i19),
  v7810 = (v7815 & i20) | (v7811 & ~i20),
  v7811 = (v7812 & i21) | (v7791 & ~i21),
  v7812 = (v7813 & i22) | (v7791 & ~i22),
  v7813 = (v7814 & i25) | (v7794 & ~i25),
  v7814 = (v7482 & i26) | (v6527 & ~i26),
  v7815 = (v7816 & i21) | (v7791 & ~i21),
  v7816 = (v7817 & i22) | (v7791 & ~i22),
  v7817 = (v7818 & i25) | (v7794 & ~i25),
  v7818 = (v7488 & i26) | (v6542 & ~i26),
  v7819 = (v7820 & i21) | (v7791 & ~i21),
  v7820 = (v7821 & i22) | (v7791 & ~i22),
  v7821 = (v7822 & i25) | (v7794 & ~i25),
  v7822 = (v7494 & i26) | (v6557 & ~i26),
  v7823 = (v7843 & i17) | (v7824 & ~i17),
  v7824 = (v7834 & i19) | (v7825 & ~i19),
  v7825 = (v7830 & i20) | (v7826 & ~i20),
  v7826 = (v7827 & i21) | (v7791 & ~i21),
  v7827 = (v7828 & i22) | (v7791 & ~i22),
  v7828 = (v7829 & i25) | (v7794 & ~i25),
  v7829 = (v7503 & i26) | (v6569 & ~i26),
  v7830 = (v7831 & i21) | (v7791 & ~i21),
  v7831 = (v7832 & i22) | (v7791 & ~i22),
  v7832 = (v7833 & i25) | (v7794 & ~i25),
  v7833 = (v7509 & i26) | (v6582 & ~i26),
  v7834 = (v7839 & i20) | (v7835 & ~i20),
  v7835 = (v7836 & i21) | (v7791 & ~i21),
  v7836 = (v7837 & i22) | (v7791 & ~i22),
  v7837 = (v7838 & i25) | (v7794 & ~i25),
  v7838 = (v7516 & i26) | (v6596 & ~i26),
  v7839 = (v7840 & i21) | (v7791 & ~i21),
  v7840 = (v7841 & i22) | (v7791 & ~i22),
  v7841 = (v7842 & i25) | (v7794 & ~i25),
  v7842 = (v7522 & i26) | (v6611 & ~i26),
  v7843 = (v7853 & i19) | (v7844 & ~i19),
  v7844 = (v7849 & i20) | (v7845 & ~i20),
  v7845 = (v7846 & i21) | (v7791 & ~i21),
  v7846 = (v7847 & i22) | (v7791 & ~i22),
  v7847 = (v7848 & i25) | (v7794 & ~i25),
  v7848 = (v7530 & i26) | (v6628 & ~i26),
  v7849 = (v7850 & i21) | (v7791 & ~i21),
  v7850 = (v7851 & i22) | (v7791 & ~i22),
  v7851 = (v7852 & i25) | (v7794 & ~i25),
  v7852 = (v7536 & i26) | (v6643 & ~i26),
  v7853 = (v7854 & i21) | (v7791 & ~i21),
  v7854 = (v7855 & i22) | (v7791 & ~i22),
  v7855 = (v7856 & i25) | (v7794 & ~i25),
  v7856 = (v7542 & i26) | (v6658 & ~i26),
  v7857 = (v7892 & i16) | (v7858 & ~i16),
  v7858 = (v7878 & i17) | (v7859 & ~i17),
  v7859 = (v7869 & i19) | (v7860 & ~i19),
  v7860 = (v7865 & i20) | (v7861 & ~i20),
  v7861 = (v7862 & i21) | (v7791 & ~i21),
  v7862 = (v7863 & i22) | (v7791 & ~i22),
  v7863 = (v7864 & i25) | (v7794 & ~i25),
  v7864 = (v7552 & i26) | (v6671 & ~i26),
  v7865 = (v7866 & i21) | (v7791 & ~i21),
  v7866 = (v7867 & i22) | (v7791 & ~i22),
  v7867 = (v7868 & i25) | (v7794 & ~i25),
  v7868 = (v7558 & i26) | (v6678 & ~i26),
  v7869 = (v7874 & i20) | (v7870 & ~i20),
  v7870 = (v7871 & i21) | (v7791 & ~i21),
  v7871 = (v7872 & i22) | (v7791 & ~i22),
  v7872 = (v7873 & i25) | (v7794 & ~i25),
  v7873 = (v7565 & i26) | (v6686 & ~i26),
  v7874 = (v7875 & i21) | (v7791 & ~i21),
  v7875 = (v7876 & i22) | (v7791 & ~i22),
  v7876 = (v7877 & i25) | (v7794 & ~i25),
  v7877 = (v7571 & i26) | (v6694 & ~i26),
  v7878 = (v7888 & i19) | (v7879 & ~i19),
  v7879 = (v7884 & i20) | (v7880 & ~i20),
  v7880 = (v7881 & i21) | (v7791 & ~i21),
  v7881 = (v7882 & i22) | (v7791 & ~i22),
  v7882 = (v7883 & i25) | (v7794 & ~i25),
  v7883 = (v7579 & i26) | (v6704 & ~i26),
  v7884 = (v7885 & i21) | (v7791 & ~i21),
  v7885 = (v7886 & i22) | (v7791 & ~i22),
  v7886 = (v7887 & i25) | (v7794 & ~i25),
  v7887 = (v7585 & i26) | (v6712 & ~i26),
  v7888 = (v7889 & i21) | (v7791 & ~i21),
  v7889 = (v7890 & i22) | (v7791 & ~i22),
  v7890 = (v7891 & i25) | (v7794 & ~i25),
  v7891 = (v7591 & i26) | (v6720 & ~i26),
  v7892 = (v7912 & i17) | (v7893 & ~i17),
  v7893 = (v7903 & i19) | (v7894 & ~i19),
  v7894 = (v7899 & i20) | (v7895 & ~i20),
  v7895 = (v7896 & i21) | (v7791 & ~i21),
  v7896 = (v7897 & i22) | (v7791 & ~i22),
  v7897 = (v7898 & i25) | (v7794 & ~i25),
  v7898 = (v7600 & i26) | (v6729 & ~i26),
  v7899 = (v7900 & i21) | (v7791 & ~i21),
  v7900 = (v7901 & i22) | (v7791 & ~i22),
  v7901 = (v7902 & i25) | (v7794 & ~i25),
  v7902 = (v7606 & i26) | (v6736 & ~i26),
  v7903 = (v7908 & i20) | (v7904 & ~i20),
  v7904 = (v7905 & i21) | (v7791 & ~i21),
  v7905 = (v7906 & i22) | (v7791 & ~i22),
  v7906 = (v7907 & i25) | (v7794 & ~i25),
  v7907 = (v7613 & i26) | (v6744 & ~i26),
  v7908 = (v7909 & i21) | (v7791 & ~i21),
  v7909 = (v7910 & i22) | (v7791 & ~i22),
  v7910 = (v7911 & i25) | (v7794 & ~i25),
  v7911 = (v7619 & i26) | (v6752 & ~i26),
  v7912 = (v7922 & i19) | (v7913 & ~i19),
  v7913 = (v7918 & i20) | (v7914 & ~i20),
  v7914 = (v7915 & i21) | (v7791 & ~i21),
  v7915 = (v7916 & i22) | (v7791 & ~i22),
  v7916 = (v7917 & i25) | (v7794 & ~i25),
  v7917 = (v7627 & i26) | (v6762 & ~i26),
  v7918 = (v7919 & i21) | (v7791 & ~i21),
  v7919 = (v7920 & i22) | (v7791 & ~i22),
  v7920 = (v7921 & i25) | (v7794 & ~i25),
  v7921 = (v7633 & i26) | (v6770 & ~i26),
  v7922 = (v7923 & i21) | (v7791 & ~i21),
  v7923 = (v7924 & i22) | (v7791 & ~i22),
  v7924 = (v7925 & i25) | (v7794 & ~i25),
  v7925 = (v7639 & i26) | (v6778 & ~i26),
  v7926 = (v8236 & i11) | (v7927 & ~i11),
  v7927 = (v7928 & i12) | (v7034 & ~i12),
  v7928 = (v7036 & i13) | (v7929 & ~i13),
  v7929 = (v8125 & i14) | (v7930 & ~i14),
  v7930 = (v8028 & i15) | (v7931 & ~i15),
  v7931 = (v7980 & i16) | (v7932 & ~i16),
  v7932 = (v7960 & i17) | (v7933 & ~i17),
  v7933 = (v7947 & i19) | (v7934 & ~i19),
  v7934 = (v7941 & i20) | (v7935 & ~i20),
  v7935 = (v7936 & i21) | (v7445 & ~i21),
  v7936 = (v7937 & i22) | (v7445 & ~i22),
  v7937 = (v7043 & i26) | (v7938 & ~i26),
  v7938 = (v7043 & i27) | (v7939 & ~i27),
  v7939 = (v7940 & i29) | (v7456 & ~i29),
  v7940 = (v7448 & i30) | (~v7045 & ~i30),
  v7941 = (v7942 & i21) | (v7445 & ~i21),
  v7942 = (v7943 & i22) | (v7445 & ~i22),
  v7943 = (v7050 & i26) | (v7944 & ~i26),
  v7944 = (v7050 & i27) | (v7945 & ~i27),
  v7945 = (v7946 & i29) | (v7462 & ~i29),
  v7946 = (v7448 & i30) | (~v7052 & ~i30),
  v7947 = (v7954 & i20) | (v7948 & ~i20),
  v7948 = (v7949 & i21) | (v7445 & ~i21),
  v7949 = (v7950 & i22) | (v7445 & ~i22),
  v7950 = (v7058 & i26) | (v7951 & ~i26),
  v7951 = (v7058 & i27) | (v7952 & ~i27),
  v7952 = (v7953 & i29) | (v7469 & ~i29),
  v7953 = (v7448 & i30) | (~v7060 & ~i30),
  v7954 = (v7955 & i21) | (v7445 & ~i21),
  v7955 = (v7956 & i22) | (v7445 & ~i22),
  v7956 = (v7065 & i26) | (v7957 & ~i26),
  v7957 = (v7065 & i27) | (v7958 & ~i27),
  v7958 = (v7959 & i29) | (v7475 & ~i29),
  v7959 = (v7448 & i30) | (~v7067 & ~i30),
  v7960 = (v7974 & i19) | (v7961 & ~i19),
  v7961 = (v7968 & i20) | (v7962 & ~i20),
  v7962 = (v7963 & i21) | (v7445 & ~i21),
  v7963 = (v7964 & i22) | (v7445 & ~i22),
  v7964 = (v7074 & i26) | (v7965 & ~i26),
  v7965 = (v7074 & i27) | (v7966 & ~i27),
  v7966 = (v7967 & i29) | (v7483 & ~i29),
  v7967 = (v7448 & i30) | (~v7076 & ~i30),
  v7968 = (v7969 & i21) | (v7445 & ~i21),
  v7969 = (v7970 & i22) | (v7445 & ~i22),
  v7970 = (v7081 & i26) | (v7971 & ~i26),
  v7971 = (v7081 & i27) | (v7972 & ~i27),
  v7972 = (v7973 & i29) | (v7489 & ~i29),
  v7973 = (v7448 & i30) | (~v7083 & ~i30),
  v7974 = (v7975 & i21) | (v7445 & ~i21),
  v7975 = (v7976 & i22) | (v7445 & ~i22),
  v7976 = (v7088 & i26) | (v7977 & ~i26),
  v7977 = (v7088 & i27) | (v7978 & ~i27),
  v7978 = (v7979 & i29) | (v7495 & ~i29),
  v7979 = (v7448 & i30) | (~v7090 & ~i30),
  v7980 = (v8008 & i17) | (v7981 & ~i17),
  v7981 = (v7995 & i19) | (v7982 & ~i19),
  v7982 = (v7989 & i20) | (v7983 & ~i20),
  v7983 = (v7984 & i21) | (v7445 & ~i21),
  v7984 = (v7985 & i22) | (v7445 & ~i22),
  v7985 = (v7098 & i26) | (v7986 & ~i26),
  v7986 = (v7098 & i27) | (v7987 & ~i27),
  v7987 = (v7988 & i29) | (v7504 & ~i29),
  v7988 = (v7448 & i30) | (~v7100 & ~i30),
  v7989 = (v7990 & i21) | (v7445 & ~i21),
  v7990 = (v7991 & i22) | (v7445 & ~i22),
  v7991 = (v7105 & i26) | (v7992 & ~i26),
  v7992 = (v7105 & i27) | (v7993 & ~i27),
  v7993 = (v7994 & i29) | (v7510 & ~i29),
  v7994 = (v7448 & i30) | (~v7107 & ~i30),
  v7995 = (v8002 & i20) | (v7996 & ~i20),
  v7996 = (v7997 & i21) | (v7445 & ~i21),
  v7997 = (v7998 & i22) | (v7445 & ~i22),
  v7998 = (v7113 & i26) | (v7999 & ~i26),
  v7999 = (v7113 & i27) | (v8000 & ~i27),
  v8000 = (v8001 & i29) | (v7517 & ~i29),
  v8001 = (v7448 & i30) | (~v7115 & ~i30),
  v8002 = (v8003 & i21) | (v7445 & ~i21),
  v8003 = (v8004 & i22) | (v7445 & ~i22),
  v8004 = (v7120 & i26) | (v8005 & ~i26),
  v8005 = (v7120 & i27) | (v8006 & ~i27),
  v8006 = (v8007 & i29) | (v7523 & ~i29),
  v8007 = (v7448 & i30) | (~v7122 & ~i30),
  v8008 = (v8022 & i19) | (v8009 & ~i19),
  v8009 = (v8016 & i20) | (v8010 & ~i20),
  v8010 = (v8011 & i21) | (v7445 & ~i21),
  v8011 = (v8012 & i22) | (v7445 & ~i22),
  v8012 = (v7129 & i26) | (v8013 & ~i26),
  v8013 = (v7129 & i27) | (v8014 & ~i27),
  v8014 = (v8015 & i29) | (v7531 & ~i29),
  v8015 = (v7448 & i30) | (~v7131 & ~i30),
  v8016 = (v8017 & i21) | (v7445 & ~i21),
  v8017 = (v8018 & i22) | (v7445 & ~i22),
  v8018 = (v7136 & i26) | (v8019 & ~i26),
  v8019 = (v7136 & i27) | (v8020 & ~i27),
  v8020 = (v8021 & i29) | (v7537 & ~i29),
  v8021 = (v7448 & i30) | (~v7138 & ~i30),
  v8022 = (v8023 & i21) | (v7445 & ~i21),
  v8023 = (v8024 & i22) | (v7445 & ~i22),
  v8024 = (v7143 & i26) | (v8025 & ~i26),
  v8025 = (v7143 & i27) | (v8026 & ~i27),
  v8026 = (v8027 & i29) | (v7543 & ~i29),
  v8027 = (v7448 & i30) | (~v7145 & ~i30),
  v8028 = (v8077 & i16) | (v8029 & ~i16),
  v8029 = (v8057 & i17) | (v8030 & ~i17),
  v8030 = (v8044 & i19) | (v8031 & ~i19),
  v8031 = (v8038 & i20) | (v8032 & ~i20),
  v8032 = (v8033 & i21) | (v7445 & ~i21),
  v8033 = (v8034 & i22) | (v7445 & ~i22),
  v8034 = (v7154 & i26) | (v8035 & ~i26),
  v8035 = (v7154 & i27) | (v8036 & ~i27),
  v8036 = (v8037 & i29) | (v7553 & ~i29),
  v8037 = (v7448 & i30) | (~v7156 & ~i30),
  v8038 = (v8039 & i21) | (v7445 & ~i21),
  v8039 = (v8040 & i22) | (v7445 & ~i22),
  v8040 = (v7161 & i26) | (v8041 & ~i26),
  v8041 = (v7161 & i27) | (v8042 & ~i27),
  v8042 = (v8043 & i29) | (v7559 & ~i29),
  v8043 = (v7448 & i30) | (~v7163 & ~i30),
  v8044 = (v8051 & i20) | (v8045 & ~i20),
  v8045 = (v8046 & i21) | (v7445 & ~i21),
  v8046 = (v8047 & i22) | (v7445 & ~i22),
  v8047 = (v7169 & i26) | (v8048 & ~i26),
  v8048 = (v7169 & i27) | (v8049 & ~i27),
  v8049 = (v8050 & i29) | (v7566 & ~i29),
  v8050 = (v7448 & i30) | (~v7171 & ~i30),
  v8051 = (v8052 & i21) | (v7445 & ~i21),
  v8052 = (v8053 & i22) | (v7445 & ~i22),
  v8053 = (v7176 & i26) | (v8054 & ~i26),
  v8054 = (v7176 & i27) | (v8055 & ~i27),
  v8055 = (v8056 & i29) | (v7572 & ~i29),
  v8056 = (v7448 & i30) | (~v7178 & ~i30),
  v8057 = (v8071 & i19) | (v8058 & ~i19),
  v8058 = (v8065 & i20) | (v8059 & ~i20),
  v8059 = (v8060 & i21) | (v7445 & ~i21),
  v8060 = (v8061 & i22) | (v7445 & ~i22),
  v8061 = (v7185 & i26) | (v8062 & ~i26),
  v8062 = (v7185 & i27) | (v8063 & ~i27),
  v8063 = (v8064 & i29) | (v7580 & ~i29),
  v8064 = (v7448 & i30) | (~v7187 & ~i30),
  v8065 = (v8066 & i21) | (v7445 & ~i21),
  v8066 = (v8067 & i22) | (v7445 & ~i22),
  v8067 = (v7192 & i26) | (v8068 & ~i26),
  v8068 = (v7192 & i27) | (v8069 & ~i27),
  v8069 = (v8070 & i29) | (v7586 & ~i29),
  v8070 = (v7448 & i30) | (~v7194 & ~i30),
  v8071 = (v8072 & i21) | (v7445 & ~i21),
  v8072 = (v8073 & i22) | (v7445 & ~i22),
  v8073 = (v7199 & i26) | (v8074 & ~i26),
  v8074 = (v7199 & i27) | (v8075 & ~i27),
  v8075 = (v8076 & i29) | (v7592 & ~i29),
  v8076 = (v7448 & i30) | (~v7201 & ~i30),
  v8077 = (v8105 & i17) | (v8078 & ~i17),
  v8078 = (v8092 & i19) | (v8079 & ~i19),
  v8079 = (v8086 & i20) | (v8080 & ~i20),
  v8080 = (v8081 & i21) | (v7445 & ~i21),
  v8081 = (v8082 & i22) | (v7445 & ~i22),
  v8082 = (v7209 & i26) | (v8083 & ~i26),
  v8083 = (v7209 & i27) | (v8084 & ~i27),
  v8084 = (v8085 & i29) | (v7601 & ~i29),
  v8085 = (v7448 & i30) | (~v7211 & ~i30),
  v8086 = (v8087 & i21) | (v7445 & ~i21),
  v8087 = (v8088 & i22) | (v7445 & ~i22),
  v8088 = (v7216 & i26) | (v8089 & ~i26),
  v8089 = (v7216 & i27) | (v8090 & ~i27),
  v8090 = (v8091 & i29) | (v7607 & ~i29),
  v8091 = (v7448 & i30) | (~v7218 & ~i30),
  v8092 = (v8099 & i20) | (v8093 & ~i20),
  v8093 = (v8094 & i21) | (v7445 & ~i21),
  v8094 = (v8095 & i22) | (v7445 & ~i22),
  v8095 = (v7224 & i26) | (v8096 & ~i26),
  v8096 = (v7224 & i27) | (v8097 & ~i27),
  v8097 = (v8098 & i29) | (v7614 & ~i29),
  v8098 = (v7448 & i30) | (~v7226 & ~i30),
  v8099 = (v8100 & i21) | (v7445 & ~i21),
  v8100 = (v8101 & i22) | (v7445 & ~i22),
  v8101 = (v7231 & i26) | (v8102 & ~i26),
  v8102 = (v7231 & i27) | (v8103 & ~i27),
  v8103 = (v8104 & i29) | (v7620 & ~i29),
  v8104 = (v7448 & i30) | (~v7233 & ~i30),
  v8105 = (v8119 & i19) | (v8106 & ~i19),
  v8106 = (v8113 & i20) | (v8107 & ~i20),
  v8107 = (v8108 & i21) | (v7445 & ~i21),
  v8108 = (v8109 & i22) | (v7445 & ~i22),
  v8109 = (v7240 & i26) | (v8110 & ~i26),
  v8110 = (v7240 & i27) | (v8111 & ~i27),
  v8111 = (v8112 & i29) | (v7628 & ~i29),
  v8112 = (v7448 & i30) | (~v7242 & ~i30),
  v8113 = (v8114 & i21) | (v7445 & ~i21),
  v8114 = (v8115 & i22) | (v7445 & ~i22),
  v8115 = (v7247 & i26) | (v8116 & ~i26),
  v8116 = (v7247 & i27) | (v8117 & ~i27),
  v8117 = (v8118 & i29) | (v7634 & ~i29),
  v8118 = (v7448 & i30) | (~v7249 & ~i30),
  v8119 = (v8120 & i21) | (v7445 & ~i21),
  v8120 = (v8121 & i22) | (v7445 & ~i22),
  v8121 = (v7254 & i26) | (v8122 & ~i26),
  v8122 = (v7254 & i27) | (v8123 & ~i27),
  v8123 = (v8124 & i29) | (v7640 & ~i29),
  v8124 = (v7448 & i30) | (~v7256 & ~i30),
  v8125 = (v8181 & i15) | (v8126 & ~i15),
  v8126 = (v8154 & i16) | (v8127 & ~i16),
  v8127 = (v8143 & i17) | (v8128 & ~i17),
  v8128 = (v8136 & i19) | (v8129 & ~i19),
  v8129 = (v8133 & i20) | (v8130 & ~i20),
  v8130 = (v8131 & i21) | (v7647 & ~i21),
  v8131 = (v8132 & i22) | (v7647 & ~i22),
  v8132 = (v7939 & i27) | (v7043 & ~i27),
  v8133 = (v8134 & i21) | (v7647 & ~i21),
  v8134 = (v8135 & i22) | (v7647 & ~i22),
  v8135 = (v7945 & i27) | (v7050 & ~i27),
  v8136 = (v8140 & i20) | (v8137 & ~i20),
  v8137 = (v8138 & i21) | (v7647 & ~i21),
  v8138 = (v8139 & i22) | (v7647 & ~i22),
  v8139 = (v7952 & i27) | (v7058 & ~i27),
  v8140 = (v8141 & i21) | (v7647 & ~i21),
  v8141 = (v8142 & i22) | (v7647 & ~i22),
  v8142 = (v7958 & i27) | (v7065 & ~i27),
  v8143 = (v8151 & i19) | (v8144 & ~i19),
  v8144 = (v8148 & i20) | (v8145 & ~i20),
  v8145 = (v8146 & i21) | (v7647 & ~i21),
  v8146 = (v8147 & i22) | (v7647 & ~i22),
  v8147 = (v7966 & i27) | (v7074 & ~i27),
  v8148 = (v8149 & i21) | (v7647 & ~i21),
  v8149 = (v8150 & i22) | (v7647 & ~i22),
  v8150 = (v7972 & i27) | (v7081 & ~i27),
  v8151 = (v8152 & i21) | (v7647 & ~i21),
  v8152 = (v8153 & i22) | (v7647 & ~i22),
  v8153 = (v7978 & i27) | (v7088 & ~i27),
  v8154 = (v8170 & i17) | (v8155 & ~i17),
  v8155 = (v8163 & i19) | (v8156 & ~i19),
  v8156 = (v8160 & i20) | (v8157 & ~i20),
  v8157 = (v8158 & i21) | (v7647 & ~i21),
  v8158 = (v8159 & i22) | (v7647 & ~i22),
  v8159 = (v7987 & i27) | (v7098 & ~i27),
  v8160 = (v8161 & i21) | (v7647 & ~i21),
  v8161 = (v8162 & i22) | (v7647 & ~i22),
  v8162 = (v7993 & i27) | (v7105 & ~i27),
  v8163 = (v8167 & i20) | (v8164 & ~i20),
  v8164 = (v8165 & i21) | (v7647 & ~i21),
  v8165 = (v8166 & i22) | (v7647 & ~i22),
  v8166 = (v8000 & i27) | (v7113 & ~i27),
  v8167 = (v8168 & i21) | (v7647 & ~i21),
  v8168 = (v8169 & i22) | (v7647 & ~i22),
  v8169 = (v8006 & i27) | (v7120 & ~i27),
  v8170 = (v8178 & i19) | (v8171 & ~i19),
  v8171 = (v8175 & i20) | (v8172 & ~i20),
  v8172 = (v8173 & i21) | (v7647 & ~i21),
  v8173 = (v8174 & i22) | (v7647 & ~i22),
  v8174 = (v8014 & i27) | (v7129 & ~i27),
  v8175 = (v8176 & i21) | (v7647 & ~i21),
  v8176 = (v8177 & i22) | (v7647 & ~i22),
  v8177 = (v8020 & i27) | (v7136 & ~i27),
  v8178 = (v8179 & i21) | (v7647 & ~i21),
  v8179 = (v8180 & i22) | (v7647 & ~i22),
  v8180 = (v8026 & i27) | (v7143 & ~i27),
  v8181 = (v8209 & i16) | (v8182 & ~i16),
  v8182 = (v8198 & i17) | (v8183 & ~i17),
  v8183 = (v8191 & i19) | (v8184 & ~i19),
  v8184 = (v8188 & i20) | (v8185 & ~i20),
  v8185 = (v8186 & i21) | (v7647 & ~i21),
  v8186 = (v8187 & i22) | (v7647 & ~i22),
  v8187 = (v8036 & i27) | (v7154 & ~i27),
  v8188 = (v8189 & i21) | (v7647 & ~i21),
  v8189 = (v8190 & i22) | (v7647 & ~i22),
  v8190 = (v8042 & i27) | (v7161 & ~i27),
  v8191 = (v8195 & i20) | (v8192 & ~i20),
  v8192 = (v8193 & i21) | (v7647 & ~i21),
  v8193 = (v8194 & i22) | (v7647 & ~i22),
  v8194 = (v8049 & i27) | (v7169 & ~i27),
  v8195 = (v8196 & i21) | (v7647 & ~i21),
  v8196 = (v8197 & i22) | (v7647 & ~i22),
  v8197 = (v8055 & i27) | (v7176 & ~i27),
  v8198 = (v8206 & i19) | (v8199 & ~i19),
  v8199 = (v8203 & i20) | (v8200 & ~i20),
  v8200 = (v8201 & i21) | (v7647 & ~i21),
  v8201 = (v8202 & i22) | (v7647 & ~i22),
  v8202 = (v8063 & i27) | (v7185 & ~i27),
  v8203 = (v8204 & i21) | (v7647 & ~i21),
  v8204 = (v8205 & i22) | (v7647 & ~i22),
  v8205 = (v8069 & i27) | (v7192 & ~i27),
  v8206 = (v8207 & i21) | (v7647 & ~i21),
  v8207 = (v8208 & i22) | (v7647 & ~i22),
  v8208 = (v8075 & i27) | (v7199 & ~i27),
  v8209 = (v8225 & i17) | (v8210 & ~i17),
  v8210 = (v8218 & i19) | (v8211 & ~i19),
  v8211 = (v8215 & i20) | (v8212 & ~i20),
  v8212 = (v8213 & i21) | (v7647 & ~i21),
  v8213 = (v8214 & i22) | (v7647 & ~i22),
  v8214 = (v8084 & i27) | (v7209 & ~i27),
  v8215 = (v8216 & i21) | (v7647 & ~i21),
  v8216 = (v8217 & i22) | (v7647 & ~i22),
  v8217 = (v8090 & i27) | (v7216 & ~i27),
  v8218 = (v8222 & i20) | (v8219 & ~i20),
  v8219 = (v8220 & i21) | (v7647 & ~i21),
  v8220 = (v8221 & i22) | (v7647 & ~i22),
  v8221 = (v8097 & i27) | (v7224 & ~i27),
  v8222 = (v8223 & i21) | (v7647 & ~i21),
  v8223 = (v8224 & i22) | (v7647 & ~i22),
  v8224 = (v8103 & i27) | (v7231 & ~i27),
  v8225 = (v8233 & i19) | (v8226 & ~i19),
  v8226 = (v8230 & i20) | (v8227 & ~i20),
  v8227 = (v8228 & i21) | (v7647 & ~i21),
  v8228 = (v8229 & i22) | (v7647 & ~i22),
  v8229 = (v8111 & i27) | (v7240 & ~i27),
  v8230 = (v8231 & i21) | (v7647 & ~i21),
  v8231 = (v8232 & i22) | (v7647 & ~i22),
  v8232 = (v8117 & i27) | (v7247 & ~i27),
  v8233 = (v8234 & i21) | (v7647 & ~i21),
  v8234 = (v8235 & i22) | (v7647 & ~i22),
  v8235 = (v8123 & i27) | (v7254 & ~i27),
  v8236 = (v7036 & i12) | (v8237 & ~i12),
  v8237 = (v7036 & i13) | (v8238 & ~i13),
  v8238 = (v8239 & i14) | (v7036 & ~i14),
  v8239 = (v8295 & i15) | (v8240 & ~i15),
  v8240 = (v8268 & i16) | (v8241 & ~i16),
  v8241 = (v8257 & i17) | (v8242 & ~i17),
  v8242 = (v8250 & i19) | (v8243 & ~i19),
  v8243 = (v8247 & i20) | (v8244 & ~i20),
  v8244 = (v8245 & i21) | (v7791 & ~i21),
  v8245 = (v8246 & i22) | (v7791 & ~i22),
  v8246 = (v7938 & i26) | (v7043 & ~i26),
  v8247 = (v8248 & i21) | (v7791 & ~i21),
  v8248 = (v8249 & i22) | (v7791 & ~i22),
  v8249 = (v7944 & i26) | (v7050 & ~i26),
  v8250 = (v8254 & i20) | (v8251 & ~i20),
  v8251 = (v8252 & i21) | (v7791 & ~i21),
  v8252 = (v8253 & i22) | (v7791 & ~i22),
  v8253 = (v7951 & i26) | (v7058 & ~i26),
  v8254 = (v8255 & i21) | (v7791 & ~i21),
  v8255 = (v8256 & i22) | (v7791 & ~i22),
  v8256 = (v7957 & i26) | (v7065 & ~i26),
  v8257 = (v8265 & i19) | (v8258 & ~i19),
  v8258 = (v8262 & i20) | (v8259 & ~i20),
  v8259 = (v8260 & i21) | (v7791 & ~i21),
  v8260 = (v8261 & i22) | (v7791 & ~i22),
  v8261 = (v7965 & i26) | (v7074 & ~i26),
  v8262 = (v8263 & i21) | (v7791 & ~i21),
  v8263 = (v8264 & i22) | (v7791 & ~i22),
  v8264 = (v7971 & i26) | (v7081 & ~i26),
  v8265 = (v8266 & i21) | (v7791 & ~i21),
  v8266 = (v8267 & i22) | (v7791 & ~i22),
  v8267 = (v7977 & i26) | (v7088 & ~i26),
  v8268 = (v8284 & i17) | (v8269 & ~i17),
  v8269 = (v8277 & i19) | (v8270 & ~i19),
  v8270 = (v8274 & i20) | (v8271 & ~i20),
  v8271 = (v8272 & i21) | (v7791 & ~i21),
  v8272 = (v8273 & i22) | (v7791 & ~i22),
  v8273 = (v7986 & i26) | (v7098 & ~i26),
  v8274 = (v8275 & i21) | (v7791 & ~i21),
  v8275 = (v8276 & i22) | (v7791 & ~i22),
  v8276 = (v7992 & i26) | (v7105 & ~i26),
  v8277 = (v8281 & i20) | (v8278 & ~i20),
  v8278 = (v8279 & i21) | (v7791 & ~i21),
  v8279 = (v8280 & i22) | (v7791 & ~i22),
  v8280 = (v7999 & i26) | (v7113 & ~i26),
  v8281 = (v8282 & i21) | (v7791 & ~i21),
  v8282 = (v8283 & i22) | (v7791 & ~i22),
  v8283 = (v8005 & i26) | (v7120 & ~i26),
  v8284 = (v8292 & i19) | (v8285 & ~i19),
  v8285 = (v8289 & i20) | (v8286 & ~i20),
  v8286 = (v8287 & i21) | (v7791 & ~i21),
  v8287 = (v8288 & i22) | (v7791 & ~i22),
  v8288 = (v8013 & i26) | (v7129 & ~i26),
  v8289 = (v8290 & i21) | (v7791 & ~i21),
  v8290 = (v8291 & i22) | (v7791 & ~i22),
  v8291 = (v8019 & i26) | (v7136 & ~i26),
  v8292 = (v8293 & i21) | (v7791 & ~i21),
  v8293 = (v8294 & i22) | (v7791 & ~i22),
  v8294 = (v8025 & i26) | (v7143 & ~i26),
  v8295 = (v8323 & i16) | (v8296 & ~i16),
  v8296 = (v8312 & i17) | (v8297 & ~i17),
  v8297 = (v8305 & i19) | (v8298 & ~i19),
  v8298 = (v8302 & i20) | (v8299 & ~i20),
  v8299 = (v8300 & i21) | (v7791 & ~i21),
  v8300 = (v8301 & i22) | (v7791 & ~i22),
  v8301 = (v8035 & i26) | (v7154 & ~i26),
  v8302 = (v8303 & i21) | (v7791 & ~i21),
  v8303 = (v8304 & i22) | (v7791 & ~i22),
  v8304 = (v8041 & i26) | (v7161 & ~i26),
  v8305 = (v8309 & i20) | (v8306 & ~i20),
  v8306 = (v8307 & i21) | (v7791 & ~i21),
  v8307 = (v8308 & i22) | (v7791 & ~i22),
  v8308 = (v8048 & i26) | (v7169 & ~i26),
  v8309 = (v8310 & i21) | (v7791 & ~i21),
  v8310 = (v8311 & i22) | (v7791 & ~i22),
  v8311 = (v8054 & i26) | (v7176 & ~i26),
  v8312 = (v8320 & i19) | (v8313 & ~i19),
  v8313 = (v8317 & i20) | (v8314 & ~i20),
  v8314 = (v8315 & i21) | (v7791 & ~i21),
  v8315 = (v8316 & i22) | (v7791 & ~i22),
  v8316 = (v8062 & i26) | (v7185 & ~i26),
  v8317 = (v8318 & i21) | (v7791 & ~i21),
  v8318 = (v8319 & i22) | (v7791 & ~i22),
  v8319 = (v8068 & i26) | (v7192 & ~i26),
  v8320 = (v8321 & i21) | (v7791 & ~i21),
  v8321 = (v8322 & i22) | (v7791 & ~i22),
  v8322 = (v8074 & i26) | (v7199 & ~i26),
  v8323 = (v8339 & i17) | (v8324 & ~i17),
  v8324 = (v8332 & i19) | (v8325 & ~i19),
  v8325 = (v8329 & i20) | (v8326 & ~i20),
  v8326 = (v8327 & i21) | (v7791 & ~i21),
  v8327 = (v8328 & i22) | (v7791 & ~i22),
  v8328 = (v8083 & i26) | (v7209 & ~i26),
  v8329 = (v8330 & i21) | (v7791 & ~i21),
  v8330 = (v8331 & i22) | (v7791 & ~i22),
  v8331 = (v8089 & i26) | (v7216 & ~i26),
  v8332 = (v8336 & i20) | (v8333 & ~i20),
  v8333 = (v8334 & i21) | (v7791 & ~i21),
  v8334 = (v8335 & i22) | (v7791 & ~i22),
  v8335 = (v8096 & i26) | (v7224 & ~i26),
  v8336 = (v8337 & i21) | (v7791 & ~i21),
  v8337 = (v8338 & i22) | (v7791 & ~i22),
  v8338 = (v8102 & i26) | (v7231 & ~i26),
  v8339 = (v8347 & i19) | (v8340 & ~i19),
  v8340 = (v8344 & i20) | (v8341 & ~i20),
  v8341 = (v8342 & i21) | (v7791 & ~i21),
  v8342 = (v8343 & i22) | (v7791 & ~i22),
  v8343 = (v8110 & i26) | (v7240 & ~i26),
  v8344 = (v8345 & i21) | (v7791 & ~i21),
  v8345 = (v8346 & i22) | (v7791 & ~i22),
  v8346 = (v8116 & i26) | (v7247 & ~i26),
  v8347 = (v8348 & i21) | (v7791 & ~i21),
  v8348 = (v8349 & i22) | (v7791 & ~i22),
  v8349 = (v8122 & i26) | (v7254 & ~i26),
  v8350 = (v8358 & i11) | (v8351 & ~i11),
  v8351 = (v8352 & i12) | (v7344 & ~i12),
  v8352 = (v7346 & i13) | (v8353 & ~i13),
  v8353 = (v8356 & i14) | (v8354 & ~i14),
  v8354 = (v8355 & i21) | (v7445 & ~i21),
  v8355 = (v7451 & i22) | (v7445 & ~i22),
  v8356 = (v8357 & i21) | (v7647 & ~i21),
  v8357 = (v7650 & i22) | (v7647 & ~i22),
  v8358 = (v7346 & i12) | (v8359 & ~i12),
  v8359 = (v7346 & i13) | (v8360 & ~i13),
  v8360 = (v8361 & i14) | (v7346 & ~i14),
  v8361 = (v8362 & i21) | (v7791 & ~i21),
  v8362 = (v7794 & i22) | (v7791 & ~i22),
  v8363 = (v8350 & i9) | (v8364 & ~i9),
  v8364 = (v8634 & i10) | (v8365 & ~i10),
  v8365 = (v8623 & i11) | (v8366 & ~i11),
  v8366 = (v8601 & i12) | (v8367 & ~i12),
  v8367 = (v8369 & i13) | (v8368 & ~i13),
  v8368 = (v8378 & i14) | (v8369 & ~i14),
  v8369 = (v8374 & i21) | (v8370 & ~i21),
  v8370 = (v6456 & i23) | (v8371 & ~i23),
  v8371 = (v6456 & i24) | (v8372 & ~i24),
  v8372 = v8373 & i30,
  v8373 = (v63 & ~i31) | i31,
  v8374 = (v8375 & i22) | (v8370 & ~i22),
  v8375 = (v6459 & i23) | (v8376 & ~i23),
  v8376 = (v6459 & i24) | (v8377 & ~i24),
  v8377 = (v8373 & i30) | (~v6460 & ~i30),
  v8378 = (v8490 & i15) | (v8379 & ~i15),
  v8379 = (v8435 & i16) | (v8380 & ~i16),
  v8380 = (v8412 & i17) | (v8381 & ~i17),
  v8381 = (v8397 & i19) | (v8382 & ~i19),
  v8382 = (v8390 & i20) | (v8383 & ~i20),
  v8383 = (v8384 & i21) | (v8370 & ~i21),
  v8384 = (v8385 & i22) | (v8370 & ~i22),
  v8385 = (v6789 & i23) | (v8386 & ~i23),
  v8386 = (v6789 & i24) | (v8387 & ~i24),
  v8387 = (v8389 & i29) | (v8388 & ~i29),
  v8388 = (v8373 & i30) | (~v6466 & ~i30),
  v8389 = (v8373 & i30) | (~v6791 & ~i30),
  v8390 = (v8391 & i21) | (v8370 & ~i21),
  v8391 = (v8392 & i22) | (v8370 & ~i22),
  v8392 = (v6797 & i23) | (v8393 & ~i23),
  v8393 = (v6797 & i24) | (v8394 & ~i24),
  v8394 = (v8396 & i29) | (v8395 & ~i29),
  v8395 = (v8373 & i30) | (~v6480 & ~i30),
  v8396 = (v8373 & i30) | (~v6799 & ~i30),
  v8397 = (v8405 & i20) | (v8398 & ~i20),
  v8398 = (v8399 & i21) | (v8370 & ~i21),
  v8399 = (v8400 & i22) | (v8370 & ~i22),
  v100 = (v102 & i31) | (~v101 & ~i31),
  v101 = (v99 & ~i32) | i32,
  v102 = (~v99 & ~i32) | i32,
  v103 = (v105 & i30) | (~v104 & ~i30),
  v104 = (v87 & i40) | (v78 & ~i40),
  v105 = (v107 & i31) | (~v106 & ~i31),
  v106 = (v104 & ~i32) | i32,
  v107 = (~v104 & ~i32) | i32,
  v108 = (v109 & i30) | (~v87 & ~i30),
  v109 = (v111 & i31) | (~v110 & ~i31),
  v110 = (v87 & ~i32) | i32,
  v111 = (~v87 & ~i32) | i32,
  v112 = (v136 & i17) | (v113 & ~i17),
  v113 = (v125 & i19) | (v114 & ~i19),
  v114 = (v120 & i20) | (v115 & ~i20),
  v115 = (v117 & i30) | (~v116 & ~i30),
  v116 = (v72 & i41) | (v70 & ~i41),
  v117 = (v119 & i31) | (~v118 & ~i31),
  v118 = (v116 & ~i32) | i32,
  v119 = (~v116 & ~i32) | i32,
  v120 = (v122 & i30) | (~v121 & ~i30),
  v121 = (v72 & i41) | (v79 & ~i41),
  v122 = (v124 & i31) | (~v123 & ~i31),
  v123 = (v121 & ~i32) | i32,
  v124 = (~v121 & ~i32) | i32,
  v125 = (v131 & i20) | (v126 & ~i20),
  v126 = (v128 & i30) | (~v127 & ~i30),
  v127 = (v116 & i40) | (v72 & ~i40),
  v128 = (v130 & i31) | (~v129 & ~i31),
  v129 = (v127 & ~i32) | i32,
  v130 = (~v127 & ~i32) | i32,
  v131 = (v133 & i30) | (~v132 & ~i30),
  v132 = (v121 & i40) | (v72 & ~i40),
  v133 = (v135 & i31) | (~v134 & ~i31),
  v134 = (v132 & ~i32) | i32,
  v135 = (~v132 & ~i32) | i32,
  v136 = (v148 & i19) | (v137 & ~i19),
  v137 = (v143 & i20) | (v138 & ~i20),
  v138 = (v140 & i30) | (~v139 & ~i30),
  v139 = (v72 & i40) | (v116 & ~i40),
  v8400 = (v6806 & i23) | (v8401 & ~i23),
  v8401 = (v6806 & i24) | (v8402 & ~i24),
  v8402 = (v8404 & i29) | (v8403 & ~i29),
  v8403 = (v8373 & i30) | (~v6495 & ~i30),
  v8404 = (v8373 & i30) | (~v6808 & ~i30),
  v8405 = (v8406 & i21) | (v8370 & ~i21),
  v8406 = (v8407 & i22) | (v8370 & ~i22),
  v140 = (v142 & i31) | (~v141 & ~i31),
  v8407 = (v6814 & i23) | (v8408 & ~i23),
  v141 = (v139 & ~i32) | i32,
  v8408 = (v6814 & i24) | (v8409 & ~i24),
  v142 = (~v139 & ~i32) | i32,
  v8409 = (v8411 & i29) | (v8410 & ~i29),
  v143 = (v145 & i30) | (~v144 & ~i30),
  v144 = (v72 & i40) | (v121 & ~i40),
  v145 = (v147 & i31) | (~v146 & ~i31),
  v146 = (v144 & ~i32) | i32,
  v147 = (~v144 & ~i32) | i32,
  v148 = (v149 & i30) | (~v72 & ~i30),
  v149 = (v151 & i31) | (~v150 & ~i31),
  v8410 = (v8373 & i30) | (~v6511 & ~i30),
  v8411 = (v8373 & i30) | (~v6816 & ~i30),
  v8412 = (v8428 & i19) | (v8413 & ~i19),
  v8413 = (v8421 & i20) | (v8414 & ~i20),
  v8414 = (v8415 & i21) | (v8370 & ~i21),
  v8415 = (v8416 & i22) | (v8370 & ~i22),
  v8416 = (v6824 & i23) | (v8417 & ~i23),
  v150 = (v72 & ~i32) | i32,
  v8417 = (v6824 & i24) | (v8418 & ~i24),
  v151 = (~v72 & ~i32) | i32,
  v8418 = (v8420 & i29) | (v8419 & ~i29),
  v152 = (v207 & i16) | (v153 & ~i16),
  v8419 = (v8373 & i30) | (~v6528 & ~i30),
  v153 = (v155 & i17) | (v154 & ~i17),
  v154 = (v174 & i18) | (v155 & ~i18),
  v155 = (v168 & i30) | (~v156 & ~i30),
  v156 = (v161 & i37) | (v157 & ~i37),
  v157 = (v161 & i38) | (~v158 & ~i38),
  v158 = (v160 & i41) | (v159 & ~i41),
  v159 = (v72 & i42) | ~i42,
  v8420 = (v8373 & i30) | (~v6826 & ~i30),
  v8421 = (v8422 & i21) | (v8370 & ~i21),
  v8422 = (v8423 & i22) | (v8370 & ~i22),
  v8423 = (v6832 & i23) | (v8424 & ~i23),
  v8424 = (v6832 & i24) | (v8425 & ~i24),
  v8425 = (v8427 & i29) | (v8426 & ~i29),
  v8426 = (v8373 & i30) | (~v6543 & ~i30),
  v160 = (~v72 & ~i42) | (v72 & i42),
  v8427 = (v8373 & i30) | (~v6834 & ~i30),
  v161 = (v165 & i39) | (~v162 & ~i39),
  v8428 = (v8429 & i21) | (v8370 & ~i21),
  v162 = (v164 & i41) | (v163 & ~i41),
  v8429 = (v8430 & i22) | (v8370 & ~i22),
  v163 = (v71 & i42) | ~i42,
  v164 = (v71 & i42) | (~v72 & ~i42),
  v165 = (v167 & i41) | (v166 & ~i41),
  v166 = v80 & i42,
  v167 = (v80 & i42) | (v72 & ~i42),
  v168 = (v173 & i31) | (~v169 & ~i31),
  v169 = (v170 & i32) | (v161 & ~i32),
  v8430 = (v6840 & i23) | (v8431 & ~i23),
  v8431 = (v6840 & i24) | (v8432 & ~i24),
  v8432 = (v8434 & i29) | (v8433 & ~i29),
  v8433 = (v8373 & i30) | (~v6558 & ~i30),
  v8434 = (v8373 & i30) | (~v6842 & ~i30),
  v8435 = (v8467 & i17) | (v8436 & ~i17),
  v8436 = (v8452 & i19) | (v8437 & ~i19),
  v170 = (v172 & i37) | (v171 & ~i37),
  v8437 = (v8445 & i20) | (v8438 & ~i20),
  v171 = v172 & i38,
  v8438 = (v8439 & i21) | (v8370 & ~i21),
  v172 = (~v60 & ~i39) | (v60 & i39),
  v8439 = (v8440 & i22) | (v8370 & ~i22),
  v173 = (~v161 & ~i32) | i32,
  v174 = (v191 & i20) | (v175 & ~i20),
  v175 = (v188 & i30) | (~v176 & ~i30),
  v176 = (v181 & i37) | (v177 & ~i37),
  v177 = (v181 & i38) | (~v178 & ~i38),
  v178 = (v179 & i40) | (v158 & ~i40),
  v179 = (v160 & i41) | (v180 & ~i41),
  v8440 = (v6851 & i23) | (v8441 & ~i23),
  v8441 = (v6851 & i24) | (v8442 & ~i24),
  v8442 = (v8444 & i29) | (v8443 & ~i29),
  v8443 = (v8373 & i30) | (~v6570 & ~i30),
  v8444 = (v8373 & i30) | (~v6853 & ~i30),
  v8445 = (v8446 & i21) | (v8370 & ~i21),
  v8446 = (v8447 & i22) | (v8370 & ~i22),
  v180 = (v72 & i42) | (v80 & ~i42),
  v8447 = (v6859 & i23) | (v8448 & ~i23),
  v181 = (v185 & i39) | (~v182 & ~i39),
  v8448 = (v6859 & i24) | (v8449 & ~i24),
  v182 = (v183 & i40) | (v162 & ~i40),
  v8449 = (v8451 & i29) | (v8450 & ~i29),
  v183 = (v164 & i41) | (v184 & ~i41),
  v184 = (v71 & i42) | (v80 & ~i42),
  v185 = (v186 & i40) | (v165 & ~i40),
  v186 = (v167 & i41) | (v187 & ~i41),
  v187 = (~v80 & ~i42) | (v80 & i42),
  v188 = (v190 & i31) | (~v189 & ~i31),
  v189 = (v170 & i32) | (v181 & ~i32),
  v8450 = (v8373 & i30) | (~v6583 & ~i30),
  v8451 = (v8373 & i30) | (~v6861 & ~i30),
  v8452 = (v8460 & i20) | (v8453 & ~i20),
  v8453 = (v8454 & i21) | (v8370 & ~i21),
  v8454 = (v8455 & i22) | (v8370 & ~i22),
  v8455 = (v6868 & i23) | (v8456 & ~i23),
  v8456 = (v6868 & i24) | (v8457 & ~i24),
  v190 = (~v181 & ~i32) | i32,
  v8457 = (v8459 & i29) | (v8458 & ~i29),
  v191 = (v204 & i30) | (~v192 & ~i30),
  v8458 = (v8373 & i30) | (~v6597 & ~i30),
  v192 = (v197 & i37) | (v193 & ~i37),
  v8459 = (v8373 & i30) | (~v6870 & ~i30),
  v193 = (v197 & i38) | (~v194 & ~i38),
  v194 = (v195 & i40) | (v158 & ~i40),
  v195 = (v160 & i41) | (v196 & ~i41),
  v196 = (v72 & i42) | (~v71 & ~i42),
  v197 = (v201 & i39) | (~v198 & ~i39),
  v198 = (v199 & i40) | (v162 & ~i40),
  v199 = (v164 & i41) | (v200 & ~i41),
  v8460 = (v8461 & i21) | (v8370 & ~i21),
  v8461 = (v8462 & i22) | (v8370 & ~i22),
  v8462 = (v6876 & i23) | (v8463 & ~i23),
  v8463 = (v6876 & i24) | (v8464 & ~i24),
  v8464 = (v8466 & i29) | (v8465 & ~i29),
  v8465 = (v8373 & i30) | (~v6612 & ~i30),
  v8466 = (v8373 & i30) | (~v6878 & ~i30),
  v8467 = (v8483 & i19) | (v8468 & ~i19),
  v8468 = (v8476 & i20) | (v8469 & ~i20),
  v8469 = (v8470 & i21) | (v8370 & ~i21),
  v8470 = (v8471 & i22) | (v8370 & ~i22),
  v8471 = (v6886 & i23) | (v8472 & ~i23),
  v8472 = (v6886 & i24) | (v8473 & ~i24),
  v8473 = (v8475 & i29) | (v8474 & ~i29),
  v8474 = (v8373 & i30) | (~v6629 & ~i30),
  v8475 = (v8373 & i30) | (~v6888 & ~i30),
  v8476 = (v8477 & i21) | (v8370 & ~i21),
  v8477 = (v8478 & i22) | (v8370 & ~i22),
  v8478 = (v6894 & i23) | (v8479 & ~i23),
  v8479 = (v6894 & i24) | (v8480 & ~i24),
  v8480 = (v8482 & i29) | (v8481 & ~i29),
  v8481 = (v8373 & i30) | (~v6644 & ~i30),
  v8482 = (v8373 & i30) | (~v6896 & ~i30),
  v8483 = (v8484 & i21) | (v8370 & ~i21),
  v8484 = (v8485 & i22) | (v8370 & ~i22),
  v8485 = (v6902 & i23) | (v8486 & ~i23),
  v8486 = (v6902 & i24) | (v8487 & ~i24),
  v8487 = (v8489 & i29) | (v8488 & ~i29),
  v8488 = (v8373 & i30) | (~v6659 & ~i30),
  v8489 = (v8373 & i30) | (~v6904 & ~i30),
  v8490 = (v8546 & i16) | (v8491 & ~i16),
  v8491 = (v8523 & i17) | (v8492 & ~i17),
  v8492 = (v8508 & i19) | (v8493 & ~i19),
  v8493 = (v8501 & i20) | (v8494 & ~i20),
  v8494 = (v8495 & i21) | (v8370 & ~i21),
  v8495 = (v8496 & i22) | (v8370 & ~i22),
  v8496 = (v6914 & i23) | (v8497 & ~i23),
  v8497 = (v6914 & i24) | (v8498 & ~i24),
  v8498 = (v8500 & i29) | (v8499 & ~i29),
  v8499 = (v8373 & i30) | (~v6672 & ~i30),
  v200 = (~v71 & ~i42) | (v71 & i42),
  v201 = (v202 & i40) | (v165 & ~i40),
  v202 = (v167 & i41) | (v203 & ~i41),
  v203 = (v80 & i42) | (v71 & ~i42),
  v204 = (v206 & i31) | (~v205 & ~i31),
  v205 = (v170 & i32) | (v197 & ~i32),
  v206 = (~v197 & ~i32) | i32,
  v207 = (v209 & i17) | (v208 & ~i17),
  v208 = (v216 & i18) | (v209 & ~i18),
  v209 = (v213 & i30) | (~v210 & ~i30),
  v210 = (v212 & i37) | (v211 & ~i37),
  v211 = (v212 & i38) | (~v159 & ~i38),
  v212 = (v166 & i39) | (~v163 & ~i39),
  v213 = (v215 & i31) | (~v214 & ~i31),
  v214 = (v170 & i32) | (v212 & ~i32),
  v215 = (~v212 & ~i32) | i32,
  v216 = (v230 & i20) | (v217 & ~i20),
  v217 = (v227 & i30) | (~v218 & ~i30),
  v218 = (v222 & i37) | (v219 & ~i37),
  v219 = (v222 & i38) | (~v220 & ~i38),
  v220 = (v221 & i40) | (v159 & ~i40),
  v221 = (v159 & i41) | (v180 & ~i41),
  v222 = (v225 & i39) | (~v223 & ~i39),
  v223 = (v224 & i40) | (v163 & ~i40),
  v224 = (v163 & i41) | (v184 & ~i41),
  v225 = (v226 & i40) | (v166 & ~i40),
  v226 = (v166 & i41) | (v187 & ~i41),
  v227 = (v229 & i31) | (~v228 & ~i31),
  v228 = (v170 & i32) | (v222 & ~i32),
  v229 = (~v222 & ~i32) | i32,
  v230 = (v240 & i30) | (~v231 & ~i30),
  v231 = (v235 & i37) | (v232 & ~i37),
  v232 = (v235 & i38) | (~v233 & ~i38),
  v233 = (v234 & i40) | (v159 & ~i40),
  v234 = (v159 & i41) | (v196 & ~i41),
  v235 = (v238 & i39) | (~v236 & ~i39),
  v236 = (v237 & i40) | (v163 & ~i40),
  v237 = (v163 & i41) | (v200 & ~i41),
  v238 = (v239 & i40) | (v166 & ~i40),
  v239 = (v166 & i41) | (v203 & ~i41),
  v8500 = (v8373 & i30) | (~v6916 & ~i30),
  v8501 = (v8502 & i21) | (v8370 & ~i21),
  v8502 = (v8503 & i22) | (v8370 & ~i22),
  v8503 = (v6922 & i23) | (v8504 & ~i23),
  v8504 = (v6922 & i24) | (v8505 & ~i24),
  v8505 = (v8507 & i29) | (v8506 & ~i29),
  v8506 = (v8373 & i30) | (~v6679 & ~i30),
  v240 = (v242 & i31) | (~v241 & ~i31),
  v8507 = (v8373 & i30) | (~v6924 & ~i30),
  v241 = (v170 & i32) | (v235 & ~i32),
  v8508 = (v8516 & i20) | (v8509 & ~i20),
  v242 = (~v235 & ~i32) | i32,
  v8509 = (v8510 & i21) | (v8370 & ~i21),
  v243 = (v254 & i2) | (v244 & ~i2),
  v244 = (v254 & i3) | (v245 & ~i3),
  v245 = (v254 & i4) | (v246 & ~i4),
  v246 = (v254 & i5) | (v247 & ~i5),
  v247 = (v254 & i6) | (v248 & ~i6),
  v248 = (v251 & i7) | (v249 & ~i7),
  v249 = (v251 & i8) | (v250 & ~i8),
  v8510 = (v8511 & i22) | (v8370 & ~i22),
  v8511 = (v6931 & i23) | (v8512 & ~i23),
  v8512 = (v6931 & i24) | (v8513 & ~i24),
  v8513 = (v8515 & i29) | (v8514 & ~i29),
  v8514 = (v8373 & i30) | (~v6687 & ~i30),
  v8515 = (v8373 & i30) | (~v6933 & ~i30),
  v8516 = (v8517 & i21) | (v8370 & ~i21),
  v250 = (v265 & i9) | (v251 & ~i9),
  v8517 = (v8518 & i22) | (v8370 & ~i22),
  v251 = (v254 & i11) | (v252 & ~i11),
  v8518 = (v6939 & i23) | (v8519 & ~i23),
  v252 = (v254 & i12) | (v253 & ~i12),
  v8519 = (v6939 & i24) | (v8520 & ~i24),
  v253 = (v255 & i13) | (v254 & ~i13),
  v254 = i41,
  v255 = (v256 & i14) | (v254 & ~i14),
  v256 = (v261 & i27) | (v257 & ~i27),
  v257 = (v258 & i30) | (v254 & ~i30),
  v258 = (v254 & i31) | (~v259 & ~i31),
  v259 = (v260 & i32) | (~v254 & ~i32),
  v8520 = (v8522 & i29) | (v8521 & ~i29),
  v8521 = (v8373 & i30) | (~v6695 & ~i30),
  v8522 = (v8373 & i30) | (~v6941 & ~i30),
  v8523 = (v8539 & i19) | (v8524 & ~i19),
  v8524 = (v8532 & i20) | (v8525 & ~i20),
  v8525 = (v8526 & i21) | (v8370 & ~i21),
  v8526 = (v8527 & i22) | (v8370 & ~i22),
  v260 = (~v254 & ~i33) | i33,
  v8527 = (v6949 & i23) | (v8528 & ~i23),
  v261 = (v262 & i30) | (v254 & ~i30),
  v8528 = (v6949 & i24) | (v8529 & ~i24),
  v262 = (v254 & i31) | (v263 & ~i31),
  v8529 = (v8531 & i29) | (v8530 & ~i29),
  v263 = (v264 & i32) | (v254 & ~i32),
  v264 = (v254 & ~i33) | i33,
  v265 = (v266 & i10) | (v251 & ~i10),
  v266 = (v269 & i11) | (v267 & ~i11),
  v267 = (v269 & i12) | (v268 & ~i12),
  v268 = (v278 & i13) | (v269 & ~i13),
  v269 = (v274 & i24) | (v270 & ~i24),
  v8530 = (v8373 & i30) | (~v6705 & ~i30),
  v8531 = (v8373 & i30) | (~v6951 & ~i30),
  v8532 = (v8533 & i21) | (v8370 & ~i21),
  v8533 = (v8534 & i22) | (v8370 & ~i22),
  v8534 = (v6957 & i23) | (v8535 & ~i23),
  v8535 = (v6957 & i24) | (v8536 & ~i24),
  v8536 = (v8538 & i29) | (v8537 & ~i29),
  v270 = (v271 & i30) | (v254 & ~i30),
  v8537 = (v8373 & i30) | (~v6713 & ~i30),
  v271 = (v254 & i31) | (v272 & ~i31),
  v8538 = (v8373 & i30) | (~v6959 & ~i30),
  v272 = (v273 & i32) | (v254 & ~i32),
  v8539 = (v8540 & i21) | (v8370 & ~i21),
  v273 = v254 & i33,
  v274 = (v275 & i30) | (v254 & ~i30),
  v275 = (v254 & i31) | (v276 & ~i31),
  v276 = (v277 & i32) | (v254 & ~i32),
  v277 = (v254 & i33) | ~i33,
  v278 = (v279 & i14) | (v269 & ~i14),
  v279 = (v287 & i24) | (v280 & ~i24),
  v8540 = (v8541 & i22) | (v8370 & ~i22),
  v8541 = (v6965 & i23) | (v8542 & ~i23),
  v8542 = (v6965 & i24) | (v8543 & ~i24),
  v8543 = (v8545 & i29) | (v8544 & ~i29),
  v8544 = (v8373 & i30) | (~v6721 & ~i30),
  v8545 = (v8373 & i30) | (~v6967 & ~i30),
  v8546 = (v8578 & i17) | (v8547 & ~i17),
  v280 = (v284 & i27) | (v281 & ~i27),
  v8547 = (v8563 & i19) | (v8548 & ~i19),
  v281 = (v282 & i30) | (v254 & ~i30),
  v8548 = (v8556 & i20) | (v8549 & ~i20),
  v282 = (v254 & i31) | (~v283 & ~i31),
  v8549 = (v8550 & i21) | (v8370 & ~i21),
  v283 = (~v254 & ~i32) | i32,
  v284 = (v285 & i30) | (v254 & ~i30),
  v285 = (v254 & i31) | (v286 & ~i31),
  v286 = (v63 & i32) | (v254 & ~i32),
  v287 = (v291 & i27) | (v288 & ~i27),
  v288 = (v289 & i30) | (v254 & ~i30),
  v289 = (v254 & i31) | (~v290 & ~i31),
  v8550 = (v8551 & i22) | (v8370 & ~i22),
  v8551 = (v6976 & i23) | (v8552 & ~i23),
  v8552 = (v6976 & i24) | (v8553 & ~i24),
  v8553 = (v8555 & i29) | (v8554 & ~i29),
  v8554 = (v8373 & i30) | (~v6730 & ~i30),
  v8555 = (v8373 & i30) | (~v6978 & ~i30),
  v8556 = (v8557 & i21) | (v8370 & ~i21),
  v290 = (v63 & i32) | (~v254 & ~i32),
  v8557 = (v8558 & i22) | (v8370 & ~i22),
  v291 = (v292 & i30) | (v254 & ~i30),
  v8558 = (v6984 & i23) | (v8559 & ~i23),
  v292 = (v254 & i31) | (v293 & ~i31),
  v8559 = (v6984 & i24) | (v8560 & ~i24),
  v293 = (v254 & ~i32) | i32,
  v294 = (v305 & i2) | (v295 & ~i2),
  v295 = (v305 & i3) | (v296 & ~i3),
  v296 = (v305 & i4) | (v297 & ~i4),
  v297 = (v305 & i5) | (v298 & ~i5),
  v298 = (v305 & i6) | (v299 & ~i6),
  v299 = (v302 & i7) | (v300 & ~i7),
  v8560 = (v8562 & i29) | (v8561 & ~i29),
  v8561 = (v8373 & i30) | (~v6737 & ~i30),
  v8562 = (v8373 & i30) | (~v6986 & ~i30),
  v8563 = (v8571 & i20) | (v8564 & ~i20),
  v8564 = (v8565 & i21) | (v8370 & ~i21),
  v8565 = (v8566 & i22) | (v8370 & ~i22),
  v8566 = (v6993 & i23) | (v8567 & ~i23),
  v8567 = (v6993 & i24) | (v8568 & ~i24),
  v8568 = (v8570 & i29) | (v8569 & ~i29),
  v8569 = (v8373 & i30) | (~v6745 & ~i30),
  v8570 = (v8373 & i30) | (~v6995 & ~i30),
  v8571 = (v8572 & i21) | (v8370 & ~i21),
  v8572 = (v8573 & i22) | (v8370 & ~i22),
  v8573 = (v7001 & i23) | (v8574 & ~i23),
  v8574 = (v7001 & i24) | (v8575 & ~i24),
  v8575 = (v8577 & i29) | (v8576 & ~i29),
  v8576 = (v8373 & i30) | (~v6753 & ~i30),
  v8577 = (v8373 & i30) | (~v7003 & ~i30),
  v8578 = (v8594 & i19) | (v8579 & ~i19),
  v8579 = (v8587 & i20) | (v8580 & ~i20),
  v8580 = (v8581 & i21) | (v8370 & ~i21),
  v8581 = (v8582 & i22) | (v8370 & ~i22),
  v8582 = (v7011 & i23) | (v8583 & ~i23),
  v8583 = (v7011 & i24) | (v8584 & ~i24),
  v8584 = (v8586 & i29) | (v8585 & ~i29),
  v8585 = (v8373 & i30) | (~v6763 & ~i30),
  v8586 = (v8373 & i30) | (~v7013 & ~i30),
  v8587 = (v8588 & i21) | (v8370 & ~i21),
  v8588 = (v8589 & i22) | (v8370 & ~i22),
  v8589 = (v7019 & i23) | (v8590 & ~i23),
  v8590 = (v7019 & i24) | (v8591 & ~i24),
  v8591 = (v8593 & i29) | (v8592 & ~i29),
  v8592 = (v8373 & i30) | (~v6771 & ~i30),
  v8593 = (v8373 & i30) | (~v7021 & ~i30),
  v8594 = (v8595 & i21) | (v8370 & ~i21),
  v8595 = (v8596 & i22) | (v8370 & ~i22),
  v8596 = (v7027 & i23) | (v8597 & ~i23),
  v8597 = (v7027 & i24) | (v8598 & ~i24),
  v8598 = (v8600 & i29) | (v8599 & ~i29),
  v8599 = (v8373 & i30) | (~v6779 & ~i30),
  v300 = (v302 & i8) | (v301 & ~i8),
  v301 = (v316 & i9) | (v302 & ~i9),
  v302 = (v305 & i11) | (v303 & ~i11),
  v303 = (v305 & i12) | (v304 & ~i12),
  v304 = (v306 & i13) | (v305 & ~i13),
  v305 = i40,
  v306 = (v307 & i14) | (v305 & ~i14),
  v307 = (v312 & i26) | (v308 & ~i26),
  v308 = (v309 & i30) | (v305 & ~i30),
  v309 = (v305 & i31) | (~v310 & ~i31),
  v310 = (v311 & i32) | (~v305 & ~i32),
  v311 = (~v305 & ~i33) | i33,
  v312 = (v313 & i30) | (v305 & ~i30),
  v313 = (v305 & i31) | (v314 & ~i31),
  v314 = (v315 & i32) | (v305 & ~i32),
  v315 = (v305 & ~i33) | i33,
  v316 = (v317 & i10) | (v302 & ~i10),
  v317 = (v320 & i11) | (v318 & ~i11),
  v318 = (v320 & i12) | (v319 & ~i12),
  v319 = (v329 & i13) | (v320 & ~i13),
  v320 = (v325 & i23) | (v321 & ~i23),
  v321 = (v322 & i30) | (v305 & ~i30),
  v322 = (v305 & i31) | (v323 & ~i31),
  v323 = (v324 & i32) | (v305 & ~i32),
  v324 = v305 & i33,
  v325 = (v326 & i30) | (v305 & ~i30),
  v326 = (v305 & i31) | (v327 & ~i31),
  v327 = (v328 & i32) | (v305 & ~i32),
  v328 = (v305 & i33) | ~i33,
  v329 = (v330 & i14) | (v320 & ~i14),
  v330 = (v338 & i23) | (v331 & ~i23),
  v331 = (v335 & i26) | (v332 & ~i26),
  v332 = (v333 & i30) | (v305 & ~i30),
  v333 = (v305 & i31) | (~v334 & ~i31),
  v334 = (~v305 & ~i32) | i32,
  i100 = \IN-i100 ,
  v335 = (v336 & i30) | (v305 & ~i30),
  i101 = \IN-i101 ,
  v336 = (v305 & i31) | (v337 & ~i31),
  i102 = \IN-i102 ,
  v337 = (v63 & i32) | (v305 & ~i32),
  i103 = \IN-i103 ,
  v338 = (v342 & i26) | (v339 & ~i26),
  i104 = \IN-i104 ,
  v339 = (v340 & i30) | (v305 & ~i30),
  v8600 = (v8373 & i30) | (~v7029 & ~i30),
  i105 = \IN-i105 ,
  v8601 = (v8369 & i13) | (v8602 & ~i13),
  i106 = \IN-i106 ,
  v8602 = (v8615 & i14) | (v8603 & ~i14),
  i107 = \IN-i107 ,
  v8603 = (v8609 & i21) | (v8604 & ~i21),
  i108 = \IN-i108 ,
  v8604 = (v7445 & i23) | (v8605 & ~i23),
  i109 = \IN-i109 ,
  v8605 = (v7445 & i24) | (v8606 & ~i24),
  v8606 = (v8372 & i26) | (v8607 & ~i26),
  v340 = (v305 & i31) | (~v341 & ~i31),
  v8607 = (v8372 & i27) | (v8608 & ~i27),
  v341 = (v63 & i32) | (~v305 & ~i32),
  v8608 = v6430 & i30,
  v342 = (v343 & i30) | (v305 & ~i30),
  v8609 = (v8610 & i22) | (v8604 & ~i22),
  v343 = (v305 & i31) | (v344 & ~i31),
  v344 = (v305 & ~i32) | i32,
  i110 = \IN-i110 ,
  v345 = (v347 & i30) | (v346 & ~i30),
  i111 = \IN-i111 ,
  v346 = i39,
  i112 = \IN-i112 ,
  v347 = (v346 & i31) | (v348 & ~i31),
  i113 = \IN-i113 ,
  v348 = (v346 & i32) | (v63 & ~i32),
  i114 = \IN-i114 ,
  v349 = (v397 & i15) | (v350 & ~i15),
  v8610 = (v7451 & i23) | (v8611 & ~i23),
  i115 = \IN-i115 ,
  v8611 = (v7451 & i24) | (v8612 & ~i24),
  i116 = \IN-i116 ,
  v8612 = (v8377 & i26) | (v8613 & ~i26),
  i117 = \IN-i117 ,
  v8613 = (v8377 & i27) | (v8614 & ~i27),
  i118 = \IN-i118 ,
  v8614 = (v6430 & i30) | (~v6460 & ~i30),
  i119 = \IN-i119 ,
  v8615 = (v8619 & i21) | (v8616 & ~i21),
  v8616 = (v7647 & i23) | (v8617 & ~i23),
  v350 = (v381 & i17) | (v351 & ~i17),
  v8617 = (v7647 & i24) | (v8618 & ~i24),
  v351 = (v369 & i19) | (v352 & ~i19),
  v8618 = (v8608 & i27) | (v8372 & ~i27),
  v352 = (v362 & i20) | (v353 & ~i20),
  v8619 = (v8620 & i22) | (v8616 & ~i22),
  v353 = (v359 & i30) | (v354 & ~i30),
  v354 = (v358 & i36) | (v355 & ~i36),
  i120 = \IN-i120 ,
  v355 = (v357 & i37) | (v356 & ~i37),
  i121 = \IN-i121 ,
  v356 = v346 & i38,
  i122 = \IN-i122 ,
  v357 = i38,
  i123 = \IN-i123 ,
  v358 = v357 & i37,
  i124 = \IN-i124 ,
  v359 = (v361 & i31) | (v360 & ~i31),
  v8620 = (v7650 & i23) | (v8621 & ~i23),
  i125 = \IN-i125 ,
  v8621 = (v7650 & i24) | (v8622 & ~i24),
  i126 = \IN-i126 ,
  v8622 = (v8614 & i27) | (v8377 & ~i27),
  i127 = \IN-i127 ,
  v8623 = (v8369 & i12) | (v8624 & ~i12),
  i128 = \IN-i128 ,
  v8624 = (v8369 & i13) | (v8625 & ~i13),
  i129 = \IN-i129 ,
  v8625 = (v8626 & i14) | (v8369 & ~i14),
  v8626 = (v8630 & i21) | (v8627 & ~i21),
  v360 = (v354 & i32) | ~i32,
  v8627 = (v7791 & i23) | (v8628 & ~i23),
  v361 = v354 & i32,
  v8628 = (v7791 & i24) | (v8629 & ~i24),
  v362 = (v366 & i30) | (v363 & ~i30),
  v8629 = (v8607 & i26) | (v8372 & ~i26),
  v363 = (v358 & i36) | (v364 & ~i36),
  v364 = (v357 & i37) | (~v365 & ~i37),
  i130 = \IN-i130 ,
  v365 = (v346 & i38) | ~i38,
  i131 = \IN-i131 ,
  v366 = (v368 & i31) | (v367 & ~i31),
  i132 = \IN-i132 ,
  v367 = (v363 & i32) | ~i32,
  i133 = \IN-i133 ,
  v368 = v363 & i32,
  i134 = \IN-i134 ,
  v369 = (v376 & i20) | (v370 & ~i20),
  v8630 = (v8631 & i22) | (v8627 & ~i22),
  i135 = \IN-i135 ,
  v8631 = (v7794 & i23) | (v8632 & ~i23),
  i136 = \IN-i136 ,
  v8632 = (v7794 & i24) | (v8633 & ~i24),
  i137 = \IN-i137 ,
  v8633 = (v8613 & i26) | (v8377 & ~i26),
  i138 = \IN-i138 ,
  v8634 = (v8763 & i11) | (v8635 & ~i11),
  i139 = \IN-i139 ,
  v8635 = (v8753 & i12) | (v8636 & ~i12),
  v8636 = (v8638 & i13) | (v8637 & ~i13),
  v370 = (v373 & i30) | (v371 & ~i30),
  v8637 = (v8642 & i14) | (v8638 & ~i14),
  v371 = (v354 & i35) | (v372 & ~i35),
  v8638 = (v8640 & i21) | (v8639 & ~i21),
  v372 = (v358 & i36) | (v357 & ~i36),
  v8639 = (v8372 & i24) | (v6456 & ~i24),
  v373 = (v375 & i31) | (v374 & ~i31),
  v374 = (v371 & i32) | ~i32,
  i140 = \IN-i140 ,
  v375 = v371 & i32,
  i141 = \IN-i141 ,
  v376 = (v378 & i30) | (v377 & ~i30),
  i142 = \IN-i142 ,
  v377 = (v363 & i35) | (v372 & ~i35),
  i143 = \IN-i143 ,
  v378 = (v380 & i31) | (v379 & ~i31),
  i144 = \IN-i144 ,
  v379 = (v377 & i32) | ~i32,
  v8640 = (v8641 & i22) | (v8639 & ~i22),
  i145 = \IN-i145 ,
  v8641 = (v8377 & i24) | (v6459 & ~i24),
  i146 = \IN-i146 ,
  v8642 = (v8698 & i15) | (v8643 & ~i15),
  i147 = \IN-i147 ,
  v8643 = (v8671 & i16) | (v8644 & ~i16),
  i148 = \IN-i148 ,
  v8644 = (v8660 & i17) | (v8645 & ~i17),
  i149 = \IN-i149 ,
  v8645 = (v8653 & i19) | (v8646 & ~i19),
  v8646 = (v8650 & i20) | (v8647 & ~i20),
  v380 = v377 & i32,
  v8647 = (v8648 & i21) | (v8639 & ~i21),
  v381 = (v393 & i19) | (v382 & ~i19),
  v8648 = (v8649 & i22) | (v8639 & ~i22),
  v382 = (v388 & i20) | (v383 & ~i20),
  v8649 = (v8387 & i24) | (v6789 & ~i24),
  v383 = (v385 & i30) | (v384 & ~i30),
  v384 = (v372 & i35) | (v354 & ~i35),
  i150 = \IN-i150 ,
  v385 = (v387 & i31) | (v386 & ~i31),
  i151 = \IN-i151 ,
  v386 = (v384 & i32) | ~i32,
  i152 = \IN-i152 ,
  v387 = v384 & i32,
  i153 = \IN-i153 ,
  v388 = (v390 & i30) | (v389 & ~i30),
  i154 = \IN-i154 ,
  v389 = (v372 & i35) | (v363 & ~i35),
  v8650 = (v8651 & i21) | (v8639 & ~i21),
  i155 = \IN-i155 ,
  v8651 = (v8652 & i22) | (v8639 & ~i22),
  i156 = \IN-i156 ,
  v8652 = (v8394 & i24) | (v6797 & ~i24),
  i157 = \IN-i157 ,
  v8653 = (v8657 & i20) | (v8654 & ~i20),
  i158 = \IN-i158 ,
  v8654 = (v8655 & i21) | (v8639 & ~i21),
  i159 = \IN-i159 ,
  v8655 = (v8656 & i22) | (v8639 & ~i22),
  v8656 = (v8402 & i24) | (v6806 & ~i24),
  v390 = (v392 & i31) | (v391 & ~i31),
  v8657 = (v8658 & i21) | (v8639 & ~i21),
  v391 = (v389 & i32) | ~i32,
  v8658 = (v8659 & i22) | (v8639 & ~i22),
  v392 = v389 & i32,
  v8659 = (v8409 & i24) | (v6814 & ~i24),
  v393 = (v394 & i30) | (v372 & ~i30),
  v394 = (v396 & i31) | (v395 & ~i31),
  i160 = \IN-i160 ,
  v395 = (v372 & i32) | ~i32,
  i161 = \IN-i161 ,
  v396 = v372 & i32,
  i162 = \IN-i162 ,
  v397 = (v421 & i17) | (v398 & ~i17),
  i163 = \IN-i163 ,
  v398 = (v410 & i19) | (v399 & ~i19),
  i164 = \IN-i164 ,
  v399 = (v405 & i20) | (v400 & ~i20),
  v8660 = (v8668 & i19) | (v8661 & ~i19),
  i165 = \IN-i165 ,
  v8661 = (v8665 & i20) | (v8662 & ~i20),
  i166 = \IN-i166 ,
  v8662 = (v8663 & i21) | (v8639 & ~i21),
  i167 = \IN-i167 ,
  v8663 = (v8664 & i22) | (v8639 & ~i22),
  i168 = \IN-i168 ,
  v8664 = (v8418 & i24) | (v6824 & ~i24),
  i169 = \IN-i169 ,
  v8665 = (v8666 & i21) | (v8639 & ~i21),
  v8666 = (v8667 & i22) | (v8639 & ~i22),
  v8667 = (v8425 & i24) | (v6832 & ~i24),
  v8668 = (v8669 & i21) | (v8639 & ~i21),
  v8669 = (v8670 & i22) | (v8639 & ~i22),
  i170 = \IN-i170 ,
  i171 = \IN-i171 ,
  i172 = \IN-i172 ,
  i173 = \IN-i173 ,
  i174 = \IN-i174 ,
  v8670 = (v8432 & i24) | (v6840 & ~i24),
  i175 = \IN-i175 ,
  v8671 = (v8687 & i17) | (v8672 & ~i17),
  i176 = \IN-i176 ,
  v8672 = (v8680 & i19) | (v8673 & ~i19),
  i177 = \IN-i177 ,
  v8673 = (v8677 & i20) | (v8674 & ~i20),
  i178 = \IN-i178 ,
  v8674 = (v8675 & i21) | (v8639 & ~i21),
  i179 = \IN-i179 ,
  v8675 = (v8676 & i22) | (v8639 & ~i22),
  v8676 = (v8442 & i24) | (v6851 & ~i24),
  v8677 = (v8678 & i21) | (v8639 & ~i21),
  v8678 = (v8679 & i22) | (v8639 & ~i22),
  v8679 = (v8449 & i24) | (v6859 & ~i24),
  i180 = \IN-i180 ,
  i181 = \IN-i181 ,
  i182 = \IN-i182 ,
  i183 = \IN-i183 ,
  i184 = \IN-i184 ,
  v8680 = (v8684 & i20) | (v8681 & ~i20),
  i185 = \IN-i185 ,
  v8681 = (v8682 & i21) | (v8639 & ~i21),
  i186 = \IN-i186 ,
  v8682 = (v8683 & i22) | (v8639 & ~i22),
  i187 = \IN-i187 ,
  v8683 = (v8457 & i24) | (v6868 & ~i24),
  i188 = \IN-i188 ,
  v8684 = (v8685 & i21) | (v8639 & ~i21),
  i189 = \IN-i189 ,
  v8685 = (v8686 & i22) | (v8639 & ~i22),
  v8686 = (v8464 & i24) | (v6876 & ~i24),
  v8687 = (v8695 & i19) | (v8688 & ~i19),
  v8688 = (v8692 & i20) | (v8689 & ~i20),
  v8689 = (v8690 & i21) | (v8639 & ~i21),
  i190 = \IN-i190 ,
  i191 = \IN-i191 ,
  i192 = \IN-i192 ,
  i193 = \IN-i193 ,
  i194 = \IN-i194 ,
  v8690 = (v8691 & i22) | (v8639 & ~i22),
  i195 = \IN-i195 ,
  v8691 = (v8473 & i24) | (v6886 & ~i24),
  i196 = \IN-i196 ,
  v8692 = (v8693 & i21) | (v8639 & ~i21),
  i197 = \IN-i197 ,
  v8693 = (v8694 & i22) | (v8639 & ~i22),
  i198 = \IN-i198 ,
  v8694 = (v8480 & i24) | (v6894 & ~i24),
  i199 = \IN-i199 ,
  v8695 = (v8696 & i21) | (v8639 & ~i21),
  v8696 = (v8697 & i22) | (v8639 & ~i22),
  v8697 = (v8487 & i24) | (v6902 & ~i24),
  v8698 = (v8726 & i16) | (v8699 & ~i16),
  v8699 = (v8715 & i17) | (v8700 & ~i17),
  v400 = (v402 & i30) | (v401 & ~i30),
  v401 = (v357 & i36) | (v355 & ~i36),
  v402 = (v404 & i31) | (v403 & ~i31),
  v403 = (v401 & i32) | ~i32,
  v404 = v401 & i32,
  v405 = (v407 & i30) | (v406 & ~i30),
  v406 = (v357 & i36) | (v364 & ~i36),
  v407 = (v409 & i31) | (v408 & ~i31),
  v408 = (v406 & i32) | ~i32,
  v409 = v406 & i32,
  v410 = (v416 & i20) | (v411 & ~i20),
  v411 = (v413 & i30) | (v412 & ~i30),
  v412 = (v401 & i35) | (v357 & ~i35),
  v413 = (v415 & i31) | (v414 & ~i31),
  v414 = (v412 & i32) | ~i32,
  v415 = v412 & i32,
  v416 = (v418 & i30) | (v417 & ~i30),
  v417 = (v406 & i35) | (v357 & ~i35),
  v418 = (v420 & i31) | (v419 & ~i31),
  v419 = (v417 & i32) | ~i32,
  v420 = v417 & i32,
  v421 = (v433 & i19) | (v422 & ~i19),
  v422 = (v428 & i20) | (v423 & ~i20),
  v423 = (v425 & i30) | (v424 & ~i30),
  v424 = (v357 & i35) | (v401 & ~i35),
  v425 = (v427 & i31) | (v426 & ~i31),
  v426 = (v424 & i32) | ~i32,
  v427 = v424 & i32,
  v428 = (v430 & i30) | (v429 & ~i30),
  v429 = (v357 & i35) | (v406 & ~i35),
  v430 = (v432 & i31) | (v431 & ~i31),
  v431 = (v429 & i32) | ~i32,
  v432 = v429 & i32,
  v433 = (v434 & i30) | (v357 & ~i30),
  v434 = (v436 & i31) | (v435 & ~i31),
  i200 = \IN-i200 ,
  v435 = (v357 & i32) | ~i32,
  i201 = \IN-i201 ,
  v436 = v357 & i32,
  i202 = \IN-i202 ,
  v437 = (v476 & i15) | (v438 & ~i15),
  i203 = \IN-i203 ,
  v438 = (v440 & i17) | (v439 & ~i17),
  i204 = \IN-i204 ,
  v439 = (v455 & i18) | (v440 & ~i18),
  v8700 = (v8708 & i19) | (v8701 & ~i19),
  i205 = \IN-i205 ,
  v8701 = (v8705 & i20) | (v8702 & ~i20),
  i206 = \IN-i206 ,
  v8702 = (v8703 & i21) | (v8639 & ~i21),
  i207 = \IN-i207 ,
  v8703 = (v8704 & i22) | (v8639 & ~i22),
  i208 = \IN-i208 ,
  v8704 = (v8498 & i24) | (v6914 & ~i24),
  i209 = \IN-i209 ,
  v8705 = (v8706 & i21) | (v8639 & ~i21),
  v8706 = (v8707 & i22) | (v8639 & ~i22),
  v440 = (v448 & i30) | (v441 & ~i30),
  v8707 = (v8505 & i24) | (v6922 & ~i24),
  v441 = (v447 & i36) | (v442 & ~i36),
  v8708 = (v8712 & i20) | (v8709 & ~i20),
  v442 = v443 & i37,
  v8709 = (v8710 & i21) | (v8639 & ~i21),
  v443 = (v444 & i38) | ~i38,
  v444 = (v446 & i39) | (~v445 & ~i39),
  i210 = \IN-i210 ,
  v445 = (v60 & i42) | (v80 & ~i42),
  i211 = \IN-i211 ,
  v446 = (v60 & i42) | (v71 & ~i42),
  i212 = \IN-i212 ,
  v447 = (v443 & i37) | (v357 & ~i37),
  i213 = \IN-i213 ,
  v448 = (v454 & i31) | (v449 & ~i31),
  i214 = \IN-i214 ,
  v449 = (v450 & i32) | (v444 & ~i32),
  v8710 = (v8711 & i22) | (v8639 & ~i22),
  i215 = \IN-i215 ,
  v8711 = (v8513 & i24) | (v6931 & ~i24),
  i216 = \IN-i216 ,
  v8712 = (v8713 & i21) | (v8639 & ~i21),
  i217 = \IN-i217 ,
  v8713 = (v8714 & i22) | (v8639 & ~i22),
  i218 = \IN-i218 ,
  v8714 = (v8520 & i24) | (v6939 & ~i24),
  i219 = \IN-i219 ,
  v8715 = (v8723 & i19) | (v8716 & ~i19),
  v8716 = (v8720 & i20) | (v8717 & ~i20),
  v450 = (v453 & i36) | (v451 & ~i36),
  v8717 = (v8718 & i21) | (v8639 & ~i21),
  v451 = v452 & i37,
  v8718 = (v8719 & i22) | (v8639 & ~i22),
  v452 = (v172 & i38) | ~i38,
  v8719 = (v8529 & i24) | (v6949 & ~i24),
  v453 = (v452 & i37) | (v357 & ~i37),
  v454 = v450 & i32,
  i220 = \IN-i220 ,
  v455 = (v466 & i20) | (v456 & ~i20),
  i221 = \IN-i221 ,
  v456 = (v460 & i30) | (v457 & ~i30),
  i222 = \IN-i222 ,
  v457 = (v458 & i35) | (v441 & ~i35),
  i223 = \IN-i223 ,
  v458 = (v447 & i36) | (v459 & ~i36),
  i224 = \IN-i224 ,
  v459 = (v443 & i37) | (~v365 & ~i37),
  v8720 = (v8721 & i21) | (v8639 & ~i21),
  i225 = \IN-i225 ,
  v8721 = (v8722 & i22) | (v8639 & ~i22),
  i226 = \IN-i226 ,
  v8722 = (v8536 & i24) | (v6957 & ~i24),
  i227 = \IN-i227 ,
  v8723 = (v8724 & i21) | (v8639 & ~i21),
  i228 = \IN-i228 ,
  v8724 = (v8725 & i22) | (v8639 & ~i22),
  i229 = \IN-i229 ,
  v8725 = (v8543 & i24) | (v6965 & ~i24),
  v8726 = (v8742 & i17) | (v8727 & ~i17),
  v460 = (v465 & i31) | (v461 & ~i31),
  v8727 = (v8735 & i19) | (v8728 & ~i19),
  v461 = (v462 & i32) | (v444 & ~i32),
  v8728 = (v8732 & i20) | (v8729 & ~i20),
  v462 = (v463 & i35) | (v450 & ~i35),
  v8729 = (v8730 & i21) | (v8639 & ~i21),
  v463 = (v453 & i36) | (v464 & ~i36),
  v464 = (v452 & i37) | (~v365 & ~i37),
  i230 = \IN-i230 ,
  v465 = v462 & i32,
  i231 = \IN-i231 ,
  v466 = (v470 & i30) | (v467 & ~i30),
  i232 = \IN-i232 ,
  v467 = (v468 & i35) | (v441 & ~i35),
  i233 = \IN-i233 ,
  v468 = (v447 & i36) | (v469 & ~i36),
  i234 = \IN-i234 ,
  v469 = (v443 & i37) | (v356 & ~i37),
  v8730 = (v8731 & i22) | (v8639 & ~i22),
  i235 = \IN-i235 ,
  v8731 = (v8553 & i24) | (v6976 & ~i24),
  i236 = \IN-i236 ,
  v8732 = (v8733 & i21) | (v8639 & ~i21),
  i237 = \IN-i237 ,
  v8733 = (v8734 & i22) | (v8639 & ~i22),
  i238 = \IN-i238 ,
  v8734 = (v8560 & i24) | (v6984 & ~i24),
  i239 = \IN-i239 ,
  v8735 = (v8739 & i20) | (v8736 & ~i20),
  v8736 = (v8737 & i21) | (v8639 & ~i21),
  v470 = (v475 & i31) | (v471 & ~i31),
  v8737 = (v8738 & i22) | (v8639 & ~i22),
  v471 = (v472 & i32) | (v444 & ~i32),
  v8738 = (v8568 & i24) | (v6993 & ~i24),
  v472 = (v473 & i35) | (v450 & ~i35),
  v8739 = (v8740 & i21) | (v8639 & ~i21),
  v473 = (v453 & i36) | (v474 & ~i36),
  v474 = (v452 & i37) | (v356 & ~i37),
  i240 = \IN-i240 ,
  v475 = v472 & i32,
  i241 = \IN-i241 ,
  v476 = (v478 & i17) | (v477 & ~i17),
  i242 = \IN-i242 ,
  v477 = (v482 & i18) | (v478 & ~i18),
  i243 = \IN-i243 ,
  v478 = (v479 & i30) | (v442 & ~i30),
  i244 = \IN-i244 ,
  v479 = (v481 & i31) | (v480 & ~i31),
  v8740 = (v8741 & i22) | (v8639 & ~i22),
  i245 = \IN-i245 ,
  v8741 = (v8575 & i24) | (v7001 & ~i24),
  i246 = \IN-i246 ,
  v8742 = (v8750 & i19) | (v8743 & ~i19),
  i247 = \IN-i247 ,
  v8743 = (v8747 & i20) | (v8744 & ~i20),
  i248 = \IN-i248 ,
  v8744 = (v8745 & i21) | (v8639 & ~i21),
  i249 = \IN-i249 ,
  v8745 = (v8746 & i22) | (v8639 & ~i22),
  v8746 = (v8584 & i24) | (v7011 & ~i24),
  v480 = (v451 & i32) | (v444 & ~i32),
  v8747 = (v8748 & i21) | (v8639 & ~i21),
  v481 = v451 & i32,
  v8748 = (v8749 & i22) | (v8639 & ~i22),
  v482 = (v491 & i20) | (v483 & ~i20),
  v8749 = (v8591 & i24) | (v7019 & ~i24),
  v483 = (v486 & i30) | (v484 & ~i30),
  v484 = (v485 & i35) | (v442 & ~i35),
  i250 = \IN-i250 ,
  v485 = (v442 & i36) | (v459 & ~i36),
  i251 = \IN-i251 ,
  v486 = (v490 & i31) | (v487 & ~i31),
  i252 = \IN-i252 ,
  v487 = (v488 & i32) | (v444 & ~i32),
  i253 = \IN-i253 ,
  v488 = (v489 & i35) | (v451 & ~i35),
  i254 = \IN-i254 ,
  v489 = (v451 & i36) | (v464 & ~i36),
  v8750 = (v8751 & i21) | (v8639 & ~i21),
  i255 = \IN-i255 ,
  v8751 = (v8752 & i22) | (v8639 & ~i22),
  i256 = \IN-i256 ,
  v8752 = (v8598 & i24) | (v7027 & ~i24),
  i257 = \IN-i257 ,
  v8753 = (v8638 & i13) | (v8754 & ~i13),
  i258 = \IN-i258 ,
  v8754 = (v8759 & i14) | (v8755 & ~i14),
  i259 = \IN-i259 ,
  v8755 = (v8757 & i21) | (v8756 & ~i21),
  v8756 = (v8606 & i24) | (v7445 & ~i24),
  v490 = v488 & i32,
  v8757 = (v8758 & i22) | (v8756 & ~i22),
  v491 = (v494 & i30) | (v492 & ~i30),
  v8758 = (v8612 & i24) | (v7451 & ~i24),
  v492 = (v493 & i35) | (v442 & ~i35),
  v8759 = (v8761 & i21) | (v8760 & ~i21),
  v493 = (v442 & i36) | (v469 & ~i36),
  v494 = (v498 & i31) | (v495 & ~i31),
  i260 = \IN-i260 ,
  v495 = (v496 & i32) | (v444 & ~i32),
  i261 = \IN-i261 ,
  v496 = (v497 & i35) | (v451 & ~i35),
  i262 = \IN-i262 ,
  v497 = (v451 & i36) | (v474 & ~i36),
  i263 = \IN-i263 ,
  v498 = v496 & i32,
  i264 = \IN-i264 ,
  v499 = (v510 & i2) | (v500 & ~i2),
  v8760 = (v8618 & i24) | (v7647 & ~i24),
  i265 = \IN-i265 ,
  v8761 = (v8762 & i22) | (v8760 & ~i22),
  i266 = \IN-i266 ,
  v8762 = (v8622 & i24) | (v7650 & ~i24),
  i267 = \IN-i267 ,
  v8763 = (v8638 & i12) | (v8764 & ~i12),
  i268 = \IN-i268 ,
  v8764 = (v8638 & i13) | (v8765 & ~i13),
  i269 = \IN-i269 ,
  v8765 = (v8766 & i14) | (v8638 & ~i14),
  v8766 = (v8768 & i21) | (v8767 & ~i21),
  v8767 = (v8629 & i24) | (v7791 & ~i24),
  v8768 = (v8769 & i22) | (v8767 & ~i22),
  v8769 = (v8633 & i24) | (v7794 & ~i24),
  i270 = \IN-i270 ,
  i271 = \IN-i271 ,
  i272 = \IN-i272 ,
  i273 = \IN-i273 ,
  i274 = \IN-i274 ,
  v8770 = (v8350 & i8) | (v8771 & ~i8),
  i275 = \IN-i275 ,
  v8771 = (v8350 & i9) | (v8772 & ~i9),
  i276 = \IN-i276 ,
  v8772 = (v8773 & i10) | (v8350 & ~i10),
  i277 = \IN-i277 ,
  v8773 = (v8902 & i11) | (v8774 & ~i11),
  i278 = \IN-i278 ,
  v8774 = (v8892 & i12) | (v8775 & ~i12),
  i279 = \IN-i279 ,
  v8775 = (v8777 & i13) | (v8776 & ~i13),
  v8776 = (v8781 & i14) | (v8777 & ~i14),
  v8777 = (v8779 & i21) | (v8778 & ~i21),
  v8778 = (v8371 & i23) | (v6456 & ~i23),
  v8779 = (v8780 & i22) | (v8778 & ~i22),
  i280 = \IN-i280 ,
  i281 = \IN-i281 ,
  i282 = \IN-i282 ,
  i283 = \IN-i283 ,
  i284 = \IN-i284 ,
  v8780 = (v8376 & i23) | (v6459 & ~i23),
  i285 = \IN-i285 ,
  v8781 = (v8837 & i15) | (v8782 & ~i15),
  i286 = \IN-i286 ,
  v8782 = (v8810 & i16) | (v8783 & ~i16),
  i287 = \IN-i287 ,
  v8783 = (v8799 & i17) | (v8784 & ~i17),
  i288 = \IN-i288 ,
  v8784 = (v8792 & i19) | (v8785 & ~i19),
  i289 = \IN-i289 ,
  v8785 = (v8789 & i20) | (v8786 & ~i20),
  v8786 = (v8787 & i21) | (v8778 & ~i21),
  v8787 = (v8788 & i22) | (v8778 & ~i22),
  v8788 = (v8386 & i23) | (v6789 & ~i23),
  v8789 = (v8790 & i21) | (v8778 & ~i21),
  i290 = \IN-i290 ,
  i291 = \IN-i291 ,
  i292 = \IN-i292 ,
  i293 = \IN-i293 ,
  i294 = \IN-i294 ,
  v8790 = (v8791 & i22) | (v8778 & ~i22),
  i295 = \IN-i295 ,
  v8791 = (v8393 & i23) | (v6797 & ~i23),
  i296 = \IN-i296 ,
  v8792 = (v8796 & i20) | (v8793 & ~i20),
  i297 = \IN-i297 ,
  v8793 = (v8794 & i21) | (v8778 & ~i21),
  i298 = \IN-i298 ,
  v8794 = (v8795 & i22) | (v8778 & ~i22),
  i299 = \IN-i299 ,
  v8795 = (v8401 & i23) | (v6806 & ~i23),
  v8796 = (v8797 & i21) | (v8778 & ~i21),
  v8797 = (v8798 & i22) | (v8778 & ~i22),
  v8798 = (v8408 & i23) | (v6814 & ~i23),
  v8799 = (v8807 & i19) | (v8800 & ~i19),
  v500 = (v510 & i3) | (v501 & ~i3),
  v501 = (v510 & i4) | (v502 & ~i4),
  v502 = (v510 & i5) | (v503 & ~i5),
  v503 = (v510 & i6) | (v504 & ~i6),
  v504 = (v507 & i7) | (v505 & ~i7),
  v505 = (v507 & i8) | (v506 & ~i8),
  v506 = (v521 & i9) | (v507 & ~i9),
  v507 = (v510 & i11) | (v508 & ~i11),
  v508 = (v510 & i12) | (v509 & ~i12),
  v509 = (v511 & i13) | (v510 & ~i13),
  v510 = i36,
  v511 = (v512 & i14) | (v510 & ~i14),
  v512 = (v517 & i27) | (v513 & ~i27),
  v513 = (v514 & i30) | (v510 & ~i30),
  v514 = (v510 & i31) | (v515 & ~i31),
  v515 = (v510 & i32) | (~v516 & ~i32),
  v516 = (~v510 & ~i33) | i33,
  v517 = (v518 & i30) | (v510 & ~i30),
  v518 = (v510 & i31) | (v519 & ~i31),
  v519 = (v510 & i32) | (v520 & ~i32),
  v520 = (v510 & ~i33) | i33,
  v521 = (v522 & i10) | (v507 & ~i10),
  v522 = (v525 & i11) | (v523 & ~i11),
  v523 = (v525 & i12) | (v524 & ~i12),
  v524 = (v534 & i13) | (v525 & ~i13),
  v525 = (v530 & i24) | (v526 & ~i24),
  v526 = (v527 & i30) | (v510 & ~i30),
  v527 = (v510 & i31) | (v528 & ~i31),
  v528 = (v510 & i32) | (v529 & ~i32),
  v529 = v510 & i33,
  v530 = (v531 & i30) | (v510 & ~i30),
  v531 = (v510 & i31) | (v532 & ~i31),
  v532 = (v510 & i32) | (v533 & ~i32),
  v533 = (v510 & i33) | ~i33,
  v534 = (v535 & i14) | (v525 & ~i14),
  i300 = \IN-i300 ,
  v535 = (v543 & i24) | (v536 & ~i24),
  i301 = \IN-i301 ,
  v536 = (v540 & i27) | (v537 & ~i27),
  i302 = \IN-i302 ,
  v537 = (v538 & i30) | (v510 & ~i30),
  i303 = \IN-i303 ,
  v538 = (v510 & i31) | (v539 & ~i31),
  i304 = \IN-i304 ,
  v539 = v510 & i32,
  v8800 = (v8804 & i20) | (v8801 & ~i20),
  i305 = \IN-i305 ,
  v8801 = (v8802 & i21) | (v8778 & ~i21),
  i306 = \IN-i306 ,
  v8802 = (v8803 & i22) | (v8778 & ~i22),
  i307 = \IN-i307 ,
  v8803 = (v8417 & i23) | (v6824 & ~i23),
  i308 = \IN-i308 ,
  v8804 = (v8805 & i21) | (v8778 & ~i21),
  i309 = \IN-i309 ,
  v8805 = (v8806 & i22) | (v8778 & ~i22),
  v8806 = (v8424 & i23) | (v6832 & ~i23),
  v540 = (v541 & i30) | (v510 & ~i30),
  v8807 = (v8808 & i21) | (v8778 & ~i21),
  v541 = (v510 & i31) | (v542 & ~i31),
  v8808 = (v8809 & i22) | (v8778 & ~i22),
  v542 = (v510 & i32) | (v63 & ~i32),
  v8809 = (v8431 & i23) | (v6840 & ~i23),
  v543 = (v547 & i27) | (v544 & ~i27),
  v544 = (v545 & i30) | (v510 & ~i30),
  i310 = \IN-i310 ,
  v545 = (v510 & i31) | (v546 & ~i31),
  i311 = \IN-i311 ,
  v546 = (v510 & i32) | (~v63 & ~i32),
  i312 = \IN-i312 ,
  v547 = (v548 & i30) | (v510 & ~i30),
  i313 = \IN-i313 ,
  v548 = (v510 & i31) | (v549 & ~i31),
  i314 = \IN-i314 ,
  v549 = (v510 & i32) | ~i32,
  v8810 = (v8826 & i17) | (v8811 & ~i17),
  i315 = \IN-i315 ,
  v8811 = (v8819 & i19) | (v8812 & ~i19),
  i316 = \IN-i316 ,
  v8812 = (v8816 & i20) | (v8813 & ~i20),
  i317 = \IN-i317 ,
  v8813 = (v8814 & i21) | (v8778 & ~i21),
  i318 = \IN-i318 ,
  v8814 = (v8815 & i22) | (v8778 & ~i22),
  i319 = \IN-i319 ,
  v8815 = (v8441 & i23) | (v6851 & ~i23),
  v8816 = (v8817 & i21) | (v8778 & ~i21),
  v550 = (v561 & i2) | (v551 & ~i2),
  v8817 = (v8818 & i22) | (v8778 & ~i22),
  v551 = (v561 & i3) | (v552 & ~i3),
  v8818 = (v8448 & i23) | (v6859 & ~i23),
  v552 = (v561 & i4) | (v553 & ~i4),
  v8819 = (v8823 & i20) | (v8820 & ~i20),
  v553 = (v561 & i5) | (v554 & ~i5),
  v554 = (v561 & i6) | (v555 & ~i6),
  i320 = \IN-i320 ,
  v555 = (v558 & i7) | (v556 & ~i7),
  i321 = \IN-i321 ,
  v556 = (v558 & i8) | (v557 & ~i8),
  i322 = \IN-i322 ,
  v557 = (v572 & i9) | (v558 & ~i9),
  i323 = \IN-i323 ,
  v558 = (v561 & i11) | (v559 & ~i11),
  i324 = \IN-i324 ,
  v559 = (v561 & i12) | (v560 & ~i12),
  v8820 = (v8821 & i21) | (v8778 & ~i21),
  i325 = \IN-i325 ,
  v8821 = (v8822 & i22) | (v8778 & ~i22),
  i326 = \IN-i326 ,
  v8822 = (v8456 & i23) | (v6868 & ~i23),
  i327 = \IN-i327 ,
  v8823 = (v8824 & i21) | (v8778 & ~i21),
  i328 = \IN-i328 ,
  v8824 = (v8825 & i22) | (v8778 & ~i22),
  i329 = \IN-i329 ,
  v8825 = (v8463 & i23) | (v6876 & ~i23),
  v8826 = (v8834 & i19) | (v8827 & ~i19),
  v560 = (v562 & i13) | (v561 & ~i13),
  v8827 = (v8831 & i20) | (v8828 & ~i20),
  v561 = i35,
  v8828 = (v8829 & i21) | (v8778 & ~i21),
  v562 = (v563 & i14) | (v561 & ~i14),
  v8829 = (v8830 & i22) | (v8778 & ~i22),
  v563 = (v568 & i26) | (v564 & ~i26),
  v564 = (v565 & i30) | (v561 & ~i30),
  i330 = \IN-i330 ,
  v565 = (v561 & i31) | (v566 & ~i31),
  i331 = \IN-i331 ,
  v566 = (v561 & i32) | (~v567 & ~i32),
  i332 = \IN-i332 ,
  v567 = (~v561 & ~i33) | i33,
  i333 = \IN-i333 ,
  v568 = (v569 & i30) | (v561 & ~i30),
  i334 = \IN-i334 ,
  v569 = (v561 & i31) | (v570 & ~i31),
  v8830 = (v8472 & i23) | (v6886 & ~i23),
  i335 = \IN-i335 ,
  v8831 = (v8832 & i21) | (v8778 & ~i21),
  i336 = \IN-i336 ,
  v8832 = (v8833 & i22) | (v8778 & ~i22),
  i337 = \IN-i337 ,
  v8833 = (v8479 & i23) | (v6894 & ~i23),
  i338 = \IN-i338 ,
  v8834 = (v8835 & i21) | (v8778 & ~i21),
  i339 = \IN-i339 ,
  v8835 = (v8836 & i22) | (v8778 & ~i22),
  v8836 = (v8486 & i23) | (v6902 & ~i23),
  v570 = (v561 & i32) | (v571 & ~i32),
  v8837 = (v8865 & i16) | (v8838 & ~i16),
  v571 = (v561 & ~i33) | i33,
  v8838 = (v8854 & i17) | (v8839 & ~i17),
  v572 = (v573 & i10) | (v558 & ~i10),
  v8839 = (v8847 & i19) | (v8840 & ~i19),
  v573 = (v576 & i11) | (v574 & ~i11),
  v574 = (v576 & i12) | (v575 & ~i12),
  i340 = \IN-i340 ,
  v575 = (v585 & i13) | (v576 & ~i13),
  i341 = \IN-i341 ,
  v576 = (v581 & i23) | (v577 & ~i23),
  i342 = \IN-i342 ,
  v577 = (v578 & i30) | (v561 & ~i30),
  i343 = \IN-i343 ,
  v578 = (v561 & i31) | (v579 & ~i31),
  i344 = \IN-i344 ,
  v579 = (v561 & i32) | (v580 & ~i32),
  v8840 = (v8844 & i20) | (v8841 & ~i20),
  i345 = \IN-i345 ,
  v8841 = (v8842 & i21) | (v8778 & ~i21),
  i346 = \IN-i346 ,
  v8842 = (v8843 & i22) | (v8778 & ~i22),
  i347 = \IN-i347 ,
  v8843 = (v8497 & i23) | (v6914 & ~i23),
  i348 = \IN-i348 ,
  v8844 = (v8845 & i21) | (v8778 & ~i21),
  i349 = \IN-i349 ,
  v8845 = (v8846 & i22) | (v8778 & ~i22),
  v8846 = (v8504 & i23) | (v6922 & ~i23),
  v580 = v561 & i33,
  v8847 = (v8851 & i20) | (v8848 & ~i20),
  v581 = (v582 & i30) | (v561 & ~i30),
  v8848 = (v8849 & i21) | (v8778 & ~i21),
  v582 = (v561 & i31) | (v583 & ~i31),
  v8849 = (v8850 & i22) | (v8778 & ~i22),
  v583 = (v561 & i32) | (v584 & ~i32),
  v584 = (v561 & i33) | ~i33,
  i350 = \IN-i350 ,
  v585 = (v586 & i14) | (v576 & ~i14),
  i351 = \IN-i351 ,
  v586 = (v594 & i23) | (v587 & ~i23),
  i352 = \IN-i352 ,
  v587 = (v591 & i26) | (v588 & ~i26),
  i353 = \IN-i353 ,
  v588 = (v589 & i30) | (v561 & ~i30),
  i354 = \IN-i354 ,
  v589 = (v561 & i31) | (v590 & ~i31),
  v8850 = (v8512 & i23) | (v6931 & ~i23),
  i355 = \IN-i355 ,
  v8851 = (v8852 & i21) | (v8778 & ~i21),
  i356 = \IN-i356 ,
  v8852 = (v8853 & i22) | (v8778 & ~i22),
  i357 = \IN-i357 ,
  v8853 = (v8519 & i23) | (v6939 & ~i23),
  i358 = \IN-i358 ,
  v8854 = (v8862 & i19) | (v8855 & ~i19),
  i359 = \IN-i359 ,
  v8855 = (v8859 & i20) | (v8856 & ~i20),
  v8856 = (v8857 & i21) | (v8778 & ~i21),
  v590 = v561 & i32,
  v8857 = (v8858 & i22) | (v8778 & ~i22),
  v591 = (v592 & i30) | (v561 & ~i30),
  v8858 = (v8528 & i23) | (v6949 & ~i23),
  v592 = (v561 & i31) | (v593 & ~i31),
  v8859 = (v8860 & i21) | (v8778 & ~i21),
  v593 = (v561 & i32) | (v63 & ~i32),
  v594 = (v598 & i26) | (v595 & ~i26),
  i360 = \IN-i360 ,
  v595 = (v596 & i30) | (v561 & ~i30),
  i361 = \IN-i361 ,
  v596 = (v561 & i31) | (v597 & ~i31),
  i362 = \IN-i362 ,
  v597 = (v561 & i32) | (~v63 & ~i32),
  i363 = \IN-i363 ,
  v598 = (v599 & i30) | (v561 & ~i30),
  i364 = \IN-i364 ,
  v599 = (v561 & i31) | (v600 & ~i31),
  v8860 = (v8861 & i22) | (v8778 & ~i22),
  i365 = \IN-i365 ,
  v8861 = (v8535 & i23) | (v6957 & ~i23),
  i366 = \IN-i366 ,
  v8862 = (v8863 & i21) | (v8778 & ~i21),
  i367 = \IN-i367 ,
  v8863 = (v8864 & i22) | (v8778 & ~i22),
  i368 = \IN-i368 ,
  v8864 = (v8542 & i23) | (v6965 & ~i23),
  i369 = \IN-i369 ,
  v8865 = (v8881 & i17) | (v8866 & ~i17),
  v8866 = (v8874 & i19) | (v8867 & ~i19),
  v8867 = (v8871 & i20) | (v8868 & ~i20),
  v8868 = (v8869 & i21) | (v8778 & ~i21),
  v8869 = (v8870 & i22) | (v8778 & ~i22),
  i370 = \IN-i370 ,
  i371 = \IN-i371 ,
  i372 = \IN-i372 ,
  i373 = \IN-i373 ,
  i374 = \IN-i374 ,
  v8870 = (v8552 & i23) | (v6976 & ~i23),
  i375 = \IN-i375 ,
  v8871 = (v8872 & i21) | (v8778 & ~i21),
  i376 = \IN-i376 ,
  v8872 = (v8873 & i22) | (v8778 & ~i22),
  i377 = \IN-i377 ,
  v8873 = (v8559 & i23) | (v6984 & ~i23),
  i378 = \IN-i378 ,
  v8874 = (v8878 & i20) | (v8875 & ~i20),
  i379 = \IN-i379 ,
  v8875 = (v8876 & i21) | (v8778 & ~i21),
  v8876 = (v8877 & i22) | (v8778 & ~i22),
  v8877 = (v8567 & i23) | (v6993 & ~i23),
  v8878 = (v8879 & i21) | (v8778 & ~i21),
  v8879 = (v8880 & i22) | (v8778 & ~i22),
  i380 = \IN-i380 ,
  i381 = \IN-i381 ,
  i382 = \IN-i382 ,
  i383 = \IN-i383 ,
  i384 = \IN-i384 ,
  v8880 = (v8574 & i23) | (v7001 & ~i23),
  i385 = \IN-i385 ,
  v8881 = (v8889 & i19) | (v8882 & ~i19),
  i386 = \IN-i386 ,
  v8882 = (v8886 & i20) | (v8883 & ~i20),
  i387 = \IN-i387 ,
  v8883 = (v8884 & i21) | (v8778 & ~i21),
  i388 = \IN-i388 ,
  v8884 = (v8885 & i22) | (v8778 & ~i22),
  i389 = \IN-i389 ,
  v8885 = (v8583 & i23) | (v7011 & ~i23),
  v8886 = (v8887 & i21) | (v8778 & ~i21),
  v8887 = (v8888 & i22) | (v8778 & ~i22),
  v8888 = (v8590 & i23) | (v7019 & ~i23),
  v8889 = (v8890 & i21) | (v8778 & ~i21),
  i390 = \IN-i390 ,
  i391 = \IN-i391 ,
  i392 = \IN-i392 ,
  i393 = \IN-i393 ,
  i394 = \IN-i394 ,
  v8890 = (v8891 & i22) | (v8778 & ~i22),
  i395 = \IN-i395 ,
  v8891 = (v8597 & i23) | (v7027 & ~i23),
  i396 = \IN-i396 ,
  v8892 = (v8777 & i13) | (v8893 & ~i13),
  i397 = \IN-i397 ,
  v8893 = (v8898 & i14) | (v8894 & ~i14),
  i398 = \IN-i398 ,
  v8894 = (v8896 & i21) | (v8895 & ~i21),
  i399 = \IN-i399 ,
  v8895 = (v8605 & i23) | (v7445 & ~i23),
  v8896 = (v8897 & i22) | (v8895 & ~i22),
  v8897 = (v8611 & i23) | (v7451 & ~i23),
  v8898 = (v8900 & i21) | (v8899 & ~i21),
  v8899 = (v8617 & i23) | (v7647 & ~i23),
  v600 = (v561 & i32) | ~i32,
  v601 = (v617 & i2) | (v602 & ~i2),
  v602 = (v617 & i3) | (v603 & ~i3),
  v603 = (v2066 & i7) | (v604 & ~i7),
  v604 = (v2066 & i8) | (v605 & ~i8),
  v605 = (v2066 & i9) | (v606 & ~i9),
  v606 = (v1616 & i10) | (v607 & ~i10),
  v607 = (v611 & i11) | (v608 & ~i11),
  v608 = (v611 & i12) | (v609 & ~i12),
  v609 = (v611 & i13) | (v610 & ~i13),
  v610 = (v1001 & i14) | (v611 & ~i14),
  v611 = (v862 & i15) | (v612 & ~i15),
  v612 = (v744 & i16) | (v613 & ~i16),
  v613 = (v694 & i17) | (v614 & ~i17),
  v614 = (v654 & i19) | (v615 & ~i19),
  v615 = (v637 & i20) | (v616 & ~i20),
  v616 = (v618 & i21) | (v617 & ~i21),
  v617 = i34,
  v618 = (v619 & i22) | (v617 & ~i22),
  v619 = (v620 & i25) | (v617 & ~i25),
  v620 = (v617 & i30) | (v621 & ~i30),
  v621 = (v617 & i31) | (v622 & ~i31),
  v622 = (v617 & i32) | (v623 & ~i32),
  v623 = (~v624 & ~i34) | i34,
  v624 = (v636 & i36) | (v625 & ~i36),
  v625 = (v635 & i37) | (v626 & ~i37),
  v626 = (v628 & i38) | (v627 & ~i38),
  v627 = (v633 & i39) | (v628 & ~i39),
  v628 = (v629 & ~i41) | i41,
  v629 = (v630 & ~i42) | i42,
  v630 = (v631 & ~i43) | i43,
  v631 = (v632 & i44) | ~i44,
  v632 = (v20 & ~i45) | i45,
  v633 = (v634 & i42) | (v632 & ~i42),
  v634 = (v632 & i43) | ~i43,
  i400 = \IN-i400 ,
  v635 = (v628 & i38) | ~i38,
  i401 = \IN-i401 ,
  v636 = (v635 & i37) | (v628 & ~i37),
  i402 = \IN-i402 ,
  v637 = (v638 & i21) | (v617 & ~i21),
  i403 = \IN-i403 ,
  v638 = (v639 & i22) | (v617 & ~i22),
  i404 = \IN-i404 ,
  v639 = (v640 & i25) | (v617 & ~i25),
  v8900 = (v8901 & i22) | (v8899 & ~i22),
  i405 = \IN-i405 ,
  v8901 = (v8621 & i23) | (v7650 & ~i23),
  i406 = \IN-i406 ,
  v8902 = (v8777 & i12) | (v8903 & ~i12),
  i407 = \IN-i407 ,
  v8903 = (v8777 & i13) | (v8904 & ~i13),
  i408 = \IN-i408 ,
  v8904 = (v8905 & i14) | (v8777 & ~i14),
  i409 = \IN-i409 ,
  v8905 = (v8907 & i21) | (v8906 & ~i21),
  v8906 = (v8628 & i23) | (v7791 & ~i23),
  v640 = (v617 & i30) | (v641 & ~i30),
  v8907 = (v8908 & i22) | (v8906 & ~i22),
  v641 = (v617 & i31) | (v642 & ~i31),
  v8908 = (v8632 & i23) | (v7794 & ~i23),
  v642 = (v617 & i32) | (v643 & ~i32),
  v8909 = (v10055 & i2) | (v8910 & ~i2),
  v643 = (~v644 & ~i34) | i34,
  v644 = (v653 & i36) | (v645 & ~i36),
  i410 = \IN-i410 ,
  v645 = (v652 & i37) | (v646 & ~i37),
  i411 = \IN-i411 ,
  v646 = (v648 & i38) | (v647 & ~i38),
  i412 = \IN-i412 ,
  v647 = (v648 & i39) | (v633 & ~i39),
  i413 = \IN-i413 ,
  v648 = (v649 & ~i41) | i41,
  i414 = \IN-i414 ,
  v649 = (v650 & ~i42) | i42,
  v8910 = (v10055 & i3) | (~v8911 & ~i3),
  i415 = \IN-i415 ,
  v8911 = (v9968 & i7) | (v8912 & ~i7),
  i416 = \IN-i416 ,
  v8912 = (v9968 & i8) | (v8913 & ~i8),
  v8913 = (v9968 & i9) | (v8914 & ~i9),
  v8914 = (v9885 & i10) | (v8915 & ~i10),
  v8915 = (v8919 & i11) | (v8916 & ~i11),
  v8916 = (v8919 & i12) | (v8917 & ~i12),
  v650 = (v651 & ~i43) | i43,
  v8917 = (v8919 & i13) | (v8918 & ~i13),
  v651 = (v632 & ~i44) | i44,
  v8918 = (v9885 & i14) | (v8919 & ~i14),
  v652 = (v648 & i38) | ~i38,
  v8919 = (v9516 & i15) | (v8920 & ~i15),
  v653 = (v652 & i37) | (v648 & ~i37),
  v654 = (v676 & i20) | (v655 & ~i20),
  v655 = (v656 & i21) | (v617 & ~i21),
  v656 = (v657 & i22) | (v617 & ~i22),
  v657 = (v658 & i25) | (v617 & ~i25),
  v658 = (v617 & i30) | (v659 & ~i30),
  v659 = (v617 & i31) | (v660 & ~i31),
  v8920 = (v9237 & i16) | (v8921 & ~i16),
  v8921 = (v9116 & i17) | (v8922 & ~i17),
  v8922 = (v9018 & i19) | (v8923 & ~i19),
  v8923 = (v8973 & i20) | (v8924 & ~i20),
  v8924 = (v8942 & i21) | (v8925 & ~i21),
  v8925 = (v8926 & i22) | ~i22,
  v8926 = (v8927 & i29) | ~i29,
  v660 = (v617 & i32) | (v661 & ~i32),
  v8927 = (v8928 & ~i30) | i30,
  v661 = (~v662 & ~i34) | i34,
  v8928 = (v8929 & i31) | ~i31,
  v662 = (v672 & i35) | (v663 & ~i35),
  v8929 = (v8930 & ~i32) | i32,
  v663 = (v671 & i36) | (v664 & ~i36),
  v664 = (v670 & i37) | (v665 & ~i37),
  v665 = (v666 & i38) | (v633 & ~i38),
  v666 = (v628 & i40) | (v667 & ~i40),
  v667 = (v668 & ~i41) | i41,
  v668 = (v669 & ~i42) | i42,
  v669 = (v632 & ~i43) | i43,
  v8930 = (v8941 & i36) | (v8931 & ~i36),
  v8931 = (v8940 & i37) | (v8932 & ~i37),
  v8932 = (v8934 & i38) | (v8933 & ~i38),
  v8933 = (v8938 & i39) | (v8934 & ~i39),
  v8934 = (v8935 & ~i41) | i41,
  v8935 = (v8936 & ~i42) | i42,
  v8936 = (v8937 & ~i43) | i43,
  v670 = (v666 & i38) | ~i38,
  v8937 = (v20 & i44) | ~i44,
  v671 = (v670 & i37) | (v666 & ~i37),
  v8938 = (v8939 & i42) | (v20 & ~i42),
  v672 = (v671 & i36) | (v673 & ~i36),
  v8939 = (v20 & i43) | ~i43,
  v673 = (v670 & i37) | (v674 & ~i37),
  v674 = (v666 & i38) | (v675 & ~i38),
  v675 = (v633 & i39) | (v666 & ~i39),
  v676 = (v677 & i21) | (v617 & ~i21),
  v677 = (v678 & i22) | (v617 & ~i22),
  v678 = (v679 & i25) | (v617 & ~i25),
  v679 = (v617 & i30) | (v680 & ~i30),
  v8940 = (v8934 & i38) | ~i38,
  v8941 = (v8940 & i37) | (v8934 & ~i37),
  v8942 = (v8959 & i22) | (v8943 & ~i22),
  v8943 = (v8944 & i29) | ~i29,
  v8944 = (v8945 & ~i30) | i30,
  v8945 = (v8946 & i31) | ~i31,
  v8946 = (v8947 & i32) | ~i32,
  v680 = (v617 & i31) | (v681 & ~i31),
  v8947 = (v8958 & i36) | (v8948 & ~i36),
  v681 = (v617 & i32) | (v682 & ~i32),
  v8948 = (v8957 & i37) | (v8949 & ~i37),
  v682 = (~v683 & ~i34) | i34,
  v8949 = (v8951 & i38) | (v8950 & ~i38),
  v683 = (v690 & i35) | (v684 & ~i35),
  v684 = (v689 & i36) | (v685 & ~i36),
  v685 = (v688 & i37) | (v686 & ~i37),
  v686 = (v687 & i38) | (v633 & ~i38),
  v687 = (v648 & i40) | (v667 & ~i40),
  v688 = (v687 & i38) | ~i38,
  v689 = (v688 & i37) | (v687 & ~i37),
  v8950 = (v8955 & i39) | (v8951 & ~i39),
  v8951 = (v8952 & ~i41) | i41,
  v8952 = (v8953 & ~i42) | i42,
  v8953 = (v8954 & ~i43) | i43,
  v8954 = (v49 & i44) | ~i44,
  v8955 = (v8956 & i42) | (v49 & ~i42),
  v8956 = (v49 & i43) | ~i43,
  v690 = (v689 & i36) | (v691 & ~i36),
  v8957 = (v8951 & i38) | ~i38,
  v691 = (v688 & i37) | (v692 & ~i37),
  v8958 = (v8957 & i37) | (v8951 & ~i37),
  v692 = (v687 & i38) | (v693 & ~i38),
  v8959 = (v8969 & i25) | (v8960 & ~i25),
  v693 = (v687 & i39) | (v633 & ~i39),
  v694 = (v732 & i19) | (v695 & ~i19),
  v695 = (v714 & i20) | (v696 & ~i20),
  v696 = (v697 & i21) | (v617 & ~i21),
  v697 = (v698 & i22) | (v617 & ~i22),
  v698 = (v699 & i25) | (v617 & ~i25),
  v699 = (v617 & i30) | (v700 & ~i30),
  v8960 = (v8961 & i29) | ~i29,
  v8961 = (v8964 & i30) | (v8962 & ~i30),
  v8962 = (v8963 & i31) | (v624 & ~i31),
  v8963 = (v8947 & i32) | (v8930 & ~i32),
  v8964 = (v8965 & i32) | (v628 & ~i32),
  v8965 = (v8966 & ~i36) | i36,
  v8966 = (v8967 & ~i37) | i37,
  v8967 = (v8968 & ~i38) | i38,
  v8968 = (v632 & i39) | ~i39,
  v8969 = (v8961 & i29) | (v8970 & ~i29),
  v8970 = (v8971 & ~i30) | i30,
  v8971 = (v8972 & ~i31) | i31,
  v8972 = (v624 & ~i32) | i32,
  v8973 = (v8989 & i21) | (v8974 & ~i21),
  v8974 = (v8975 & i22) | ~i22,
  v8975 = (v8976 & i29) | ~i29,
  v8976 = (v8977 & ~i30) | i30,
  v8977 = (v8978 & i31) | ~i31,
  v8978 = (v8979 & ~i32) | i32,
  v8979 = (v8988 & i36) | (v8980 & ~i36),
  v8980 = (v8987 & i37) | (v8981 & ~i37),
  v8981 = (v8983 & i38) | (v8982 & ~i38),
  v8982 = (v8983 & i39) | (v8938 & ~i39),
  v8983 = (v8984 & ~i41) | i41,
  v8984 = (v8985 & ~i42) | i42,
  v8985 = (v8986 & ~i43) | i43,
  v8986 = (v20 & ~i44) | i44,
  v8987 = (v8983 & i38) | ~i38,
  v8988 = (v8987 & i37) | (v8983 & ~i37),
  v8989 = (v9004 & i22) | (v8990 & ~i22),
  v8990 = (v8991 & i29) | ~i29,
  v8991 = (v8992 & ~i30) | i30,
  v8992 = (v8993 & i31) | ~i31,
  v8993 = (v8994 & i32) | ~i32,
  v8994 = (v9003 & i36) | (v8995 & ~i36),
  v8995 = (v9002 & i37) | (v8996 & ~i37),
  v8996 = (v8998 & i38) | (v8997 & ~i38),
  v8997 = (v8998 & i39) | (v8955 & ~i39),
  v8998 = (v8999 & ~i41) | i41,
  v8999 = (v9000 & ~i42) | i42,
  v700 = (v617 & i31) | (v701 & ~i31),
  v701 = (v617 & i32) | (v702 & ~i32),
  v702 = (~v703 & ~i34) | i34,
  v703 = (v711 & i35) | (v704 & ~i35),
  v704 = (v710 & i36) | (v705 & ~i36),
  v705 = (v709 & i37) | (v706 & ~i37),
  v706 = (v708 & i38) | (v707 & ~i38),
  v707 = (v633 & i39) | (v708 & ~i39),
  v708 = (v667 & i40) | (v628 & ~i40),
  v709 = (v708 & i38) | ~i38,
  v710 = (v709 & i37) | (v708 & ~i37),
  v711 = (v710 & i36) | (v712 & ~i36),
  v712 = (v709 & i37) | (v713 & ~i37),
  v713 = (v708 & i38) | (v633 & ~i38),
  v714 = (v715 & i21) | (v617 & ~i21),
  v715 = (v716 & i22) | (v617 & ~i22),
  v716 = (v717 & i25) | (v617 & ~i25),
  v717 = (v617 & i30) | (v718 & ~i30),
  v718 = (v617 & i31) | (v719 & ~i31),
  v719 = (v617 & i32) | (v720 & ~i32),
  v720 = (~v721 & ~i34) | i34,
  v721 = (v729 & i35) | (v722 & ~i35),
  v722 = (v728 & i36) | (v723 & ~i36),
  v723 = (v727 & i37) | (v724 & ~i37),
  v724 = (v726 & i38) | (v725 & ~i38),
  v725 = (v726 & i39) | (v633 & ~i39),
  v726 = (v667 & i40) | (v648 & ~i40),
  v727 = (v726 & i38) | ~i38,
  v728 = (v727 & i37) | (v726 & ~i37),
  v729 = (v728 & i36) | (v730 & ~i36),
  v730 = (v727 & i37) | (v731 & ~i37),
  v731 = (v726 & i38) | (v633 & ~i38),
  v732 = (v733 & i21) | (v617 & ~i21),
  v733 = (v734 & i22) | (v617 & ~i22),
  v734 = (v735 & i25) | (v617 & ~i25),
  v735 = (v617 & i30) | (v736 & ~i30),
  v736 = (v617 & i31) | (v737 & ~i31),
  v737 = (v617 & i32) | (v738 & ~i32),
  v738 = (~v739 & ~i34) | i34,
  v739 = (v743 & i36) | (v740 & ~i36),
  v740 = (v742 & i37) | (v741 & ~i37),
  v741 = (v667 & i38) | (v633 & ~i38),
  v742 = (v667 & i38) | ~i38,
  v743 = (v742 & i37) | (v667 & ~i37),
  v744 = (v812 & i17) | (v745 & ~i17),
  v745 = (v775 & i19) | (v746 & ~i19),
  v746 = (v761 & i20) | (v747 & ~i20),
  v747 = (v748 & i21) | (v617 & ~i21),
  v748 = (v749 & i22) | (v617 & ~i22),
  v749 = (v750 & i25) | (v617 & ~i25),
  v750 = (v617 & i30) | (v751 & ~i30),
  v751 = (v617 & i31) | (v752 & ~i31),
  v752 = (v617 & i32) | (v753 & ~i32),
  v753 = (~v754 & ~i34) | i34,
  v754 = (v760 & i36) | (v755 & ~i36),
  v755 = (v759 & i37) | (v756 & ~i37),
  v756 = (v758 & i38) | (v757 & ~i38),
  v757 = (v633 & i39) | (v758 & ~i39),
  v758 = (v668 & i41) | (v629 & ~i41),
  v759 = (v758 & i38) | ~i38,
  v760 = (v759 & i37) | (v758 & ~i37),
  v761 = (v762 & i21) | (v617 & ~i21),
  v762 = (v763 & i22) | (v617 & ~i22),
  v763 = (v764 & i25) | (v617 & ~i25),
  v764 = (v617 & i30) | (v765 & ~i30),
  v765 = (v617 & i31) | (v766 & ~i31),
  v766 = (v617 & i32) | (v767 & ~i32),
  v767 = (~v768 & ~i34) | i34,
  v768 = (v774 & i36) | (v769 & ~i36),
  v769 = (v773 & i37) | (v770 & ~i37),
  v770 = (v772 & i38) | (v771 & ~i38),
  v771 = (v772 & i39) | (v633 & ~i39),
  v772 = (v668 & i41) | (v649 & ~i41),
  v773 = (v772 & i38) | ~i38,
  v774 = (v773 & i37) | (v772 & ~i37),
  v775 = (v794 & i20) | (v776 & ~i20),
  v776 = (v777 & i21) | (v617 & ~i21),
  v777 = (v778 & i22) | (v617 & ~i22),
  v778 = (v779 & i25) | (v617 & ~i25),
  v779 = (v617 & i30) | (v780 & ~i30),
  v780 = (v617 & i31) | (v781 & ~i31),
  v781 = (v617 & i32) | (v782 & ~i32),
  v782 = (~v783 & ~i34) | i34,
  v783 = (v790 & i35) | (v784 & ~i35),
  v784 = (v789 & i36) | (v785 & ~i36),
  v785 = (v788 & i37) | (v786 & ~i37),
  v786 = (v787 & i38) | (v633 & ~i38),
  v787 = (v758 & i40) | (v668 & ~i40),
  v788 = (v787 & i38) | ~i38,
  v789 = (v788 & i37) | (v787 & ~i37),
  v790 = (v789 & i36) | (v791 & ~i36),
  v791 = (v788 & i37) | (v792 & ~i37),
  v792 = (v787 & i38) | (v793 & ~i38),
  v793 = (v633 & i39) | (v787 & ~i39),
  v794 = (v795 & i21) | (v617 & ~i21),
  v795 = (v796 & i22) | (v617 & ~i22),
  v796 = (v797 & i25) | (v617 & ~i25),
  v797 = (v617 & i30) | (v798 & ~i30),
  v798 = (v617 & i31) | (v799 & ~i31),
  v799 = (v617 & i32) | (v800 & ~i32),
  v800 = (~v801 & ~i34) | i34,
  v801 = (v808 & i35) | (v802 & ~i35),
  v802 = (v807 & i36) | (v803 & ~i36),
  v803 = (v806 & i37) | (v804 & ~i37),
  v804 = (v805 & i38) | (v633 & ~i38),
  v805 = (v772 & i40) | (v668 & ~i40),
  v806 = (v805 & i38) | ~i38,
  v807 = (v806 & i37) | (v805 & ~i37),
  v808 = (v807 & i36) | (v809 & ~i36),
  v809 = (v806 & i37) | (v810 & ~i37),
  v810 = (v805 & i38) | (v811 & ~i38),
  v811 = (v805 & i39) | (v633 & ~i39),
  v812 = (v850 & i19) | (v813 & ~i19),
  v813 = (v832 & i20) | (v814 & ~i20),
  v814 = (v815 & i21) | (v617 & ~i21),
  v815 = (v816 & i22) | (v617 & ~i22),
  v816 = (v817 & i25) | (v617 & ~i25),
  v817 = (v617 & i30) | (v818 & ~i30),
  v818 = (v617 & i31) | (v819 & ~i31),
  v819 = (v617 & i32) | (v820 & ~i32),
  v820 = (~v821 & ~i34) | i34,
  v821 = (v829 & i35) | (v822 & ~i35),
  v822 = (v828 & i36) | (v823 & ~i36),
  v823 = (v827 & i37) | (v824 & ~i37),
  v824 = (v826 & i38) | (v825 & ~i38),
  v825 = (v633 & i39) | (v826 & ~i39),
  v826 = (v668 & i40) | (v758 & ~i40),
  v827 = (v826 & i38) | ~i38,
  v828 = (v827 & i37) | (v826 & ~i37),
  v829 = (v828 & i36) | (v830 & ~i36),
  v830 = (v827 & i37) | (v831 & ~i37),
  v831 = (v826 & i38) | (v633 & ~i38),
  v832 = (v833 & i21) | (v617 & ~i21),
  v833 = (v834 & i22) | (v617 & ~i22),
  v834 = (v835 & i25) | (v617 & ~i25),
  v835 = (v617 & i30) | (v836 & ~i30),
  v836 = (v617 & i31) | (v837 & ~i31),
  v837 = (v617 & i32) | (v838 & ~i32),
  v838 = (~v839 & ~i34) | i34,
  v839 = (v847 & i35) | (v840 & ~i35),
  v840 = (v846 & i36) | (v841 & ~i36),
  v841 = (v845 & i37) | (v842 & ~i37),
  v842 = (v844 & i38) | (v843 & ~i38),
  v843 = (v844 & i39) | (v633 & ~i39),
  v844 = (v668 & i40) | (v772 & ~i40),
  v845 = (v844 & i38) | ~i38,
  v846 = (v845 & i37) | (v844 & ~i37),
  v847 = (v846 & i36) | (v848 & ~i36),
  v848 = (v845 & i37) | (v849 & ~i37),
  v849 = (v844 & i38) | (v633 & ~i38),
  v850 = (v851 & i21) | (v617 & ~i21),
  v851 = (v852 & i22) | (v617 & ~i22),
  v852 = (v853 & i25) | (v617 & ~i25),
  v853 = (v617 & i30) | (v854 & ~i30),
  v854 = (v617 & i31) | (v855 & ~i31),
  v855 = (v617 & i32) | (v856 & ~i32),
  v856 = (~v857 & ~i34) | i34,
  v857 = (v861 & i36) | (v858 & ~i36),
  v858 = (v860 & i37) | (v859 & ~i37),
  v859 = (v668 & i38) | (v633 & ~i38),
  v860 = (v668 & i38) | ~i38,
  v861 = (v860 & i37) | (v668 & ~i37),
  v862 = (v932 & i16) | (v863 & ~i16),
  v863 = (v905 & i17) | (v864 & ~i17),
  v864 = (v886 & i19) | (v865 & ~i19),
  v865 = (v876 & i20) | (v866 & ~i20),
  v866 = (v867 & i21) | (v617 & ~i21),
  v867 = (v868 & i22) | (v617 & ~i22),
  v868 = (v869 & i25) | (v617 & ~i25),
  v869 = (v617 & i30) | (v870 & ~i30),
  v870 = (v617 & i31) | (v871 & ~i31),
  v871 = (v617 & i32) | (v872 & ~i32),
  v872 = (~v873 & ~i34) | i34,
  v873 = (v874 & i36) | (v625 & ~i36),
  v874 = (v635 & i37) | (v875 & ~i37),
  v875 = (v628 & i38) | (v633 & ~i38),
  v876 = (v877 & i21) | (v617 & ~i21),
  v877 = (v878 & i22) | (v617 & ~i22),
  v878 = (v879 & i25) | (v617 & ~i25),
  v879 = (v617 & i30) | (v880 & ~i30),
  v880 = (v617 & i31) | (v881 & ~i31),
  v881 = (v617 & i32) | (v882 & ~i32),
  v882 = (~v883 & ~i34) | i34,
  v883 = (v884 & i36) | (v645 & ~i36),
  v884 = (v652 & i37) | (v885 & ~i37),
  v885 = (v648 & i38) | (v633 & ~i38),
  v886 = (v896 & i20) | (v887 & ~i20),
  v887 = (v888 & i21) | (v617 & ~i21),
  v888 = (v889 & i22) | (v617 & ~i22),
  v889 = (v890 & i25) | (v617 & ~i25),
  v890 = (v617 & i30) | (v891 & ~i30),
  v891 = (v617 & i31) | (v892 & ~i31),
  v892 = (v617 & i32) | (v893 & ~i32),
  v893 = (~v894 & ~i34) | i34,
  v894 = (v895 & i35) | (v664 & ~i35),
  v895 = (v664 & i36) | (v673 & ~i36),
  v896 = (v897 & i21) | (v617 & ~i21),
  v897 = (v898 & i22) | (v617 & ~i22),
  v898 = (v899 & i25) | (v617 & ~i25),
  v899 = (v617 & i30) | (v900 & ~i30),
  v900 = (v617 & i31) | (v901 & ~i31),
  v901 = (v617 & i32) | (v902 & ~i32),
  v902 = (~v903 & ~i34) | i34,
  v903 = (v904 & i35) | (v685 & ~i35),
  v904 = (v685 & i36) | (v691 & ~i36),
  v905 = (v925 & i19) | (v906 & ~i19),
  v906 = (v916 & i20) | (v907 & ~i20),
  v907 = (v908 & i21) | (v617 & ~i21),
  v908 = (v909 & i22) | (v617 & ~i22),
  v909 = (v910 & i25) | (v617 & ~i25),
  v910 = (v617 & i30) | (v911 & ~i30),
  v911 = (v617 & i31) | (v912 & ~i31),
  v912 = (v617 & i32) | (v913 & ~i32),
  v913 = (~v914 & ~i34) | i34,
  v914 = (v712 & i35) | (v915 & ~i35),
  v915 = (v712 & i36) | (v705 & ~i36),
  v916 = (v917 & i21) | (v617 & ~i21),
  v917 = (v918 & i22) | (v617 & ~i22),
  v918 = (v919 & i25) | (v617 & ~i25),
  v919 = (v617 & i30) | (v920 & ~i30),
  v920 = (v617 & i31) | (v921 & ~i31),
  v921 = (v617 & i32) | (v922 & ~i32),
  v922 = (~v923 & ~i34) | i34,
  v923 = (v730 & i35) | (v924 & ~i35),
  v924 = (v730 & i36) | (v723 & ~i36),
  v925 = (v926 & i21) | (v617 & ~i21),
  v926 = (v927 & i22) | (v617 & ~i22),
  v927 = (v928 & i25) | (v617 & ~i25),
  v928 = (v617 & i30) | (v929 & ~i30),
  v929 = (v617 & i31) | (v930 & ~i31),
  v930 = (v617 & i32) | (v931 & ~i32),
  v931 = (~v740 & ~i34) | i34,
  v932 = (v974 & i17) | (v933 & ~i17),
  v933 = (v955 & i19) | (v934 & ~i19),
  v934 = (v945 & i20) | (v935 & ~i20),
  v935 = (v936 & i21) | (v617 & ~i21),
  v936 = (v937 & i22) | (v617 & ~i22),
  v937 = (v938 & i25) | (v617 & ~i25),
  v938 = (v617 & i30) | (v939 & ~i30),
  v939 = (v617 & i31) | (v940 & ~i31),
  v940 = (v617 & i32) | (v941 & ~i32),
  v941 = (~v942 & ~i34) | i34,
  v942 = (v943 & i36) | (v755 & ~i36),
  v943 = (v759 & i37) | (v944 & ~i37),
  v944 = (v758 & i38) | (v633 & ~i38),
  v945 = (v946 & i21) | (v617 & ~i21),
  v946 = (v947 & i22) | (v617 & ~i22),
  v947 = (v948 & i25) | (v617 & ~i25),
  v948 = (v617 & i30) | (v949 & ~i30),
  v949 = (v617 & i31) | (v950 & ~i31),
  v950 = (v617 & i32) | (v951 & ~i32),
  v951 = (~v952 & ~i34) | i34,
  v952 = (v953 & i36) | (v769 & ~i36),
  v953 = (v773 & i37) | (v954 & ~i37),
  v954 = (v772 & i38) | (v633 & ~i38),
  v955 = (v965 & i20) | (v956 & ~i20),
  v956 = (v957 & i21) | (v617 & ~i21),
  v957 = (v958 & i22) | (v617 & ~i22),
  v958 = (v959 & i25) | (v617 & ~i25),
  v959 = (v617 & i30) | (v960 & ~i30),
  v960 = (v617 & i31) | (v961 & ~i31),
  v961 = (v617 & i32) | (v962 & ~i32),
  v962 = (~v963 & ~i34) | i34,
  v963 = (v964 & i35) | (v785 & ~i35),
  v964 = (v785 & i36) | (v791 & ~i36),
  v965 = (v966 & i21) | (v617 & ~i21),
  v966 = (v967 & i22) | (v617 & ~i22),
  v967 = (v968 & i25) | (v617 & ~i25),
  v968 = (v617 & i30) | (v969 & ~i30),
  v969 = (v617 & i31) | (v970 & ~i31),
  v970 = (v617 & i32) | (v971 & ~i32),
  v971 = (~v972 & ~i34) | i34,
  v972 = (v973 & i35) | (v803 & ~i35),
  v973 = (v803 & i36) | (v809 & ~i36),
  v974 = (v994 & i19) | (v975 & ~i19),
  v975 = (v985 & i20) | (v976 & ~i20),
  v976 = (v977 & i21) | (v617 & ~i21),
  v977 = (v978 & i22) | (v617 & ~i22),
  v978 = (v979 & i25) | (v617 & ~i25),
  v979 = (v617 & i30) | (v980 & ~i30),
  v980 = (v617 & i31) | (v981 & ~i31),
  v981 = (v617 & i32) | (v982 & ~i32),
  v982 = (~v983 & ~i34) | i34,
  v983 = (v830 & i35) | (v984 & ~i35),
  v984 = (v830 & i36) | (v823 & ~i36),
  v985 = (v986 & i21) | (v617 & ~i21),
  v986 = (v987 & i22) | (v617 & ~i22),
  v987 = (v988 & i25) | (v617 & ~i25),
  v988 = (v617 & i30) | (v989 & ~i30),
  v989 = (v617 & i31) | (v990 & ~i31),
  v990 = (v617 & i32) | (v991 & ~i32),
  v991 = (~v992 & ~i34) | i34,
  v992 = (v848 & i35) | (v993 & ~i35),
  v993 = (v848 & i36) | (v841 & ~i36),
  v994 = (v995 & i21) | (v617 & ~i21),
  v995 = (v996 & i22) | (v617 & ~i22),
  v996 = (v997 & i25) | (v617 & ~i25),
  v997 = (v617 & i30) | (v998 & ~i30),
  v998 = (v617 & i31) | (v999 & ~i31),
  v999 = (v617 & i32) | (v1000 & ~i32),
  v9000 = (v9001 & ~i43) | i43,
  v9001 = (v49 & ~i44) | i44,
  v9002 = (v8998 & i38) | ~i38,
  v9003 = (v9002 & i37) | (v8998 & ~i37),
  v9004 = (v9014 & i25) | (v9005 & ~i25),
  v9005 = (v9006 & i29) | ~i29,
  v9006 = (v9009 & i30) | (v9007 & ~i30),
  v9007 = (v9008 & i31) | (v644 & ~i31),
  v9008 = (v8994 & i32) | (v8979 & ~i32),
  v9009 = (v9010 & i32) | (v648 & ~i32),
  v9010 = (v9011 & ~i36) | i36,
  v9011 = (v9012 & ~i37) | i37,
  v9012 = (v9013 & ~i38) | i38,
  v9013 = (v632 & ~i39) | i39,
  v9014 = (v9006 & i29) | (v9015 & ~i29),
  v9015 = (v9016 & ~i30) | i30,
  v9016 = (v9017 & ~i31) | i31,
  v9017 = (v644 & ~i32) | i32,
  v9018 = (v9072 & i20) | (v9019 & ~i20),
  v9019 = (v9039 & i21) | (v9020 & ~i21),
  v9020 = (v9021 & i22) | ~i22,
  v9021 = (v9022 & i29) | ~i29,
  v9022 = (v9023 & ~i30) | i30,
  v9023 = (v9024 & i31) | ~i31,
  v9024 = (v9025 & ~i32) | i32,
  v9025 = (v9035 & i35) | (v9026 & ~i35),
  v9026 = (v9034 & i36) | (v9027 & ~i36),
  v9027 = (v9033 & i37) | (v9028 & ~i37),
  v9028 = (v9029 & i38) | (v8938 & ~i38),
  v9029 = (v8934 & i40) | (v9030 & ~i40),
  v9030 = (v9031 & ~i41) | i41,
  v9031 = (v9032 & ~i42) | i42,
  v9032 = (v20 & ~i43) | i43,
  v9033 = (v9029 & i38) | ~i38,
  v9034 = (v9033 & i37) | (v9029 & ~i37),
  v9035 = (v9034 & i36) | (v9036 & ~i36),
  v9036 = (v9033 & i37) | (v9037 & ~i37),
  v9037 = (v9029 & i38) | (v9038 & ~i38),
  v9038 = (v8938 & i39) | (v9029 & ~i39),
  v9039 = (v9058 & i22) | (v9040 & ~i22),
  v9040 = (v9041 & i29) | ~i29,
  v9041 = (v9042 & ~i30) | i30,
  v9042 = (v9043 & i31) | ~i31,
  v9043 = (v9044 & i32) | ~i32,
  v9044 = (v9054 & i35) | (v9045 & ~i35),
  v9045 = (v9053 & i36) | (v9046 & ~i36),
  v9046 = (v9052 & i37) | (v9047 & ~i37),
  v9047 = (v9048 & i38) | (v8955 & ~i38),
  v9048 = (v8951 & i40) | (v9049 & ~i40),
  v9049 = (v9050 & ~i41) | i41,
  v9050 = (v9051 & ~i42) | i42,
  v9051 = (v49 & ~i43) | i43,
  v9052 = (v9048 & i38) | ~i38,
  v9053 = (v9052 & i37) | (v9048 & ~i37),
  v9054 = (v9053 & i36) | (v9055 & ~i36),
  v9055 = (v9052 & i37) | (v9056 & ~i37),
  v9056 = (v9048 & i38) | (v9057 & ~i38),
  v9057 = (v8955 & i39) | (v9048 & ~i39),
  v9058 = (v9068 & i25) | (v9059 & ~i25),
  v9059 = (v9060 & i29) | ~i29,
  v9060 = (v9063 & i30) | (v9061 & ~i30),
  v9061 = (v9062 & i31) | (v662 & ~i31),
  v9062 = (v9044 & i32) | (v9025 & ~i32),
  v9063 = (v9064 & i32) | (v666 & ~i32),
  v9064 = (v8965 & i35) | (v9065 & ~i35),
  v9065 = (v9066 & ~i36) | i36,
  v9066 = (v9067 & ~i37) | i37,
  v9067 = (v632 & ~i38) | i38,
  v9068 = (v9060 & i29) | (v9069 & ~i29),
  v9069 = (v9070 & ~i30) | i30,
  v9070 = (v9071 & ~i31) | i31,
  v9071 = (v662 & ~i32) | i32,
  v9072 = (v9089 & i21) | (v9073 & ~i21),
  v9073 = (v9074 & i22) | ~i22,
  v9074 = (v9075 & i29) | ~i29,
  v9075 = (v9076 & ~i30) | i30,
  v9076 = (v9077 & i31) | ~i31,
  v9077 = (v9078 & ~i32) | i32,
  v9078 = (v9085 & i35) | (v9079 & ~i35),
  v9079 = (v9084 & i36) | (v9080 & ~i36),
  v9080 = (v9083 & i37) | (v9081 & ~i37),
  v9081 = (v9082 & i38) | (v8938 & ~i38),
  v9082 = (v8983 & i40) | (v9030 & ~i40),
  v9083 = (v9082 & i38) | ~i38,
  v9084 = (v9083 & i37) | (v9082 & ~i37),
  v9085 = (v9084 & i36) | (v9086 & ~i36),
  v9086 = (v9083 & i37) | (v9087 & ~i37),
  v9087 = (v9082 & i38) | (v9088 & ~i38),
  v9088 = (v9082 & i39) | (v8938 & ~i39),
  v9089 = (v9105 & i22) | (v9090 & ~i22),
  v9090 = (v9091 & i29) | ~i29,
  v9091 = (v9092 & ~i30) | i30,
  v9092 = (v9093 & i31) | ~i31,
  v9093 = (v9094 & i32) | ~i32,
  v9094 = (v9101 & i35) | (v9095 & ~i35),
  v9095 = (v9100 & i36) | (v9096 & ~i36),
  v9096 = (v9099 & i37) | (v9097 & ~i37),
  v9097 = (v9098 & i38) | (v8955 & ~i38),
  v9098 = (v8998 & i40) | (v9049 & ~i40),
  v9099 = (v9098 & i38) | ~i38,
  v9100 = (v9099 & i37) | (v9098 & ~i37),
  v9101 = (v9100 & i36) | (v9102 & ~i36),
  v9102 = (v9099 & i37) | (v9103 & ~i37),
  v9103 = (v9098 & i38) | (v9104 & ~i38),
  v9104 = (v9098 & i39) | (v8955 & ~i39),
  v9105 = (v9112 & i25) | (v9106 & ~i25),
  v9106 = (v9107 & i29) | ~i29,
  v9107 = (v9110 & i30) | (v9108 & ~i30),
  v9108 = (v9109 & i31) | (v683 & ~i31),
  v9109 = (v9094 & i32) | (v9078 & ~i32),
  v9110 = (v9111 & i32) | (v687 & ~i32),
  v9111 = (v9010 & i35) | (v9065 & ~i35),
  v9112 = (v9107 & i29) | (v9113 & ~i29),
  v9113 = (v9114 & ~i30) | i30,
  v9114 = (v9115 & ~i31) | i31,
  v9115 = (v683 & ~i32) | i32,
  v9116 = (v9206 & i19) | (v9117 & ~i19),
  v9117 = (v9162 & i20) | (v9118 & ~i20),
  v9118 = (v9135 & i21) | (v9119 & ~i21),
  v9119 = (v9120 & i22) | ~i22,
  v9120 = (v9121 & i29) | ~i29,
  v9121 = (v9122 & ~i30) | i30,
  v9122 = (v9123 & i31) | ~i31,
  v9123 = (v9124 & ~i32) | i32,
  v9124 = (v9132 & i35) | (v9125 & ~i35),
  v9125 = (v9131 & i36) | (v9126 & ~i36),
  v9126 = (v9130 & i37) | (v9127 & ~i37),
  v9127 = (v9129 & i38) | (v9128 & ~i38),
  v9128 = (v8938 & i39) | (v9129 & ~i39),
  v9129 = (v9030 & i40) | (v8934 & ~i40),
  v9130 = (v9129 & i38) | ~i38,
  v9131 = (v9130 & i37) | (v9129 & ~i37),
  v9132 = (v9131 & i36) | (v9133 & ~i36),
  v9133 = (v9130 & i37) | (v9134 & ~i37),
  v9134 = (v9129 & i38) | (v8938 & ~i38),
  v9135 = (v9151 & i22) | (v9136 & ~i22),
  v9136 = (v9137 & i29) | ~i29,
  v9137 = (v9138 & ~i30) | i30,
  v9138 = (v9139 & i31) | ~i31,
  v9139 = (v9140 & i32) | ~i32,
  v9140 = (v9148 & i35) | (v9141 & ~i35),
  v9141 = (v9147 & i36) | (v9142 & ~i36),
  v9142 = (v9146 & i37) | (v9143 & ~i37),
  v9143 = (v9145 & i38) | (v9144 & ~i38),
  v9144 = (v8955 & i39) | (v9145 & ~i39),
  v9145 = (v9049 & i40) | (v8951 & ~i40),
  v9146 = (v9145 & i38) | ~i38,
  v9147 = (v9146 & i37) | (v9145 & ~i37),
  v9148 = (v9147 & i36) | (v9149 & ~i36),
  v9149 = (v9146 & i37) | (v9150 & ~i37),
  v9150 = (v9145 & i38) | (v8955 & ~i38),
  v9151 = (v9158 & i25) | (v9152 & ~i25),
  v9152 = (v9153 & i29) | ~i29,
  v9153 = (v9156 & i30) | (v9154 & ~i30),
  v9154 = (v9155 & i31) | (v703 & ~i31),
  v9155 = (v9140 & i32) | (v9124 & ~i32),
  v9156 = (v9157 & i32) | (v708 & ~i32),
  v9157 = (v9065 & i35) | (v8965 & ~i35),
  v9158 = (v9153 & i29) | (v9159 & ~i29),
  v9159 = (v9160 & ~i30) | i30,
  v9160 = (v9161 & ~i31) | i31,
  v9161 = (v703 & ~i32) | i32,
  v9162 = (v9179 & i21) | (v9163 & ~i21),
  v9163 = (v9164 & i22) | ~i22,
  v9164 = (v9165 & i29) | ~i29,
  v9165 = (v9166 & ~i30) | i30,
  v9166 = (v9167 & i31) | ~i31,
  v9167 = (v9168 & ~i32) | i32,
  v9168 = (v9176 & i35) | (v9169 & ~i35),
  v9169 = (v9175 & i36) | (v9170 & ~i36),
  v9170 = (v9174 & i37) | (v9171 & ~i37),
  v9171 = (v9173 & i38) | (v9172 & ~i38),
  v9172 = (v9173 & i39) | (v8938 & ~i39),
  v9173 = (v9030 & i40) | (v8983 & ~i40),
  v9174 = (v9173 & i38) | ~i38,
  v9175 = (v9174 & i37) | (v9173 & ~i37),
  v9176 = (v9175 & i36) | (v9177 & ~i36),
  v9177 = (v9174 & i37) | (v9178 & ~i37),
  v9178 = (v9173 & i38) | (v8938 & ~i38),
  v9179 = (v9195 & i22) | (v9180 & ~i22),
  v9180 = (v9181 & i29) | ~i29,
  v9181 = (v9182 & ~i30) | i30,
  v9182 = (v9183 & i31) | ~i31,
  v9183 = (v9184 & i32) | ~i32,
  v9184 = (v9192 & i35) | (v9185 & ~i35),
  v9185 = (v9191 & i36) | (v9186 & ~i36),
  v9186 = (v9190 & i37) | (v9187 & ~i37),
  v9187 = (v9189 & i38) | (v9188 & ~i38),
  v9188 = (v9189 & i39) | (v8955 & ~i39),
  v9189 = (v9049 & i40) | (v8998 & ~i40),
  v9190 = (v9189 & i38) | ~i38,
  v9191 = (v9190 & i37) | (v9189 & ~i37),
  v9192 = (v9191 & i36) | (v9193 & ~i36),
  v9193 = (v9190 & i37) | (v9194 & ~i37),
  v9194 = (v9189 & i38) | (v8955 & ~i38),
  v9195 = (v9202 & i25) | (v9196 & ~i25),
  v9196 = (v9197 & i29) | ~i29,
  v9197 = (v9200 & i30) | (v9198 & ~i30),
  v9198 = (v9199 & i31) | (v721 & ~i31),
  v9199 = (v9184 & i32) | (v9168 & ~i32),
  v9200 = (v9201 & i32) | (v726 & ~i32),
  v9201 = (v9065 & i35) | (v9010 & ~i35),
  v9202 = (v9197 & i29) | (v9203 & ~i29),
  v9203 = (v9204 & ~i30) | i30,
  v9204 = (v9205 & ~i31) | i31,
  v9205 = (v721 & ~i32) | i32,
  v9206 = (v9217 & i21) | (v9207 & ~i21),
  v9207 = (v9208 & i22) | ~i22,
  v9208 = (v9209 & i29) | ~i29,
  v9209 = (v9210 & ~i30) | i30,
  v9210 = (v9211 & i31) | ~i31,
  v9211 = (v9212 & ~i32) | i32,
  v9212 = (v9216 & i36) | (v9213 & ~i36),
  v9213 = (v9215 & i37) | (v9214 & ~i37),
  v9214 = (v9030 & i38) | (v8938 & ~i38),
  v9215 = (v9030 & i38) | ~i38,
  v9216 = (v9215 & i37) | (v9030 & ~i37),
  v9217 = (v9227 & i22) | (v9218 & ~i22),
  v9218 = (v9219 & i29) | ~i29,
  v9219 = (v9220 & ~i30) | i30,
  v9220 = (v9221 & i31) | ~i31,
  v9221 = (v9222 & i32) | ~i32,
  v9222 = (v9226 & i36) | (v9223 & ~i36),
  v9223 = (v9225 & i37) | (v9224 & ~i37),
  v9224 = (v9049 & i38) | (v8955 & ~i38),
  v9225 = (v9049 & i38) | ~i38,
  v9226 = (v9225 & i37) | (v9049 & ~i37),
  v9227 = (v9233 & i25) | (v9228 & ~i25),
  v9228 = (v9229 & i29) | ~i29,
  v9229 = (v9232 & i30) | (v9230 & ~i30),
  v9230 = (v9231 & i31) | (v739 & ~i31),
  v9231 = (v9222 & i32) | (v9212 & ~i32),
  v9232 = (v9065 & i32) | (v667 & ~i32),
  v9233 = (v9229 & i29) | (v9234 & ~i29),
  v9234 = (v9235 & ~i30) | i30,
  v9235 = (v9236 & ~i31) | i31,
  v9236 = (v739 & ~i32) | i32,
  v9237 = (v9397 & i17) | (v9238 & ~i17),
  v9238 = (v9310 & i19) | (v9239 & ~i19),
  v9239 = (v9275 & i20) | (v9240 & ~i20),
  v9240 = (v9253 & i21) | (v9241 & ~i21),
  v9241 = (v9242 & i22) | ~i22,
  v9242 = (v9243 & i29) | ~i29,
  v9243 = (v9244 & ~i30) | i30,
  v9244 = (v9245 & i31) | ~i31,
  v9245 = (v9246 & ~i32) | i32,
  v9246 = (v9252 & i36) | (v9247 & ~i36),
  v9247 = (v9251 & i37) | (v9248 & ~i37),
  v9248 = (v9250 & i38) | (v9249 & ~i38),
  v9249 = (v8938 & i39) | (v9250 & ~i39),
  v9250 = (v9031 & i41) | (v8935 & ~i41),
  v9251 = (v9250 & i38) | ~i38,
  v9252 = (v9251 & i37) | (v9250 & ~i37),
  v9253 = (v9265 & i22) | (v9254 & ~i22),
  v9254 = (v9255 & i29) | ~i29,
  v9255 = (v9256 & ~i30) | i30,
  v9256 = (v9257 & i31) | ~i31,
  v9257 = (v9258 & i32) | ~i32,
  v9258 = (v9264 & i36) | (v9259 & ~i36),
  v9259 = (v9263 & i37) | (v9260 & ~i37),
  v9260 = (v9262 & i38) | (v9261 & ~i38),
  v9261 = (v8955 & i39) | (v9262 & ~i39),
  v9262 = (v9050 & i41) | (v8952 & ~i41),
  v9263 = (v9262 & i38) | ~i38,
  v9264 = (v9263 & i37) | (v9262 & ~i37),
  v9265 = (v9271 & i25) | (v9266 & ~i25),
  v9266 = (v9267 & i29) | ~i29,
  v9267 = (v9270 & i30) | (v9268 & ~i30),
  v9268 = (v9269 & i31) | (v754 & ~i31),
  v9269 = (v9258 & i32) | (v9246 & ~i32),
  v9270 = (v8965 & i32) | (v758 & ~i32),
  v9271 = (v9267 & i29) | (v9272 & ~i29),
  v9272 = (v9273 & ~i30) | i30,
  v9273 = (v9274 & ~i31) | i31,
  v9274 = (v754 & ~i32) | i32,
  v9275 = (v9288 & i21) | (v9276 & ~i21),
  v9276 = (v9277 & i22) | ~i22,
  v9277 = (v9278 & i29) | ~i29,
  v9278 = (v9279 & ~i30) | i30,
  v9279 = (v9280 & i31) | ~i31,
  v9280 = (v9281 & ~i32) | i32,
  v9281 = (v9287 & i36) | (v9282 & ~i36),
  v9282 = (v9286 & i37) | (v9283 & ~i37),
  v9283 = (v9285 & i38) | (v9284 & ~i38),
  v9284 = (v9285 & i39) | (v8938 & ~i39),
  v9285 = (v9031 & i41) | (v8984 & ~i41),
  v9286 = (v9285 & i38) | ~i38,
  v9287 = (v9286 & i37) | (v9285 & ~i37),
  v9288 = (v9300 & i22) | (v9289 & ~i22),
  v9289 = (v9290 & i29) | ~i29,
  v9290 = (v9291 & ~i30) | i30,
  v9291 = (v9292 & i31) | ~i31,
  v9292 = (v9293 & i32) | ~i32,
  v9293 = (v9299 & i36) | (v9294 & ~i36),
  v9294 = (v9298 & i37) | (v9295 & ~i37),
  v9295 = (v9297 & i38) | (v9296 & ~i38),
  v9296 = (v9297 & i39) | (v8955 & ~i39),
  v9297 = (v9050 & i41) | (v8999 & ~i41),
  v9298 = (v9297 & i38) | ~i38,
  v9299 = (v9298 & i37) | (v9297 & ~i37),
  v9300 = (v9306 & i25) | (v9301 & ~i25),
  v9301 = (v9302 & i29) | ~i29,
  v9302 = (v9305 & i30) | (v9303 & ~i30),
  v9303 = (v9304 & i31) | (v768 & ~i31),
  v9304 = (v9293 & i32) | (v9281 & ~i32),
  v9305 = (v9010 & i32) | (v772 & ~i32),
  v9306 = (v9302 & i29) | (v9307 & ~i29),
  v9307 = (v9308 & ~i30) | i30,
  v9308 = (v9309 & ~i31) | i31,
  v9309 = (v768 & ~i32) | i32,
  v9310 = (v9354 & i20) | (v9311 & ~i20),
  v9311 = (v9328 & i21) | (v9312 & ~i21),
  v9312 = (v9313 & i22) | ~i22,
  v9313 = (v9314 & i29) | ~i29,
  v9314 = (v9315 & ~i30) | i30,
  v9315 = (v9316 & i31) | ~i31,
  v9316 = (v9317 & ~i32) | i32,
  v9317 = (v9324 & i35) | (v9318 & ~i35),
  v9318 = (v9323 & i36) | (v9319 & ~i36),
  v9319 = (v9322 & i37) | (v9320 & ~i37),
  v9320 = (v9321 & i38) | (v8938 & ~i38),
  v9321 = (v9250 & i40) | (v9031 & ~i40),
  v9322 = (v9321 & i38) | ~i38,
  v9323 = (v9322 & i37) | (v9321 & ~i37),
  v9324 = (v9323 & i36) | (v9325 & ~i36),
  v9325 = (v9322 & i37) | (v9326 & ~i37),
  v9326 = (v9321 & i38) | (v9327 & ~i38),
  v9327 = (v8938 & i39) | (v9321 & ~i39),
  v9328 = (v9344 & i22) | (v9329 & ~i22),
  v9329 = (v9330 & i29) | ~i29,
  v9330 = (v9331 & ~i30) | i30,
  v9331 = (v9332 & i31) | ~i31,
  v9332 = (v9333 & i32) | ~i32,
  v9333 = (v9340 & i35) | (v9334 & ~i35),
  v9334 = (v9339 & i36) | (v9335 & ~i36),
  v9335 = (v9338 & i37) | (v9336 & ~i37),
  v9336 = (v9337 & i38) | (v8955 & ~i38),
  v9337 = (v9262 & i40) | (v9050 & ~i40),
  v9338 = (v9337 & i38) | ~i38,
  v9339 = (v9338 & i37) | (v9337 & ~i37),
  v9340 = (v9339 & i36) | (v9341 & ~i36),
  v9341 = (v9338 & i37) | (v9342 & ~i37),
  v9342 = (v9337 & i38) | (v9343 & ~i38),
  v9343 = (v8955 & i39) | (v9337 & ~i39),
  v9344 = (v9350 & i25) | (v9345 & ~i25),
  v9345 = (v9346 & i29) | ~i29,
  v9346 = (v9349 & i30) | (v9347 & ~i30),
  v9347 = (v9348 & i31) | (v783 & ~i31),
  v9348 = (v9333 & i32) | (v9317 & ~i32),
  v9349 = (v9064 & i32) | (v787 & ~i32),
  v9350 = (v9346 & i29) | (v9351 & ~i29),
  v9351 = (v9352 & ~i30) | i30,
  v9352 = (v9353 & ~i31) | i31,
  v9353 = (v783 & ~i32) | i32,
  v9354 = (v9371 & i21) | (v9355 & ~i21),
  v9355 = (v9356 & i22) | ~i22,
  v9356 = (v9357 & i29) | ~i29,
  v9357 = (v9358 & ~i30) | i30,
  v9358 = (v9359 & i31) | ~i31,
  v9359 = (v9360 & ~i32) | i32,
  v9360 = (v9367 & i35) | (v9361 & ~i35),
  v9361 = (v9366 & i36) | (v9362 & ~i36),
  v9362 = (v9365 & i37) | (v9363 & ~i37),
  v9363 = (v9364 & i38) | (v8938 & ~i38),
  v9364 = (v9285 & i40) | (v9031 & ~i40),
  v9365 = (v9364 & i38) | ~i38,
  v9366 = (v9365 & i37) | (v9364 & ~i37),
  v9367 = (v9366 & i36) | (v9368 & ~i36),
  v9368 = (v9365 & i37) | (v9369 & ~i37),
  v9369 = (v9364 & i38) | (v9370 & ~i38),
  v9370 = (v9364 & i39) | (v8938 & ~i39),
  v9371 = (v9387 & i22) | (v9372 & ~i22),
  v9372 = (v9373 & i29) | ~i29,
  v9373 = (v9374 & ~i30) | i30,
  v9374 = (v9375 & i31) | ~i31,
  v9375 = (v9376 & i32) | ~i32,
  v9376 = (v9383 & i35) | (v9377 & ~i35),
  v9377 = (v9382 & i36) | (v9378 & ~i36),
  v9378 = (v9381 & i37) | (v9379 & ~i37),
  v9379 = (v9380 & i38) | (v8955 & ~i38),
  v9380 = (v9297 & i40) | (v9050 & ~i40),
  v9381 = (v9380 & i38) | ~i38,
  v9382 = (v9381 & i37) | (v9380 & ~i37),
  v9383 = (v9382 & i36) | (v9384 & ~i36),
  v9384 = (v9381 & i37) | (v9385 & ~i37),
  v9385 = (v9380 & i38) | (v9386 & ~i38),
  v9386 = (v9380 & i39) | (v8955 & ~i39),
  v9387 = (v9393 & i25) | (v9388 & ~i25),
  v9388 = (v9389 & i29) | ~i29,
  v9389 = (v9392 & i30) | (v9390 & ~i30),
  v9390 = (v9391 & i31) | (v801 & ~i31),
  v9391 = (v9376 & i32) | (v9360 & ~i32),
  v9392 = (v9111 & i32) | (v805 & ~i32),
  v9393 = (v9389 & i29) | (v9394 & ~i29),
  v9394 = (v9395 & ~i30) | i30,
  v9395 = (v9396 & ~i31) | i31,
  v9396 = (v801 & ~i32) | i32,
  v9397 = (v9485 & i19) | (v9398 & ~i19),
  v9398 = (v9442 & i20) | (v9399 & ~i20),
  v9399 = (v9416 & i21) | (v9400 & ~i21),
  v9400 = (v9401 & i22) | ~i22,
  v9401 = (v9402 & i29) | ~i29,
  v9402 = (v9403 & ~i30) | i30,
  v9403 = (v9404 & i31) | ~i31,
  v9404 = (v9405 & ~i32) | i32,
  v9405 = (v9413 & i35) | (v9406 & ~i35),
  v9406 = (v9412 & i36) | (v9407 & ~i36),
  v9407 = (v9411 & i37) | (v9408 & ~i37),
  v9408 = (v9410 & i38) | (v9409 & ~i38),
  v9409 = (v8938 & i39) | (v9410 & ~i39),
  v9410 = (v9031 & i40) | (v9250 & ~i40),
  v9411 = (v9410 & i38) | ~i38,
  v9412 = (v9411 & i37) | (v9410 & ~i37),
  v9413 = (v9412 & i36) | (v9414 & ~i36),
  v9414 = (v9411 & i37) | (v9415 & ~i37),
  v9415 = (v9410 & i38) | (v8938 & ~i38),
  v9416 = (v9432 & i22) | (v9417 & ~i22),
  v9417 = (v9418 & i29) | ~i29,
  v9418 = (v9419 & ~i30) | i30,
  v9419 = (v9420 & i31) | ~i31,
  v9420 = (v9421 & i32) | ~i32,
  v9421 = (v9429 & i35) | (v9422 & ~i35),
  v9422 = (v9428 & i36) | (v9423 & ~i36),
  v9423 = (v9427 & i37) | (v9424 & ~i37),
  v9424 = (v9426 & i38) | (v9425 & ~i38),
  v9425 = (v8955 & i39) | (v9426 & ~i39),
  v9426 = (v9050 & i40) | (v9262 & ~i40),
  v9427 = (v9426 & i38) | ~i38,
  v9428 = (v9427 & i37) | (v9426 & ~i37),
  v9429 = (v9428 & i36) | (v9430 & ~i36),
  v9430 = (v9427 & i37) | (v9431 & ~i37),
  v9431 = (v9426 & i38) | (v8955 & ~i38),
  v9432 = (v9438 & i25) | (v9433 & ~i25),
  v9433 = (v9434 & i29) | ~i29,
  v9434 = (v9437 & i30) | (v9435 & ~i30),
  v9435 = (v9436 & i31) | (v821 & ~i31),
  v9436 = (v9421 & i32) | (v9405 & ~i32),
  v9437 = (v9157 & i32) | (v826 & ~i32),
  v9438 = (v9434 & i29) | (v9439 & ~i29),
  v9439 = (v9440 & ~i30) | i30,
  v9440 = (v9441 & ~i31) | i31,
  v9441 = (v821 & ~i32) | i32,
  v9442 = (v9459 & i21) | (v9443 & ~i21),
  v9443 = (v9444 & i22) | ~i22,
  v9444 = (v9445 & i29) | ~i29,
  v9445 = (v9446 & ~i30) | i30,
  v9446 = (v9447 & i31) | ~i31,
  v9447 = (v9448 & ~i32) | i32,
  v9448 = (v9456 & i35) | (v9449 & ~i35),
  v9449 = (v9455 & i36) | (v9450 & ~i36),
  v9450 = (v9454 & i37) | (v9451 & ~i37),
  v9451 = (v9453 & i38) | (v9452 & ~i38),
  v9452 = (v9453 & i39) | (v8938 & ~i39),
  v9453 = (v9031 & i40) | (v9285 & ~i40),
  v9454 = (v9453 & i38) | ~i38,
  v9455 = (v9454 & i37) | (v9453 & ~i37),
  v9456 = (v9455 & i36) | (v9457 & ~i36),
  v9457 = (v9454 & i37) | (v9458 & ~i37),
  v9458 = (v9453 & i38) | (v8938 & ~i38),
  v9459 = (v9475 & i22) | (v9460 & ~i22),
  v9460 = (v9461 & i29) | ~i29,
  v9461 = (v9462 & ~i30) | i30,
  v9462 = (v9463 & i31) | ~i31,
  v9463 = (v9464 & i32) | ~i32,
  v9464 = (v9472 & i35) | (v9465 & ~i35),
  v9465 = (v9471 & i36) | (v9466 & ~i36),
  v9466 = (v9470 & i37) | (v9467 & ~i37),
  v9467 = (v9469 & i38) | (v9468 & ~i38),
  v9468 = (v9469 & i39) | (v8955 & ~i39),
  v9469 = (v9050 & i40) | (v9297 & ~i40),
  v9470 = (v9469 & i38) | ~i38,
  v9471 = (v9470 & i37) | (v9469 & ~i37),
  v9472 = (v9471 & i36) | (v9473 & ~i36),
  v9473 = (v9470 & i37) | (v9474 & ~i37),
  v9474 = (v9469 & i38) | (v8955 & ~i38),
  v9475 = (v9481 & i25) | (v9476 & ~i25),
  v9476 = (v9477 & i29) | ~i29,
  v9477 = (v9480 & i30) | (v9478 & ~i30),
  v9478 = (v9479 & i31) | (v839 & ~i31),
  v9479 = (v9464 & i32) | (v9448 & ~i32),
  v9480 = (v9201 & i32) | (v844 & ~i32),
  v9481 = (v9477 & i29) | (v9482 & ~i29),
  v9482 = (v9483 & ~i30) | i30,
  v9483 = (v9484 & ~i31) | i31,
  v9484 = (v839 & ~i32) | i32,
  v9485 = (v9496 & i21) | (v9486 & ~i21),
  v9486 = (v9487 & i22) | ~i22,
  v9487 = (v9488 & i29) | ~i29,
  v9488 = (v9489 & ~i30) | i30,
  v9489 = (v9490 & i31) | ~i31,
  v9490 = (v9491 & ~i32) | i32,
  v9491 = (v9495 & i36) | (v9492 & ~i36),
  v9492 = (v9494 & i37) | (v9493 & ~i37),
  v9493 = (v9031 & i38) | (v8938 & ~i38),
  v9494 = (v9031 & i38) | ~i38,
  v9495 = (v9494 & i37) | (v9031 & ~i37),
  v9496 = (v9506 & i22) | (v9497 & ~i22),
  v9497 = (v9498 & i29) | ~i29,
  v9498 = (v9499 & ~i30) | i30,
  v9499 = (v9500 & i31) | ~i31,
  v9500 = (v9501 & i32) | ~i32,
  v9501 = (v9505 & i36) | (v9502 & ~i36),
  v9502 = (v9504 & i37) | (v9503 & ~i37),
  v9503 = (v9050 & i38) | (v8955 & ~i38),
  v9504 = (v9050 & i38) | ~i38,
  v9505 = (v9504 & i37) | (v9050 & ~i37),
  v9506 = (v9512 & i25) | (v9507 & ~i25),
  v9507 = (v9508 & i29) | ~i29,
  v9508 = (v9511 & i30) | (v9509 & ~i30),
  v9509 = (v9510 & i31) | (v857 & ~i31),
  v9510 = (v9501 & i32) | (v9491 & ~i32),
  v9511 = (v9065 & i32) | (v668 & ~i32),
  v9512 = (v9508 & i29) | (v9513 & ~i29),
  v9513 = (v9514 & ~i30) | i30,
  v9514 = (v9515 & ~i31) | i31,
  v9515 = (v857 & ~i32) | i32,
  v9516 = (v9704 & i16) | (v9517 & ~i16),
  v9517 = (v9629 & i17) | (v9518 & ~i17),
  v9518 = (v9576 & i19) | (v9519 & ~i19),
  v9519 = (v9548 & i20) | (v9520 & ~i20),
  v9520 = (v9529 & i21) | (v9521 & ~i21),
  v9521 = (v9522 & i22) | ~i22,
  v9522 = (v9523 & i29) | ~i29,
  v9523 = (v9524 & ~i30) | i30,
  v9524 = (v9525 & i31) | ~i31,
  v9525 = (v9526 & ~i32) | i32,
  v9526 = (v9527 & i36) | (v8931 & ~i36),
  v9527 = (v8940 & i37) | (v9528 & ~i37),
  v9528 = (v8934 & i38) | (v8938 & ~i38),
  v9529 = (v9537 & i22) | (v9530 & ~i22),
  v9530 = (v9531 & i29) | ~i29,
  v9531 = (v9532 & ~i30) | i30,
  v9532 = (v9533 & i31) | ~i31,
  v9533 = (v9534 & i32) | ~i32,
  v9534 = (v9535 & i36) | (v8948 & ~i36),
  v9535 = (v8957 & i37) | (v9536 & ~i37),
  v9536 = (v8951 & i38) | (v8955 & ~i38),
  v9537 = (v9544 & i25) | (v9538 & ~i25),
  v9538 = (v9539 & i29) | ~i29,
  v9539 = (v9542 & i30) | (v9540 & ~i30),
  v9540 = (v9541 & i31) | (v873 & ~i31),
  v9541 = (v9534 & i32) | (v9526 & ~i32),
  v9542 = (v9543 & i32) | (v628 & ~i32),
  v9543 = (v9066 & i36) | (v8966 & ~i36),
  v9544 = (v9539 & i29) | (v9545 & ~i29),
  v9545 = (v9546 & ~i30) | i30,
  v9546 = (v9547 & ~i31) | i31,
  v9547 = (v873 & ~i32) | i32,
  v9548 = (v9557 & i21) | (v9549 & ~i21),
  v9549 = (v9550 & i22) | ~i22,
  v9550 = (v9551 & i29) | ~i29,
  v9551 = (v9552 & ~i30) | i30,
  v9552 = (v9553 & i31) | ~i31,
  v9553 = (v9554 & ~i32) | i32,
  v9554 = (v9555 & i36) | (v8980 & ~i36),
  v9555 = (v8987 & i37) | (v9556 & ~i37),
  v9556 = (v8983 & i38) | (v8938 & ~i38),
  v9557 = (v9565 & i22) | (v9558 & ~i22),
  v9558 = (v9559 & i29) | ~i29,
  v9559 = (v9560 & ~i30) | i30,
  v9560 = (v9561 & i31) | ~i31,
  v9561 = (v9562 & i32) | ~i32,
  v9562 = (v9563 & i36) | (v8995 & ~i36),
  v9563 = (v9002 & i37) | (v9564 & ~i37),
  v9564 = (v8998 & i38) | (v8955 & ~i38),
  v9565 = (v9572 & i25) | (v9566 & ~i25),
  v9566 = (v9567 & i29) | ~i29,
  v9567 = (v9570 & i30) | (v9568 & ~i30),
  v9568 = (v9569 & i31) | (v883 & ~i31),
  v9569 = (v9562 & i32) | (v9554 & ~i32),
  v9570 = (v9571 & i32) | (v648 & ~i32),
  v9571 = (v9066 & i36) | (v9011 & ~i36),
  v9572 = (v9567 & i29) | (v9573 & ~i29),
  v9573 = (v9574 & ~i30) | i30,
  v9574 = (v9575 & ~i31) | i31,
  v9575 = (v883 & ~i32) | i32,
  v9576 = (v9603 & i20) | (v9577 & ~i20),
  v9577 = (v9585 & i21) | (v9578 & ~i21),
  v9578 = (v9579 & i22) | ~i22,
  v9579 = (v9580 & i29) | ~i29,
  v9580 = (v9581 & ~i30) | i30,
  v9581 = (v9582 & i31) | ~i31,
  v9582 = (v9583 & ~i32) | i32,
  v9583 = (v9584 & i35) | (v9027 & ~i35),
  v9584 = (v9027 & i36) | (v9036 & ~i36),
  v9585 = (v9592 & i22) | (v9586 & ~i22),
  v9586 = (v9587 & i29) | ~i29,
  v9587 = (v9588 & ~i30) | i30,
  v9588 = (v9589 & i31) | ~i31,
  v9589 = (v9590 & i32) | ~i32,
  v9590 = (v9591 & i35) | (v9046 & ~i35),
  v9591 = (v9046 & i36) | (v9055 & ~i36),
  v9592 = (v9599 & i25) | (v9593 & ~i25),
  v9593 = (v9594 & i29) | ~i29,
  v9594 = (v9597 & i30) | (v9595 & ~i30),
  v9595 = (v9596 & i31) | (v894 & ~i31),
  v9596 = (v9590 & i32) | (v9583 & ~i32),
  v9597 = (v9598 & i32) | (v666 & ~i32),
  v9598 = (v9543 & i35) | (v9066 & ~i35),
  v9599 = (v9594 & i29) | (v9600 & ~i29),
  v9600 = (v9601 & ~i30) | i30,
  v9601 = (v9602 & ~i31) | i31,
  v9602 = (v894 & ~i32) | i32,
  v9603 = (v9611 & i21) | (v9604 & ~i21),
  v9604 = (v9605 & i22) | ~i22,
  v9605 = (v9606 & i29) | ~i29,
  v9606 = (v9607 & ~i30) | i30,
  v9607 = (v9608 & i31) | ~i31,
  v9608 = (v9609 & ~i32) | i32,
  v9609 = (v9610 & i35) | (v9080 & ~i35),
  v9610 = (v9080 & i36) | (v9086 & ~i36),
  v9611 = (v9618 & i22) | (v9612 & ~i22),
  v9612 = (v9613 & i29) | ~i29,
  v9613 = (v9614 & ~i30) | i30,
  v9614 = (v9615 & i31) | ~i31,
  v9615 = (v9616 & i32) | ~i32,
  v9616 = (v9617 & i35) | (v9096 & ~i35),
  v9617 = (v9096 & i36) | (v9102 & ~i36),
  v9618 = (v9625 & i25) | (v9619 & ~i25),
  v9619 = (v9620 & i29) | ~i29,
  v9620 = (v9623 & i30) | (v9621 & ~i30),
  v9621 = (v9622 & i31) | (v903 & ~i31),
  v9622 = (v9616 & i32) | (v9609 & ~i32),
  v9623 = (v9624 & i32) | (v687 & ~i32),
  v9624 = (v9571 & i35) | (v9066 & ~i35),
  v9625 = (v9620 & i29) | (v9626 & ~i29),
  v9626 = (v9627 & ~i30) | i30,
  v9627 = (v9628 & ~i31) | i31,
  v9628 = (v903 & ~i32) | i32,
  v9629 = (v9683 & i19) | (v9630 & ~i19),
  v9630 = (v9657 & i20) | (v9631 & ~i20),
  v9631 = (v9639 & i21) | (v9632 & ~i21),
  v9632 = (v9633 & i22) | ~i22,
  v9633 = (v9634 & i29) | ~i29,
  v9634 = (v9635 & ~i30) | i30,
  v9635 = (v9636 & i31) | ~i31,
  v9636 = (v9637 & ~i32) | i32,
  v9637 = (v9133 & i35) | (v9638 & ~i35),
  v9638 = (v9133 & i36) | (v9126 & ~i36),
  v9639 = (v9646 & i22) | (v9640 & ~i22),
  v9640 = (v9641 & i29) | ~i29,
  v9641 = (v9642 & ~i30) | i30,
  v9642 = (v9643 & i31) | ~i31,
  v9643 = (v9644 & i32) | ~i32,
  v9644 = (v9149 & i35) | (v9645 & ~i35),
  v9645 = (v9149 & i36) | (v9142 & ~i36),
  v9646 = (v9653 & i25) | (v9647 & ~i25),
  v9647 = (v9648 & i29) | ~i29,
  v9648 = (v9651 & i30) | (v9649 & ~i30),
  v9649 = (v9650 & i31) | (v914 & ~i31),
  v9650 = (v9644 & i32) | (v9637 & ~i32),
  v9651 = (v9652 & i32) | (v708 & ~i32),
  v9652 = (v9066 & i35) | (v9543 & ~i35),
  v9653 = (v9648 & i29) | (v9654 & ~i29),
  v9654 = (v9655 & ~i30) | i30,
  v9655 = (v9656 & ~i31) | i31,
  v9656 = (v914 & ~i32) | i32,
  v9657 = (v9665 & i21) | (v9658 & ~i21),
  v9658 = (v9659 & i22) | ~i22,
  v9659 = (v9660 & i29) | ~i29,
  v9660 = (v9661 & ~i30) | i30,
  v9661 = (v9662 & i31) | ~i31,
  v9662 = (v9663 & ~i32) | i32,
  v9663 = (v9177 & i35) | (v9664 & ~i35),
  v9664 = (v9177 & i36) | (v9170 & ~i36),
  v9665 = (v9672 & i22) | (v9666 & ~i22),
  v9666 = (v9667 & i29) | ~i29,
  v9667 = (v9668 & ~i30) | i30,
  v9668 = (v9669 & i31) | ~i31,
  v9669 = (v9670 & i32) | ~i32,
  v9670 = (v9193 & i35) | (v9671 & ~i35),
  v9671 = (v9193 & i36) | (v9186 & ~i36),
  v9672 = (v9679 & i25) | (v9673 & ~i25),
  v9673 = (v9674 & i29) | ~i29,
  v9674 = (v9677 & i30) | (v9675 & ~i30),
  v9675 = (v9676 & i31) | (v923 & ~i31),
  v9676 = (v9670 & i32) | (v9663 & ~i32),
  v9677 = (v9678 & i32) | (v726 & ~i32),
  v9678 = (v9066 & i35) | (v9571 & ~i35),
  v9679 = (v9674 & i29) | (v9680 & ~i29),
  v9680 = (v9681 & ~i30) | i30,
  v9681 = (v9682 & ~i31) | i31,
  v9682 = (v923 & ~i32) | i32,
  v9683 = (v9689 & i21) | (v9684 & ~i21),
  v9684 = (v9685 & i22) | ~i22,
  v9685 = (v9686 & i29) | ~i29,
  v9686 = (v9687 & ~i30) | i30,
  v9687 = (v9688 & i31) | ~i31,
  v9688 = (v9213 & ~i32) | i32,
  v9689 = (v9694 & i22) | (v9690 & ~i22),
  v9690 = (v9691 & i29) | ~i29,
  v9691 = (v9692 & ~i30) | i30,
  v9692 = (v9693 & i31) | ~i31,
  v9693 = (v9223 & i32) | ~i32,
  v9694 = (v9700 & i25) | (v9695 & ~i25),
  v9695 = (v9696 & i29) | ~i29,
  v9696 = (v9699 & i30) | (v9697 & ~i30),
  v9697 = (v9698 & i31) | (v740 & ~i31),
  v9698 = (v9223 & i32) | (v9213 & ~i32),
  v9699 = (v9066 & i32) | (v667 & ~i32),
  v9700 = (v9696 & i29) | (v9701 & ~i29),
  v9701 = (v9702 & ~i30) | i30,
  v9702 = (v9703 & ~i31) | i31,
  v9703 = (v740 & ~i32) | i32,
  v9704 = (v9812 & i17) | (v9705 & ~i17),
  v9705 = (v9761 & i19) | (v9706 & ~i19),
  v9706 = (v9734 & i20) | (v9707 & ~i20),
  v9707 = (v9716 & i21) | (v9708 & ~i21),
  v9708 = (v9709 & i22) | ~i22,
  v9709 = (v9710 & i29) | ~i29,
  v9710 = (v9711 & ~i30) | i30,
  v9711 = (v9712 & i31) | ~i31,
  v9712 = (v9713 & ~i32) | i32,
  v9713 = (v9714 & i36) | (v9247 & ~i36),
  v9714 = (v9251 & i37) | (v9715 & ~i37),
  v9715 = (v9250 & i38) | (v8938 & ~i38),
  v9716 = (v9724 & i22) | (v9717 & ~i22),
  v9717 = (v9718 & i29) | ~i29,
  v9718 = (v9719 & ~i30) | i30,
  v9719 = (v9720 & i31) | ~i31,
  v9720 = (v9721 & i32) | ~i32,
  v9721 = (v9722 & i36) | (v9259 & ~i36),
  v9722 = (v9263 & i37) | (v9723 & ~i37),
  v9723 = (v9262 & i38) | (v8955 & ~i38),
  v9724 = (v9730 & i25) | (v9725 & ~i25),
  v9725 = (v9726 & i29) | ~i29,
  v9726 = (v9729 & i30) | (v9727 & ~i30),
  v9727 = (v9728 & i31) | (v942 & ~i31),
  v9728 = (v9721 & i32) | (v9713 & ~i32),
  v9729 = (v9543 & i32) | (v758 & ~i32),
  v9730 = (v9726 & i29) | (v9731 & ~i29),
  v9731 = (v9732 & ~i30) | i30,
  v9732 = (v9733 & ~i31) | i31,
  v9733 = (v942 & ~i32) | i32,
  v9734 = (v9743 & i21) | (v9735 & ~i21),
  v9735 = (v9736 & i22) | ~i22,
  v9736 = (v9737 & i29) | ~i29,
  v9737 = (v9738 & ~i30) | i30,
  v9738 = (v9739 & i31) | ~i31,
  v9739 = (v9740 & ~i32) | i32,
  v9740 = (v9741 & i36) | (v9282 & ~i36),
  v9741 = (v9286 & i37) | (v9742 & ~i37),
  v9742 = (v9285 & i38) | (v8938 & ~i38),
  v9743 = (v9751 & i22) | (v9744 & ~i22),
  v9744 = (v9745 & i29) | ~i29,
  v9745 = (v9746 & ~i30) | i30,
  v9746 = (v9747 & i31) | ~i31,
  v9747 = (v9748 & i32) | ~i32,
  v9748 = (v9749 & i36) | (v9294 & ~i36),
  v9749 = (v9298 & i37) | (v9750 & ~i37),
  v9750 = (v9297 & i38) | (v8955 & ~i38),
  v9751 = (v9757 & i25) | (v9752 & ~i25),
  v9752 = (v9753 & i29) | ~i29,
  v9753 = (v9756 & i30) | (v9754 & ~i30),
  v9754 = (v9755 & i31) | (v952 & ~i31),
  v9755 = (v9748 & i32) | (v9740 & ~i32),
  v9756 = (v9571 & i32) | (v772 & ~i32),
  v9757 = (v9753 & i29) | (v9758 & ~i29),
  v9758 = (v9759 & ~i30) | i30,
  v9759 = (v9760 & ~i31) | i31,
  v9760 = (v952 & ~i32) | i32,
  v9761 = (v9787 & i20) | (v9762 & ~i20),
  v9762 = (v9770 & i21) | (v9763 & ~i21),
  v9763 = (v9764 & i22) | ~i22,
  v9764 = (v9765 & i29) | ~i29,
  v9765 = (v9766 & ~i30) | i30,
  v9766 = (v9767 & i31) | ~i31,
  v9767 = (v9768 & ~i32) | i32,
  v9768 = (v9769 & i35) | (v9319 & ~i35),
  v9769 = (v9319 & i36) | (v9325 & ~i36),
  v9770 = (v9777 & i22) | (v9771 & ~i22),
  v9771 = (v9772 & i29) | ~i29,
  v9772 = (v9773 & ~i30) | i30,
  v9773 = (v9774 & i31) | ~i31,
  v9774 = (v9775 & i32) | ~i32,
  v9775 = (v9776 & i35) | (v9335 & ~i35),
  v9776 = (v9335 & i36) | (v9341 & ~i36),
  v9777 = (v9783 & i25) | (v9778 & ~i25),
  v9778 = (v9779 & i29) | ~i29,
  v9779 = (v9782 & i30) | (v9780 & ~i30),
  v9780 = (v9781 & i31) | (v963 & ~i31),
  v9781 = (v9775 & i32) | (v9768 & ~i32),
  v9782 = (v9598 & i32) | (v787 & ~i32),
  v9783 = (v9779 & i29) | (v9784 & ~i29),
  v9784 = (v9785 & ~i30) | i30,
  v9785 = (v9786 & ~i31) | i31,
  v9786 = (v963 & ~i32) | i32,
  v9787 = (v9795 & i21) | (v9788 & ~i21),
  v9788 = (v9789 & i22) | ~i22,
  v9789 = (v9790 & i29) | ~i29,
  v9790 = (v9791 & ~i30) | i30,
  v9791 = (v9792 & i31) | ~i31,
  v9792 = (v9793 & ~i32) | i32,
  v9793 = (v9794 & i35) | (v9362 & ~i35),
  v9794 = (v9362 & i36) | (v9368 & ~i36),
  v9795 = (v9802 & i22) | (v9796 & ~i22),
  v9796 = (v9797 & i29) | ~i29,
  v9797 = (v9798 & ~i30) | i30,
  v9798 = (v9799 & i31) | ~i31,
  v9799 = (v9800 & i32) | ~i32,
  v9800 = (v9801 & i35) | (v9378 & ~i35),
  v9801 = (v9378 & i36) | (v9384 & ~i36),
  v9802 = (v9808 & i25) | (v9803 & ~i25),
  v9803 = (v9804 & i29) | ~i29,
  v9804 = (v9807 & i30) | (v9805 & ~i30),
  v9805 = (v9806 & i31) | (v972 & ~i31),
  v9806 = (v9800 & i32) | (v9793 & ~i32),
  v9807 = (v9624 & i32) | (v805 & ~i32),
  v9808 = (v9804 & i29) | (v9809 & ~i29),
  v9809 = (v9810 & ~i30) | i30,
  v9810 = (v9811 & ~i31) | i31,
  v9811 = (v972 & ~i32) | i32,
  v9812 = (v9864 & i19) | (v9813 & ~i19),
  v9813 = (v9839 & i20) | (v9814 & ~i20),
  v9814 = (v9822 & i21) | (v9815 & ~i21),
  v9815 = (v9816 & i22) | ~i22,
  v9816 = (v9817 & i29) | ~i29,
  v9817 = (v9818 & ~i30) | i30,
  v9818 = (v9819 & i31) | ~i31,
  v9819 = (v9820 & ~i32) | i32,
  v9820 = (v9414 & i35) | (v9821 & ~i35),
  v9821 = (v9414 & i36) | (v9407 & ~i36),
  v9822 = (v9829 & i22) | (v9823 & ~i22),
  v9823 = (v9824 & i29) | ~i29,
  v9824 = (v9825 & ~i30) | i30,
  v9825 = (v9826 & i31) | ~i31,
  v9826 = (v9827 & i32) | ~i32,
  v9827 = (v9430 & i35) | (v9828 & ~i35),
  v9828 = (v9430 & i36) | (v9423 & ~i36),
  v9829 = (v9835 & i25) | (v9830 & ~i25),
  v9830 = (v9831 & i29) | ~i29,
  v9831 = (v9834 & i30) | (v9832 & ~i30),
  v9832 = (v9833 & i31) | (v983 & ~i31),
  v9833 = (v9827 & i32) | (v9820 & ~i32),
  v9834 = (v9652 & i32) | (v826 & ~i32),
  v9835 = (v9831 & i29) | (v9836 & ~i29),
  v9836 = (v9837 & ~i30) | i30,
  v9837 = (v9838 & ~i31) | i31,
  v9838 = (v983 & ~i32) | i32,
  v9839 = (v9847 & i21) | (v9840 & ~i21),
  v9840 = (v9841 & i22) | ~i22,
  v9841 = (v9842 & i29) | ~i29,
  v9842 = (v9843 & ~i30) | i30,
  v9843 = (v9844 & i31) | ~i31,
  v9844 = (v9845 & ~i32) | i32,
  v9845 = (v9457 & i35) | (v9846 & ~i35),
  v9846 = (v9457 & i36) | (v9450 & ~i36),
  v9847 = (v9854 & i22) | (v9848 & ~i22),
  v9848 = (v9849 & i29) | ~i29,
  v9849 = (v9850 & ~i30) | i30,
  v9850 = (v9851 & i31) | ~i31,
  v9851 = (v9852 & i32) | ~i32,
  v9852 = (v9473 & i35) | (v9853 & ~i35),
  v9853 = (v9473 & i36) | (v9466 & ~i36),
  v9854 = (v9860 & i25) | (v9855 & ~i25),
  v9855 = (v9856 & i29) | ~i29,
  v9856 = (v9859 & i30) | (v9857 & ~i30),
  v9857 = (v9858 & i31) | (v992 & ~i31),
  v9858 = (v9852 & i32) | (v9845 & ~i32),
  v9859 = (v9678 & i32) | (v844 & ~i32),
  v9860 = (v9856 & i29) | (v9861 & ~i29),
  v9861 = (v9862 & ~i30) | i30,
  v9862 = (v9863 & ~i31) | i31,
  v9863 = (v992 & ~i32) | i32,
  v9864 = (v9870 & i21) | (v9865 & ~i21),
  v9865 = (v9866 & i22) | ~i22,
  v9866 = (v9867 & i29) | ~i29,
  v9867 = (v9868 & ~i30) | i30,
  v9868 = (v9869 & i31) | ~i31,
  v9869 = (v9492 & ~i32) | i32,
  v9870 = (v9875 & i22) | (v9871 & ~i22),
  v9871 = (v9872 & i29) | ~i29,
  v9872 = (v9873 & ~i30) | i30,
  v9873 = (v9874 & i31) | ~i31,
  v9874 = (v9502 & i32) | ~i32,
  v9875 = (v9881 & i25) | (v9876 & ~i25),
  v9876 = (v9877 & i29) | ~i29,
  v9877 = (v9880 & i30) | (v9878 & ~i30),
  v9878 = (v9879 & i31) | (v858 & ~i31),
  v9879 = (v9502 & i32) | (v9492 & ~i32),
  v9880 = (v9066 & i32) | (v668 & ~i32),
  v9881 = (v9877 & i29) | (v9882 & ~i29),
  v9882 = (v9883 & ~i30) | i30,
  v9883 = (v9884 & ~i31) | i31,
  v9884 = (v858 & ~i32) | i32,
  v9885 = (v9927 & i15) | (v9886 & ~i15),
  v9886 = (v9907 & i16) | (v9887 & ~i16),
  v9887 = (v9899 & i17) | (v9888 & ~i17),
  v9888 = (v9894 & i19) | (v9889 & ~i19),
  v9889 = (v9892 & i20) | (v9890 & ~i20),
  v9890 = (v9891 & i21) | (v8925 & ~i21),
  v9891 = (v8969 & i22) | (v8943 & ~i22),
  v9892 = (v9893 & i21) | (v8974 & ~i21),
  v9893 = (v9014 & i22) | (v8990 & ~i22),
  v9894 = (v9897 & i20) | (v9895 & ~i20),
  v9895 = (v9896 & i21) | (v9020 & ~i21),
  v9896 = (v9068 & i22) | (v9040 & ~i22),
  v9897 = (v9898 & i21) | (v9073 & ~i21),
  v9898 = (v9112 & i22) | (v9090 & ~i22),
  v9899 = (v9905 & i19) | (v9900 & ~i19),
  v9900 = (v9903 & i20) | (v9901 & ~i20),
  v9901 = (v9902 & i21) | (v9119 & ~i21),
  v9902 = (v9158 & i22) | (v9136 & ~i22),
  v9903 = (v9904 & i21) | (v9163 & ~i21),
  v9904 = (v9202 & i22) | (v9180 & ~i22),
  v9905 = (v9906 & i21) | (v9207 & ~i21),
  v9906 = (v9233 & i22) | (v9218 & ~i22),
  v9907 = (v9919 & i17) | (v9908 & ~i17),
  v9908 = (v9914 & i19) | (v9909 & ~i19),
  v9909 = (v9912 & i20) | (v9910 & ~i20),
  v9910 = (v9911 & i21) | (v9241 & ~i21),
  v9911 = (v9271 & i22) | (v9254 & ~i22),
  v9912 = (v9913 & i21) | (v9276 & ~i21),
  v9913 = (v9306 & i22) | (v9289 & ~i22),
  v9914 = (v9917 & i20) | (v9915 & ~i20),
  v9915 = (v9916 & i21) | (v9312 & ~i21),
  v9916 = (v9350 & i22) | (v9329 & ~i22),
  v9917 = (v9918 & i21) | (v9355 & ~i21),
  v9918 = (v9393 & i22) | (v9372 & ~i22),
  v9919 = (v9925 & i19) | (v9920 & ~i19),
  v9920 = (v9923 & i20) | (v9921 & ~i20),
  v9921 = (v9922 & i21) | (v9400 & ~i21),
  v9922 = (v9438 & i22) | (v9417 & ~i22),
  v9923 = (v9924 & i21) | (v9443 & ~i21),
  v9924 = (v9481 & i22) | (v9460 & ~i22),
  v9925 = (v9926 & i21) | (v9486 & ~i21),
  v9926 = (v9512 & i22) | (v9497 & ~i22),
  v9927 = (v9948 & i16) | (v9928 & ~i16),
  v9928 = (v9940 & i17) | (v9929 & ~i17),
  v9929 = (v9935 & i19) | (v9930 & ~i19),
  v9930 = (v9933 & i20) | (v9931 & ~i20),
  v9931 = (v9932 & i21) | (v9521 & ~i21),
  v9932 = (v9544 & i22) | (v9530 & ~i22),
  v9933 = (v9934 & i21) | (v9549 & ~i21),
  v9934 = (v9572 & i22) | (v9558 & ~i22),
  v9935 = (v9938 & i20) | (v9936 & ~i20),
  v9936 = (v9937 & i21) | (v9578 & ~i21),
  v9937 = (v9599 & i22) | (v9586 & ~i22),
  v9938 = (v9939 & i21) | (v9604 & ~i21),
  v9939 = (v9625 & i22) | (v9612 & ~i22),
  v9940 = (v9946 & i19) | (v9941 & ~i19),
  v9941 = (v9944 & i20) | (v9942 & ~i20),
  v9942 = (v9943 & i21) | (v9632 & ~i21),
  v9943 = (v9653 & i22) | (v9640 & ~i22),
  v9944 = (v9945 & i21) | (v9658 & ~i21),
  v9945 = (v9679 & i22) | (v9666 & ~i22),
  v9946 = (v9947 & i21) | (v9684 & ~i21),
  v9947 = (v9700 & i22) | (v9690 & ~i22),
  v9948 = (v9960 & i17) | (v9949 & ~i17),
  v9949 = (v9955 & i19) | (v9950 & ~i19),
  v9950 = (v9953 & i20) | (v9951 & ~i20),
  v9951 = (v9952 & i21) | (v9708 & ~i21),
  v9952 = (v9730 & i22) | (v9717 & ~i22),
  v9953 = (v9954 & i21) | (v9735 & ~i21),
  v9954 = (v9757 & i22) | (v9744 & ~i22),
  v9955 = (v9958 & i20) | (v9956 & ~i20),
  v9956 = (v9957 & i21) | (v9763 & ~i21),
  v9957 = (v9783 & i22) | (v9771 & ~i22),
  v9958 = (v9959 & i21) | (v9788 & ~i21),
  v9959 = (v9808 & i22) | (v9796 & ~i22),
  v9960 = (v9966 & i19) | (v9961 & ~i19),
  v9961 = (v9964 & i20) | (v9962 & ~i20),
  v9962 = (v9963 & i21) | (v9815 & ~i21),
  v9963 = (v9835 & i22) | (v9823 & ~i22),
  v9964 = (v9965 & i21) | (v9840 & ~i21),
  v9965 = (v9860 & i22) | (v9848 & ~i22),
  v9966 = (v9967 & i21) | (v9865 & ~i21),
  v9967 = (v9881 & i22) | (v9871 & ~i22),
  v9968 = (v9972 & i11) | (v9969 & ~i11),
  v9969 = (v9972 & i12) | (v9970 & ~i12),
  v9970 = (v9972 & i13) | (v9971 & ~i13),
  v9971 = (v9885 & i14) | (v9972 & ~i14),
  v9972 = (v10014 & i15) | (v9973 & ~i15),
  v9973 = (v9994 & i16) | (v9974 & ~i16),
  v9974 = (v9986 & i17) | (v9975 & ~i17),
  v9975 = (v9981 & i19) | (v9976 & ~i19),
  v9976 = (v9979 & i20) | (v9977 & ~i20),
  v9977 = (v9978 & i21) | (v8925 & ~i21),
  v9978 = (v8960 & i22) | (v8943 & ~i22),
  v9979 = (v9980 & i21) | (v8974 & ~i21),
  v9980 = (v9005 & i22) | (v8990 & ~i22),
  v9981 = (v9984 & i20) | (v9982 & ~i20),
  v9982 = (v9983 & i21) | (v9020 & ~i21),
  v9983 = (v9059 & i22) | (v9040 & ~i22),
  v9984 = (v9985 & i21) | (v9073 & ~i21),
  v9985 = (v9106 & i22) | (v9090 & ~i22),
  v9986 = (v9992 & i19) | (v9987 & ~i19),
  v9987 = (v9990 & i20) | (v9988 & ~i20),
  v9988 = (v9989 & i21) | (v9119 & ~i21),
  v9989 = (v9152 & i22) | (v9136 & ~i22),
  v9990 = (v9991 & i21) | (v9163 & ~i21),
  v9991 = (v9196 & i22) | (v9180 & ~i22),
  v9992 = (v9993 & i21) | (v9207 & ~i21),
  v9993 = (v9228 & i22) | (v9218 & ~i22),
  v9994 = (v10006 & i17) | (v9995 & ~i17),
  v9995 = (v10001 & i19) | (v9996 & ~i19),
  v9996 = (v9999 & i20) | (v9997 & ~i20),
  v9997 = (v9998 & i21) | (v9241 & ~i21),
  v9998 = (v9266 & i22) | (v9254 & ~i22),
  v9999 = (v10000 & i21) | (v9276 & ~i21),
  i28 = \IN-i28 ,
  i49 = \IN-i49 ,
  i50 = \IN-i50 ,
  i51 = \IN-i51 ,
  i52 = \IN-i52 ,
  i53 = \IN-i53 ,
  i54 = \IN-i54 ,
  i55 = \IN-i55 ,
  i56 = \IN-i56 ,
  i57 = \IN-i57 ,
  i58 = \IN-i58 ,
  i59 = \IN-i59 ,
  i60 = \IN-i60 ,
  i61 = \IN-i61 ,
  i62 = \IN-i62 ,
  i63 = \IN-i63 ,
  i64 = \IN-i64 ,
  i65 = \IN-i65 ,
  i66 = \IN-i66 ,
  i67 = \IN-i67 ,
  i68 = \IN-i68 ,
  i69 = \IN-i69 ,
  i70 = \IN-i70 ,
  i71 = \IN-i71 ,
  i72 = \IN-i72 ,
  i73 = \IN-i73 ,
  i74 = \IN-i74 ,
  i75 = \IN-i75 ,
  i76 = \IN-i76 ,
  i77 = \IN-i77 ,
  i78 = \IN-i78 ,
  i79 = \IN-i79 ,
  i80 = \IN-i80 ,
  i81 = \IN-i81 ,
  i82 = \IN-i82 ,
  i83 = \IN-i83 ,
  i84 = \IN-i84 ,
  i85 = \IN-i85 ,
  i86 = \IN-i86 ,
  i87 = \IN-i87 ,
  i88 = \IN-i88 ,
  i89 = \IN-i89 ,
  i90 = \IN-i90 ,
  i91 = \IN-i91 ,
  i92 = \IN-i92 ,
  i93 = \IN-i93 ,
  i94 = \IN-i94 ,
  i95 = \IN-i95 ,
  i96 = \IN-i96 ,
  i97 = \IN-i97 ,
  i98 = \IN-i98 ,
  i99 = \IN-i99 ,
  v10 = (v12 & i30) | (v11 & ~i30),
  v11 = (v13 & i31) | (v12 & ~i31),
  v12 = (v7 & i47) | ~i47,
  v13 = (v7 & i32) | (v12 & ~i32),
  v14 = (v16 & i2) | (v15 & ~i2),
  v15 = (v21 & i3) | (v16 & ~i3),
  v16 = (v20 & i22) | (v17 & ~i22),
  v17 = (v18 & ~i30) | i30,
  v18 = (v19 & i31) | ~i31,
  v19 = (v20 & i32) | ~i32,
  v20 = i47,
  v21 = (v16 & i4) | (v22 & ~i4),
  v22 = (v16 & i5) | (v23 & ~i5),
  v23 = (v24 & i6) | (v16 & ~i6),
  v24 = (v28 & i22) | (v25 & ~i22),
  v25 = (~v26 & ~i30) | i30,
  v26 = v27 & i31,
  v27 = i32,
  v28 = (v20 & i30) | (~v29 & ~i30),
  v29 = (v30 & i31) | (~v20 & ~i31),
  v30 = (~v20 & ~i32) | i32,
  v31 = (v38 & i20) | (v32 & ~i20),
  v32 = (v36 & i21) | (v33 & ~i21),
  v33 = (v35 & i30) | (v34 & ~i30),
  v34 = (v37 & i31) | (v35 & ~i31),
  v35 = v36 & i45,
  v36 = i46,
  v37 = (v35 & i32) | (v36 & ~i32),
  v38 = (v36 & i21) | (v39 & ~i21),
  v39 = (v41 & i30) | (v40 & ~i30),
  v40 = (v42 & i31) | (v41 & ~i31),
  v41 = (v36 & i45) | ~i45,
  v42 = (v41 & i32) | (v36 & ~i32),
  v43 = (v45 & i2) | (v44 & ~i2),
  v44 = (v50 & i3) | (v45 & ~i3),
  v45 = (v49 & i21) | (v46 & ~i21),
  v46 = (v47 & ~i30) | i30,
  v47 = (v48 & i31) | ~i31,
  v48 = (v49 & ~i32) | i32,
  v49 = i45,
  v50 = (v45 & i4) | (v51 & ~i4),
  v51 = (v45 & i5) | (v52 & ~i5),
  v52 = (v53 & i6) | (v45 & ~i6),
  v53 = (v56 & i21) | (v54 & ~i21),
  v54 = (v55 & ~i30) | i30,
  v55 = (v27 & i31) | ~i31,
  v56 = (v49 & i30) | (v57 & ~i30),
  v57 = (v58 & i31) | (v49 & ~i31),
  v58 = v49 & i32,
  v59 = (v61 & i30) | (v60 & ~i30),
  v60 = i44,
  v61 = (v60 & i31) | (v62 & ~i31),
  v62 = (v63 & i32) | (v60 & ~i32),
  v63 = i33,
  v64 = (v112 & i16) | (v65 & ~i16),
  v65 = (v96 & i17) | (v66 & ~i17),
  v66 = (v84 & i19) | (v67 & ~i19),
  v67 = (v77 & i20) | (v68 & ~i20),
  v68 = (v74 & i30) | (~v69 & ~i30),
  v69 = (v73 & i41) | (v70 & ~i41),
  v70 = (v72 & i42) | (v71 & ~i42),
  v71 = v60 & i43,
  v72 = i43,
  v73 = v72 & i42,
  v74 = (v76 & i31) | (~v75 & ~i31),
  v75 = (v69 & ~i32) | i32,
  v76 = (~v69 & ~i32) | i32,
  v77 = (v81 & i30) | (~v78 & ~i30),
  v78 = (v73 & i41) | (v79 & ~i41),
  v79 = (v72 & i42) | (~v80 & ~i42),
  v80 = (v60 & i43) | ~i43,
  v81 = (v83 & i31) | (~v82 & ~i31),
  v82 = (v78 & ~i32) | i32,
  v83 = (~v78 & ~i32) | i32,
  v84 = (v91 & i20) | (v85 & ~i20),
  v85 = (v88 & i30) | (~v86 & ~i30),
  v86 = (v69 & i40) | (v87 & ~i40),
  v87 = (v73 & i41) | (v72 & ~i41),
  v88 = (v90 & i31) | (~v89 & ~i31),
  v89 = (v86 & ~i32) | i32,
  v90 = (~v86 & ~i32) | i32,
  v91 = (v93 & i30) | (~v92 & ~i30),
  v92 = (v78 & i40) | (v87 & ~i40),
  v93 = (v95 & i31) | (~v94 & ~i31),
  v94 = (v92 & ~i32) | i32,
  v95 = (~v92 & ~i32) | i32,
  v96 = (v108 & i19) | (v97 & ~i19),
  v97 = (v103 & i20) | (v98 & ~i20),
  v98 = (v100 & i30) | (~v99 & ~i30),
  v99 = (v87 & i40) | (v69 & ~i40),
  v1000 = (~v858 & ~i34) | i34,
  v1001 = (v1309 & i15) | (v1002 & ~i15),
  v1002 = (v1156 & i16) | (v1003 & ~i16),
  v1003 = (v1091 & i17) | (v1004 & ~i17),
  v1004 = (v1048 & i19) | (v1005 & ~i19),
  v1005 = (v1027 & i20) | (v1006 & ~i20),
  v1006 = (v1007 & i21) | (v617 & ~i21),
  v1007 = (v1008 & i22) | (v617 & ~i22),
  v1008 = (v1018 & i25) | (v1009 & ~i25),
  v1009 = (v1014 & i29) | (v1010 & ~i29),
  v1010 = (v617 & i30) | (v1011 & ~i30),
  v1011 = (v617 & i31) | (v1012 & ~i31),
  v1012 = (v617 & i32) | (v1013 & ~i32),
  v1013 = v624 & i34,
  v1014 = (v617 & i30) | (v1015 & ~i30),
  v1015 = (v617 & i31) | (v1016 & ~i31),
  v1016 = (v617 & i32) | (v1017 & ~i32),
  v1017 = (v617 & i33) | (v1013 & ~i33),
  v1018 = (v1023 & i29) | (v1019 & ~i29),
  v1019 = (v617 & i30) | (v1020 & ~i30),
  v1020 = (v617 & i31) | (v1021 & ~i31),
  v1021 = (v617 & i32) | (v1022 & ~i32),
  v1022 = (~v624 & ~i34) | (v624 & i34),
  v1023 = (v617 & i30) | (v1024 & ~i30),
  v1024 = (v617 & i31) | (v1025 & ~i31),
  v1025 = (v617 & i32) | (v1026 & ~i32),
  v1026 = (v623 & i33) | (v1022 & ~i33),
  v1027 = (v1028 & i21) | (v617 & ~i21),
  v1028 = (v1029 & i22) | (v617 & ~i22),
  v1029 = (v1039 & i25) | (v1030 & ~i25),
  v1030 = (v1035 & i29) | (v1031 & ~i29),
  v1031 = (v617 & i30) | (v1032 & ~i30),
  v1032 = (v617 & i31) | (v1033 & ~i31),
  v1033 = (v617 & i32) | (v1034 & ~i32),
  v1034 = v644 & i34,
  v1035 = (v617 & i30) | (v1036 & ~i30),
  v1036 = (v617 & i31) | (v1037 & ~i31),
  v1037 = (v617 & i32) | (v1038 & ~i32),
  v1038 = (v617 & i33) | (v1034 & ~i33),
  v1039 = (v1044 & i29) | (v1040 & ~i29),
  v1040 = (v617 & i30) | (v1041 & ~i30),
  v1041 = (v617 & i31) | (v1042 & ~i31),
  v1042 = (v617 & i32) | (v1043 & ~i32),
  v1043 = (~v644 & ~i34) | (v644 & i34),
  v1044 = (v617 & i30) | (v1045 & ~i30),
  v1045 = (v617 & i31) | (v1046 & ~i31),
  v1046 = (v617 & i32) | (v1047 & ~i32),
  v1047 = (v643 & i33) | (v1043 & ~i33),
  v1048 = (v1070 & i20) | (v1049 & ~i20),
  v1049 = (v1050 & i21) | (v617 & ~i21),
  v1050 = (v1051 & i22) | (v617 & ~i22),
  v1051 = (v1061 & i25) | (v1052 & ~i25),
  v1052 = (v1057 & i29) | (v1053 & ~i29),
  v1053 = (v617 & i30) | (v1054 & ~i30),
  v1054 = (v617 & i31) | (v1055 & ~i31),
  v1055 = (v617 & i32) | (v1056 & ~i32),
  v1056 = v662 & i34,
  v1057 = (v617 & i30) | (v1058 & ~i30),
  v1058 = (v617 & i31) | (v1059 & ~i31),
  v1059 = (v617 & i32) | (v1060 & ~i32),
  v1060 = (v617 & i33) | (v1056 & ~i33),
  v1061 = (v1066 & i29) | (v1062 & ~i29),
  v1062 = (v617 & i30) | (v1063 & ~i30),
  v1063 = (v617 & i31) | (v1064 & ~i31),
  v1064 = (v617 & i32) | (v1065 & ~i32),
  v1065 = (~v662 & ~i34) | (v662 & i34),
  v1066 = (v617 & i30) | (v1067 & ~i30),
  v1067 = (v617 & i31) | (v1068 & ~i31),
  v1068 = (v617 & i32) | (v1069 & ~i32),
  v1069 = (v661 & i33) | (v1065 & ~i33),
  v1070 = (v1071 & i21) | (v617 & ~i21),
  v1071 = (v1072 & i22) | (v617 & ~i22),
  v1072 = (v1082 & i25) | (v1073 & ~i25),
  v1073 = (v1078 & i29) | (v1074 & ~i29),
  v1074 = (v617 & i30) | (v1075 & ~i30),
  v1075 = (v617 & i31) | (v1076 & ~i31),
  v1076 = (v617 & i32) | (v1077 & ~i32),
  v1077 = v683 & i34,
  v1078 = (v617 & i30) | (v1079 & ~i30),
  v1079 = (v617 & i31) | (v1080 & ~i31),
  v1080 = (v617 & i32) | (v1081 & ~i32),
  v1081 = (v617 & i33) | (v1077 & ~i33),
  v1082 = (v1087 & i29) | (v1083 & ~i29),
  v1083 = (v617 & i30) | (v1084 & ~i30),
  v1084 = (v617 & i31) | (v1085 & ~i31),
  v1085 = (v617 & i32) | (v1086 & ~i32),
  v1086 = (~v683 & ~i34) | (v683 & i34),
  v1087 = (v617 & i30) | (v1088 & ~i30),
  v1088 = (v617 & i31) | (v1089 & ~i31),
  v1089 = (v617 & i32) | (v1090 & ~i32),
  v1090 = (v682 & i33) | (v1086 & ~i33),
  v1091 = (v1135 & i19) | (v1092 & ~i19),
  v1092 = (v1114 & i20) | (v1093 & ~i20),
  v1093 = (v1094 & i21) | (v617 & ~i21),
  v1094 = (v1095 & i22) | (v617 & ~i22),
  v1095 = (v1105 & i25) | (v1096 & ~i25),
  v1096 = (v1101 & i29) | (v1097 & ~i29),
  v1097 = (v617 & i30) | (v1098 & ~i30),
  v1098 = (v617 & i31) | (v1099 & ~i31),
  v1099 = (v617 & i32) | (v1100 & ~i32),
  v1100 = v703 & i34,
  v1101 = (v617 & i30) | (v1102 & ~i30),
  v1102 = (v617 & i31) | (v1103 & ~i31),
  v1103 = (v617 & i32) | (v1104 & ~i32),
  v1104 = (v617 & i33) | (v1100 & ~i33),
  v1105 = (v1110 & i29) | (v1106 & ~i29),
  v1106 = (v617 & i30) | (v1107 & ~i30),
  v1107 = (v617 & i31) | (v1108 & ~i31),
  v1108 = (v617 & i32) | (v1109 & ~i32),
  v1109 = (~v703 & ~i34) | (v703 & i34),
  v1110 = (v617 & i30) | (v1111 & ~i30),
  v1111 = (v617 & i31) | (v1112 & ~i31),
  v1112 = (v617 & i32) | (v1113 & ~i32),
  v1113 = (v702 & i33) | (v1109 & ~i33),
  v1114 = (v1115 & i21) | (v617 & ~i21),
  v1115 = (v1116 & i22) | (v617 & ~i22),
  v1116 = (v1126 & i25) | (v1117 & ~i25),
  v1117 = (v1122 & i29) | (v1118 & ~i29),
  v1118 = (v617 & i30) | (v1119 & ~i30),
  v1119 = (v617 & i31) | (v1120 & ~i31),
  v1120 = (v617 & i32) | (v1121 & ~i32),
  v1121 = v721 & i34,
  v1122 = (v617 & i30) | (v1123 & ~i30),
  v1123 = (v617 & i31) | (v1124 & ~i31),
  v1124 = (v617 & i32) | (v1125 & ~i32),
  v1125 = (v617 & i33) | (v1121 & ~i33),
  v1126 = (v1131 & i29) | (v1127 & ~i29),
  v1127 = (v617 & i30) | (v1128 & ~i30),
  v1128 = (v617 & i31) | (v1129 & ~i31),
  v1129 = (v617 & i32) | (v1130 & ~i32),
  v1130 = (~v721 & ~i34) | (v721 & i34),
  v1131 = (v617 & i30) | (v1132 & ~i30),
  v1132 = (v617 & i31) | (v1133 & ~i31),
  v1133 = (v617 & i32) | (v1134 & ~i32),
  v1134 = (v720 & i33) | (v1130 & ~i33),
  v1135 = (v1136 & i21) | (v617 & ~i21),
  v1136 = (v1137 & i22) | (v617 & ~i22),
  v1137 = (v1147 & i25) | (v1138 & ~i25),
  v1138 = (v1143 & i29) | (v1139 & ~i29),
  v1139 = (v617 & i30) | (v1140 & ~i30),
  v1140 = (v617 & i31) | (v1141 & ~i31),
  v1141 = (v617 & i32) | (v1142 & ~i32),
  v1142 = v739 & i34,
  v1143 = (v617 & i30) | (v1144 & ~i30),
  v1144 = (v617 & i31) | (v1145 & ~i31),
  v1145 = (v617 & i32) | (v1146 & ~i32),
  v1146 = (v617 & i33) | (v1142 & ~i33),
  v1147 = (v1152 & i29) | (v1148 & ~i29),
  v1148 = (v617 & i30) | (v1149 & ~i30),
  v1149 = (v617 & i31) | (v1150 & ~i31),
  v1150 = (v617 & i32) | (v1151 & ~i32),
  v1151 = (~v739 & ~i34) | (v739 & i34),
  v1152 = (v617 & i30) | (v1153 & ~i30),
  v1153 = (v617 & i31) | (v1154 & ~i31),
  v1154 = (v617 & i32) | (v1155 & ~i32),
  v1155 = (v738 & i33) | (v1151 & ~i33),
  v1156 = (v1244 & i17) | (v1157 & ~i17),
  v1157 = (v1201 & i19) | (v1158 & ~i19),
  v1158 = (v1180 & i20) | (v1159 & ~i20),
  v1159 = (v1160 & i21) | (v617 & ~i21),
  v1160 = (v1161 & i22) | (v617 & ~i22),
  v1161 = (v1171 & i25) | (v1162 & ~i25),
  v1162 = (v1167 & i29) | (v1163 & ~i29),
  v1163 = (v617 & i30) | (v1164 & ~i30),
  v1164 = (v617 & i31) | (v1165 & ~i31),
  v1165 = (v617 & i32) | (v1166 & ~i32),
  v1166 = v754 & i34,
  v1167 = (v617 & i30) | (v1168 & ~i30),
  v1168 = (v617 & i31) | (v1169 & ~i31),
  v1169 = (v617 & i32) | (v1170 & ~i32),
  v1170 = (v617 & i33) | (v1166 & ~i33),
  v1171 = (v1176 & i29) | (v1172 & ~i29),
  v1172 = (v617 & i30) | (v1173 & ~i30),
  v1173 = (v617 & i31) | (v1174 & ~i31),
  v1174 = (v617 & i32) | (v1175 & ~i32),
  v1175 = (~v754 & ~i34) | (v754 & i34),
  v1176 = (v617 & i30) | (v1177 & ~i30),
  v1177 = (v617 & i31) | (v1178 & ~i31),
  v1178 = (v617 & i32) | (v1179 & ~i32),
  v1179 = (v753 & i33) | (v1175 & ~i33),
  v1180 = (v1181 & i21) | (v617 & ~i21),
  v1181 = (v1182 & i22) | (v617 & ~i22),
  v1182 = (v1192 & i25) | (v1183 & ~i25),
  v1183 = (v1188 & i29) | (v1184 & ~i29),
  v1184 = (v617 & i30) | (v1185 & ~i30),
  v1185 = (v617 & i31) | (v1186 & ~i31),
  v1186 = (v617 & i32) | (v1187 & ~i32),
  v1187 = v768 & i34,
  v1188 = (v617 & i30) | (v1189 & ~i30),
  v1189 = (v617 & i31) | (v1190 & ~i31),
  v1190 = (v617 & i32) | (v1191 & ~i32),
  v1191 = (v617 & i33) | (v1187 & ~i33),
  v1192 = (v1197 & i29) | (v1193 & ~i29),
  v1193 = (v617 & i30) | (v1194 & ~i30),
  v1194 = (v617 & i31) | (v1195 & ~i31),
  v1195 = (v617 & i32) | (v1196 & ~i32),
  v1196 = (~v768 & ~i34) | (v768 & i34),
  v1197 = (v617 & i30) | (v1198 & ~i30),
  v1198 = (v617 & i31) | (v1199 & ~i31),
  v1199 = (v617 & i32) | (v1200 & ~i32),
  v1200 = (v767 & i33) | (v1196 & ~i33),
  v1201 = (v1223 & i20) | (v1202 & ~i20),
  v1202 = (v1203 & i21) | (v617 & ~i21),
  v1203 = (v1204 & i22) | (v617 & ~i22),
  v1204 = (v1214 & i25) | (v1205 & ~i25),
  v1205 = (v1210 & i29) | (v1206 & ~i29),
  v1206 = (v617 & i30) | (v1207 & ~i30),
  v1207 = (v617 & i31) | (v1208 & ~i31),
  v1208 = (v617 & i32) | (v1209 & ~i32),
  v1209 = v783 & i34,
  v1210 = (v617 & i30) | (v1211 & ~i30),
  v1211 = (v617 & i31) | (v1212 & ~i31),
  v1212 = (v617 & i32) | (v1213 & ~i32),
  v1213 = (v617 & i33) | (v1209 & ~i33),
  v1214 = (v1219 & i29) | (v1215 & ~i29),
  v1215 = (v617 & i30) | (v1216 & ~i30),
  v1216 = (v617 & i31) | (v1217 & ~i31),
  v1217 = (v617 & i32) | (v1218 & ~i32),
  v1218 = (~v783 & ~i34) | (v783 & i34),
  v1219 = (v617 & i30) | (v1220 & ~i30),
  v1220 = (v617 & i31) | (v1221 & ~i31),
  v1221 = (v617 & i32) | (v1222 & ~i32),
  v1222 = (v782 & i33) | (v1218 & ~i33),
  v1223 = (v1224 & i21) | (v617 & ~i21),
  v1224 = (v1225 & i22) | (v617 & ~i22),
  v1225 = (v1235 & i25) | (v1226 & ~i25),
  v1226 = (v1231 & i29) | (v1227 & ~i29),
  v1227 = (v617 & i30) | (v1228 & ~i30),
  v1228 = (v617 & i31) | (v1229 & ~i31),
  v1229 = (v617 & i32) | (v1230 & ~i32),
  v1230 = v801 & i34,
  v1231 = (v617 & i30) | (v1232 & ~i30),
  v1232 = (v617 & i31) | (v1233 & ~i31),
  v1233 = (v617 & i32) | (v1234 & ~i32),
  v1234 = (v617 & i33) | (v1230 & ~i33),
  v1235 = (v1240 & i29) | (v1236 & ~i29),
  v1236 = (v617 & i30) | (v1237 & ~i30),
  v1237 = (v617 & i31) | (v1238 & ~i31),
  v1238 = (v617 & i32) | (v1239 & ~i32),
  v1239 = (~v801 & ~i34) | (v801 & i34),
  v1240 = (v617 & i30) | (v1241 & ~i30),
  v1241 = (v617 & i31) | (v1242 & ~i31),
  v1242 = (v617 & i32) | (v1243 & ~i32),
  v1243 = (v800 & i33) | (v1239 & ~i33),
  v1244 = (v1288 & i19) | (v1245 & ~i19),
  v1245 = (v1267 & i20) | (v1246 & ~i20),
  v1246 = (v1247 & i21) | (v617 & ~i21),
  v1247 = (v1248 & i22) | (v617 & ~i22),
  v1248 = (v1258 & i25) | (v1249 & ~i25),
  v1249 = (v1254 & i29) | (v1250 & ~i29),
  v1250 = (v617 & i30) | (v1251 & ~i30),
  v1251 = (v617 & i31) | (v1252 & ~i31),
  v1252 = (v617 & i32) | (v1253 & ~i32),
  v1253 = v821 & i34,
  v1254 = (v617 & i30) | (v1255 & ~i30),
  v1255 = (v617 & i31) | (v1256 & ~i31),
  v1256 = (v617 & i32) | (v1257 & ~i32),
  v1257 = (v617 & i33) | (v1253 & ~i33),
  v1258 = (v1263 & i29) | (v1259 & ~i29),
  v1259 = (v617 & i30) | (v1260 & ~i30),
  v1260 = (v617 & i31) | (v1261 & ~i31),
  v1261 = (v617 & i32) | (v1262 & ~i32),
  v1262 = (~v821 & ~i34) | (v821 & i34),
  v1263 = (v617 & i30) | (v1264 & ~i30),
  v1264 = (v617 & i31) | (v1265 & ~i31),
  v1265 = (v617 & i32) | (v1266 & ~i32),
  v1266 = (v820 & i33) | (v1262 & ~i33),
  v1267 = (v1268 & i21) | (v617 & ~i21),
  v1268 = (v1269 & i22) | (v617 & ~i22),
  v1269 = (v1279 & i25) | (v1270 & ~i25),
  v1270 = (v1275 & i29) | (v1271 & ~i29),
  v1271 = (v617 & i30) | (v1272 & ~i30),
  v1272 = (v617 & i31) | (v1273 & ~i31),
  v1273 = (v617 & i32) | (v1274 & ~i32),
  v1274 = v839 & i34,
  v1275 = (v617 & i30) | (v1276 & ~i30),
  v1276 = (v617 & i31) | (v1277 & ~i31),
  v1277 = (v617 & i32) | (v1278 & ~i32),
  v1278 = (v617 & i33) | (v1274 & ~i33),
  v1279 = (v1284 & i29) | (v1280 & ~i29),
  v1280 = (v617 & i30) | (v1281 & ~i30),
  v1281 = (v617 & i31) | (v1282 & ~i31),
  v1282 = (v617 & i32) | (v1283 & ~i32),
  v1283 = (~v839 & ~i34) | (v839 & i34),
  v1284 = (v617 & i30) | (v1285 & ~i30),
  v1285 = (v617 & i31) | (v1286 & ~i31),
  v1286 = (v617 & i32) | (v1287 & ~i32),
  v1287 = (v838 & i33) | (v1283 & ~i33),
  v1288 = (v1289 & i21) | (v617 & ~i21),
  v1289 = (v1290 & i22) | (v617 & ~i22),
  v1290 = (v1300 & i25) | (v1291 & ~i25),
  v1291 = (v1296 & i29) | (v1292 & ~i29),
  v1292 = (v617 & i30) | (v1293 & ~i30),
  v1293 = (v617 & i31) | (v1294 & ~i31),
  v1294 = (v617 & i32) | (v1295 & ~i32),
  v1295 = v857 & i34,
  v1296 = (v617 & i30) | (v1297 & ~i30),
  v1297 = (v617 & i31) | (v1298 & ~i31),
  v1298 = (v617 & i32) | (v1299 & ~i32),
  v1299 = (v617 & i33) | (v1295 & ~i33),
  v1300 = (v1305 & i29) | (v1301 & ~i29),
  v1301 = (v617 & i30) | (v1302 & ~i30),
  v1302 = (v617 & i31) | (v1303 & ~i31),
  v1303 = (v617 & i32) | (v1304 & ~i32),
  v1304 = (~v857 & ~i34) | (v857 & i34),
  v1305 = (v617 & i30) | (v1306 & ~i30),
  v1306 = (v617 & i31) | (v1307 & ~i31),
  v1307 = (v617 & i32) | (v1308 & ~i32),
  v1308 = (v856 & i33) | (v1304 & ~i33),
  v1309 = (v1463 & i16) | (v1310 & ~i16),
  v1310 = (v1398 & i17) | (v1311 & ~i17),
  v1311 = (v1355 & i19) | (v1312 & ~i19),
  v1312 = (v1334 & i20) | (v1313 & ~i20),
  v1313 = (v1314 & i21) | (v617 & ~i21),
  v1314 = (v1315 & i22) | (v617 & ~i22),
  v1315 = (v1325 & i25) | (v1316 & ~i25),
  v1316 = (v1321 & i29) | (v1317 & ~i29),
  v1317 = (v617 & i30) | (v1318 & ~i30),
  v1318 = (v617 & i31) | (v1319 & ~i31),
  v1319 = (v617 & i32) | (v1320 & ~i32),
  v1320 = v873 & i34,
  v1321 = (v617 & i30) | (v1322 & ~i30),
  v1322 = (v617 & i31) | (v1323 & ~i31),
  v1323 = (v617 & i32) | (v1324 & ~i32),
  v1324 = (v617 & i33) | (v1320 & ~i33),
  v1325 = (v1330 & i29) | (v1326 & ~i29),
  v1326 = (v617 & i30) | (v1327 & ~i30),
  v1327 = (v617 & i31) | (v1328 & ~i31),
  v1328 = (v617 & i32) | (v1329 & ~i32),
  v1329 = (~v873 & ~i34) | (v873 & i34),
  v1330 = (v617 & i30) | (v1331 & ~i30),
  v1331 = (v617 & i31) | (v1332 & ~i31),
  v1332 = (v617 & i32) | (v1333 & ~i32),
  v1333 = (v872 & i33) | (v1329 & ~i33),
  v1334 = (v1335 & i21) | (v617 & ~i21),
  v1335 = (v1336 & i22) | (v617 & ~i22),
  v1336 = (v1346 & i25) | (v1337 & ~i25),
  v1337 = (v1342 & i29) | (v1338 & ~i29),
  v1338 = (v617 & i30) | (v1339 & ~i30),
  v1339 = (v617 & i31) | (v1340 & ~i31),
  v1340 = (v617 & i32) | (v1341 & ~i32),
  v1341 = v883 & i34,
  v1342 = (v617 & i30) | (v1343 & ~i30),
  v1343 = (v617 & i31) | (v1344 & ~i31),
  v1344 = (v617 & i32) | (v1345 & ~i32),
  v1345 = (v617 & i33) | (v1341 & ~i33),
  v1346 = (v1351 & i29) | (v1347 & ~i29),
  v1347 = (v617 & i30) | (v1348 & ~i30),
  v1348 = (v617 & i31) | (v1349 & ~i31),
  v1349 = (v617 & i32) | (v1350 & ~i32),
  v1350 = (~v883 & ~i34) | (v883 & i34),
  v1351 = (v617 & i30) | (v1352 & ~i30),
  v1352 = (v617 & i31) | (v1353 & ~i31),
  v1353 = (v617 & i32) | (v1354 & ~i32),
  v1354 = (v882 & i33) | (v1350 & ~i33),
  v1355 = (v1377 & i20) | (v1356 & ~i20),
  v1356 = (v1357 & i21) | (v617 & ~i21),
  v1357 = (v1358 & i22) | (v617 & ~i22),
  v1358 = (v1368 & i25) | (v1359 & ~i25),
  v1359 = (v1364 & i29) | (v1360 & ~i29),
  v1360 = (v617 & i30) | (v1361 & ~i30),
  v1361 = (v617 & i31) | (v1362 & ~i31),
  v1362 = (v617 & i32) | (v1363 & ~i32),
  v1363 = v894 & i34,
  v1364 = (v617 & i30) | (v1365 & ~i30),
  v1365 = (v617 & i31) | (v1366 & ~i31),
  v1366 = (v617 & i32) | (v1367 & ~i32),
  v1367 = (v617 & i33) | (v1363 & ~i33),
  v1368 = (v1373 & i29) | (v1369 & ~i29),
  v1369 = (v617 & i30) | (v1370 & ~i30),
  v1370 = (v617 & i31) | (v1371 & ~i31),
  v1371 = (v617 & i32) | (v1372 & ~i32),
  v1372 = (~v894 & ~i34) | (v894 & i34),
  v1373 = (v617 & i30) | (v1374 & ~i30),
  v1374 = (v617 & i31) | (v1375 & ~i31),
  v1375 = (v617 & i32) | (v1376 & ~i32),
  v1376 = (v893 & i33) | (v1372 & ~i33),
  v1377 = (v1378 & i21) | (v617 & ~i21),
  v1378 = (v1379 & i22) | (v617 & ~i22),
  v1379 = (v1389 & i25) | (v1380 & ~i25),
  v1380 = (v1385 & i29) | (v1381 & ~i29),
  v1381 = (v617 & i30) | (v1382 & ~i30),
  v1382 = (v617 & i31) | (v1383 & ~i31),
  v1383 = (v617 & i32) | (v1384 & ~i32),
  v1384 = v903 & i34,
  v1385 = (v617 & i30) | (v1386 & ~i30),
  v1386 = (v617 & i31) | (v1387 & ~i31),
  v1387 = (v617 & i32) | (v1388 & ~i32),
  v1388 = (v617 & i33) | (v1384 & ~i33),
  v1389 = (v1394 & i29) | (v1390 & ~i29),
  v1390 = (v617 & i30) | (v1391 & ~i30),
  v1391 = (v617 & i31) | (v1392 & ~i31),
  v1392 = (v617 & i32) | (v1393 & ~i32),
  v1393 = (~v903 & ~i34) | (v903 & i34),
  v1394 = (v617 & i30) | (v1395 & ~i30),
  v1395 = (v617 & i31) | (v1396 & ~i31),
  v1396 = (v617 & i32) | (v1397 & ~i32),
  v1397 = (v902 & i33) | (v1393 & ~i33),
  v1398 = (v1442 & i19) | (v1399 & ~i19),
  v1399 = (v1421 & i20) | (v1400 & ~i20),
  v1400 = (v1401 & i21) | (v617 & ~i21),
  v1401 = (v1402 & i22) | (v617 & ~i22),
  v1402 = (v1412 & i25) | (v1403 & ~i25),
  v1403 = (v1408 & i29) | (v1404 & ~i29),
  v1404 = (v617 & i30) | (v1405 & ~i30),
  v1405 = (v617 & i31) | (v1406 & ~i31),
  v1406 = (v617 & i32) | (v1407 & ~i32),
  v1407 = v914 & i34,
  v1408 = (v617 & i30) | (v1409 & ~i30),
  v1409 = (v617 & i31) | (v1410 & ~i31),
  v1410 = (v617 & i32) | (v1411 & ~i32),
  v1411 = (v617 & i33) | (v1407 & ~i33),
  v1412 = (v1417 & i29) | (v1413 & ~i29),
  v1413 = (v617 & i30) | (v1414 & ~i30),
  v1414 = (v617 & i31) | (v1415 & ~i31),
  v1415 = (v617 & i32) | (v1416 & ~i32),
  v1416 = (~v914 & ~i34) | (v914 & i34),
  v1417 = (v617 & i30) | (v1418 & ~i30),
  v1418 = (v617 & i31) | (v1419 & ~i31),
  v1419 = (v617 & i32) | (v1420 & ~i32),
  v1420 = (v913 & i33) | (v1416 & ~i33),
  v1421 = (v1422 & i21) | (v617 & ~i21),
  v1422 = (v1423 & i22) | (v617 & ~i22),
  v1423 = (v1433 & i25) | (v1424 & ~i25),
  v1424 = (v1429 & i29) | (v1425 & ~i29),
  v1425 = (v617 & i30) | (v1426 & ~i30),
  v1426 = (v617 & i31) | (v1427 & ~i31),
  v1427 = (v617 & i32) | (v1428 & ~i32),
  v1428 = v923 & i34,
  v1429 = (v617 & i30) | (v1430 & ~i30),
  v1430 = (v617 & i31) | (v1431 & ~i31),
  v1431 = (v617 & i32) | (v1432 & ~i32),
  v1432 = (v617 & i33) | (v1428 & ~i33),
  v1433 = (v1438 & i29) | (v1434 & ~i29),
  v1434 = (v617 & i30) | (v1435 & ~i30),
  v1435 = (v617 & i31) | (v1436 & ~i31),
  v1436 = (v617 & i32) | (v1437 & ~i32),
  v1437 = (~v923 & ~i34) | (v923 & i34),
  v1438 = (v617 & i30) | (v1439 & ~i30),
  v1439 = (v617 & i31) | (v1440 & ~i31),
  v1440 = (v617 & i32) | (v1441 & ~i32),
  v1441 = (v922 & i33) | (v1437 & ~i33),
  v1442 = (v1443 & i21) | (v617 & ~i21),
  v1443 = (v1444 & i22) | (v617 & ~i22),
  v1444 = (v1454 & i25) | (v1445 & ~i25),
  v1445 = (v1450 & i29) | (v1446 & ~i29),
  v1446 = (v617 & i30) | (v1447 & ~i30),
  v1447 = (v617 & i31) | (v1448 & ~i31),
  v1448 = (v617 & i32) | (v1449 & ~i32),
  v1449 = v740 & i34,
  v1450 = (v617 & i30) | (v1451 & ~i30),
  v1451 = (v617 & i31) | (v1452 & ~i31),
  v1452 = (v617 & i32) | (v1453 & ~i32),
  v1453 = (v617 & i33) | (v1449 & ~i33),
  v1454 = (v1459 & i29) | (v1455 & ~i29),
  v1455 = (v617 & i30) | (v1456 & ~i30),
  v1456 = (v617 & i31) | (v1457 & ~i31),
  v1457 = (v617 & i32) | (v1458 & ~i32),
  v1458 = (~v740 & ~i34) | (v740 & i34),
  v1459 = (v617 & i30) | (v1460 & ~i30),
  v1460 = (v617 & i31) | (v1461 & ~i31),
  v1461 = (v617 & i32) | (v1462 & ~i32),
  v1462 = (v931 & i33) | (v1458 & ~i33),
  v1463 = (v1551 & i17) | (v1464 & ~i17),
  v1464 = (v1508 & i19) | (v1465 & ~i19),
  v1465 = (v1487 & i20) | (v1466 & ~i20),
  v1466 = (v1467 & i21) | (v617 & ~i21),
  v1467 = (v1468 & i22) | (v617 & ~i22),
  v1468 = (v1478 & i25) | (v1469 & ~i25),
  v1469 = (v1474 & i29) | (v1470 & ~i29),
  v1470 = (v617 & i30) | (v1471 & ~i30),
  v1471 = (v617 & i31) | (v1472 & ~i31),
  v1472 = (v617 & i32) | (v1473 & ~i32),
  v1473 = v942 & i34,
  v1474 = (v617 & i30) | (v1475 & ~i30),
  v1475 = (v617 & i31) | (v1476 & ~i31),
  v1476 = (v617 & i32) | (v1477 & ~i32),
  v1477 = (v617 & i33) | (v1473 & ~i33),
  v1478 = (v1483 & i29) | (v1479 & ~i29),
  v1479 = (v617 & i30) | (v1480 & ~i30),
  v1480 = (v617 & i31) | (v1481 & ~i31),
  v1481 = (v617 & i32) | (v1482 & ~i32),
  v1482 = (~v942 & ~i34) | (v942 & i34),
  v1483 = (v617 & i30) | (v1484 & ~i30),
  v1484 = (v617 & i31) | (v1485 & ~i31),
  v1485 = (v617 & i32) | (v1486 & ~i32),
  v1486 = (v941 & i33) | (v1482 & ~i33),
  v1487 = (v1488 & i21) | (v617 & ~i21),
  v1488 = (v1489 & i22) | (v617 & ~i22),
  v1489 = (v1499 & i25) | (v1490 & ~i25),
  v1490 = (v1495 & i29) | (v1491 & ~i29),
  v1491 = (v617 & i30) | (v1492 & ~i30),
  v1492 = (v617 & i31) | (v1493 & ~i31),
  v1493 = (v617 & i32) | (v1494 & ~i32),
  v1494 = v952 & i34,
  v1495 = (v617 & i30) | (v1496 & ~i30),
  v1496 = (v617 & i31) | (v1497 & ~i31),
  v1497 = (v617 & i32) | (v1498 & ~i32),
  v1498 = (v617 & i33) | (v1494 & ~i33),
  v1499 = (v1504 & i29) | (v1500 & ~i29),
  v1500 = (v617 & i30) | (v1501 & ~i30),
  v1501 = (v617 & i31) | (v1502 & ~i31),
  v1502 = (v617 & i32) | (v1503 & ~i32),
  v1503 = (~v952 & ~i34) | (v952 & i34),
  v1504 = (v617 & i30) | (v1505 & ~i30),
  v1505 = (v617 & i31) | (v1506 & ~i31),
  v1506 = (v617 & i32) | (v1507 & ~i32),
  v1507 = (v951 & i33) | (v1503 & ~i33),
  v1508 = (v1530 & i20) | (v1509 & ~i20),
  v1509 = (v1510 & i21) | (v617 & ~i21),
  v1510 = (v1511 & i22) | (v617 & ~i22),
  v1511 = (v1521 & i25) | (v1512 & ~i25),
  v1512 = (v1517 & i29) | (v1513 & ~i29),
  v1513 = (v617 & i30) | (v1514 & ~i30),
  v1514 = (v617 & i31) | (v1515 & ~i31),
  v1515 = (v617 & i32) | (v1516 & ~i32),
  v1516 = v963 & i34,
  v1517 = (v617 & i30) | (v1518 & ~i30),
  v1518 = (v617 & i31) | (v1519 & ~i31),
  v1519 = (v617 & i32) | (v1520 & ~i32),
  v1520 = (v617 & i33) | (v1516 & ~i33),
  v1521 = (v1526 & i29) | (v1522 & ~i29),
  v1522 = (v617 & i30) | (v1523 & ~i30),
  v1523 = (v617 & i31) | (v1524 & ~i31),
  v1524 = (v617 & i32) | (v1525 & ~i32),
  v1525 = (~v963 & ~i34) | (v963 & i34),
  v1526 = (v617 & i30) | (v1527 & ~i30),
  v1527 = (v617 & i31) | (v1528 & ~i31),
  v1528 = (v617 & i32) | (v1529 & ~i32),
  v1529 = (v962 & i33) | (v1525 & ~i33),
  v1530 = (v1531 & i21) | (v617 & ~i21),
  v1531 = (v1532 & i22) | (v617 & ~i22),
  v1532 = (v1542 & i25) | (v1533 & ~i25),
  v1533 = (v1538 & i29) | (v1534 & ~i29),
  v1534 = (v617 & i30) | (v1535 & ~i30),
  v1535 = (v617 & i31) | (v1536 & ~i31),
  v1536 = (v617 & i32) | (v1537 & ~i32),
  v1537 = v972 & i34,
  v1538 = (v617 & i30) | (v1539 & ~i30),
  v1539 = (v617 & i31) | (v1540 & ~i31),
  v1540 = (v617 & i32) | (v1541 & ~i32),
  v1541 = (v617 & i33) | (v1537 & ~i33),
  v1542 = (v1547 & i29) | (v1543 & ~i29),
  v1543 = (v617 & i30) | (v1544 & ~i30),
  v1544 = (v617 & i31) | (v1545 & ~i31),
  v1545 = (v617 & i32) | (v1546 & ~i32),
  v1546 = (~v972 & ~i34) | (v972 & i34),
  v1547 = (v617 & i30) | (v1548 & ~i30),
  v1548 = (v617 & i31) | (v1549 & ~i31),
  v1549 = (v617 & i32) | (v1550 & ~i32),
  v1550 = (v971 & i33) | (v1546 & ~i33),
  v1551 = (v1595 & i19) | (v1552 & ~i19),
  v1552 = (v1574 & i20) | (v1553 & ~i20),
  v1553 = (v1554 & i21) | (v617 & ~i21),
  v1554 = (v1555 & i22) | (v617 & ~i22),
  v1555 = (v1565 & i25) | (v1556 & ~i25),
  v1556 = (v1561 & i29) | (v1557 & ~i29),
  v1557 = (v617 & i30) | (v1558 & ~i30),
  v1558 = (v617 & i31) | (v1559 & ~i31),
  v1559 = (v617 & i32) | (v1560 & ~i32),
  v1560 = v983 & i34,
  v1561 = (v617 & i30) | (v1562 & ~i30),
  v1562 = (v617 & i31) | (v1563 & ~i31),
  v1563 = (v617 & i32) | (v1564 & ~i32),
  v1564 = (v617 & i33) | (v1560 & ~i33),
  v1565 = (v1570 & i29) | (v1566 & ~i29),
  v1566 = (v617 & i30) | (v1567 & ~i30),
  v1567 = (v617 & i31) | (v1568 & ~i31),
  v1568 = (v617 & i32) | (v1569 & ~i32),
  v1569 = (~v983 & ~i34) | (v983 & i34),
  v1570 = (v617 & i30) | (v1571 & ~i30),
  v1571 = (v617 & i31) | (v1572 & ~i31),
  v1572 = (v617 & i32) | (v1573 & ~i32),
  v1573 = (v982 & i33) | (v1569 & ~i33),
  v1574 = (v1575 & i21) | (v617 & ~i21),
  v1575 = (v1576 & i22) | (v617 & ~i22),
  v1576 = (v1586 & i25) | (v1577 & ~i25),
  v1577 = (v1582 & i29) | (v1578 & ~i29),
  v1578 = (v617 & i30) | (v1579 & ~i30),
  v1579 = (v617 & i31) | (v1580 & ~i31),
  v1580 = (v617 & i32) | (v1581 & ~i32),
  v1581 = v992 & i34,
  v1582 = (v617 & i30) | (v1583 & ~i30),
  v1583 = (v617 & i31) | (v1584 & ~i31),
  v1584 = (v617 & i32) | (v1585 & ~i32),
  v1585 = (v617 & i33) | (v1581 & ~i33),
  v1586 = (v1591 & i29) | (v1587 & ~i29),
  v1587 = (v617 & i30) | (v1588 & ~i30),
  v1588 = (v617 & i31) | (v1589 & ~i31),
  v1589 = (v617 & i32) | (v1590 & ~i32),
  v1590 = (~v992 & ~i34) | (v992 & i34),
  v1591 = (v617 & i30) | (v1592 & ~i30),
  v1592 = (v617 & i31) | (v1593 & ~i31),
  v1593 = (v617 & i32) | (v1594 & ~i32),
  v1594 = (v991 & i33) | (v1590 & ~i33),
  v1595 = (v1596 & i21) | (v617 & ~i21),
  v1596 = (v1597 & i22) | (v617 & ~i22),
  v1597 = (v1607 & i25) | (v1598 & ~i25),
  v1598 = (v1603 & i29) | (v1599 & ~i29),
  v1599 = (v617 & i30) | (v1600 & ~i30),
  v1600 = (v617 & i31) | (v1601 & ~i31),
  v1601 = (v617 & i32) | (v1602 & ~i32),
  v1602 = v858 & i34,
  v1603 = (v617 & i30) | (v1604 & ~i30),
  v1604 = (v617 & i31) | (v1605 & ~i31),
  v1605 = (v617 & i32) | (v1606 & ~i32),
  v1606 = (v617 & i33) | (v1602 & ~i33),
  v1607 = (v1612 & i29) | (v1608 & ~i29),
  v1608 = (v617 & i30) | (v1609 & ~i30),
  v1609 = (v617 & i31) | (v1610 & ~i31),
  v1610 = (v617 & i32) | (v1611 & ~i32),
  v1611 = (~v858 & ~i34) | (v858 & i34),
  v1612 = (v617 & i30) | (v1613 & ~i30),
  v1613 = (v617 & i31) | (v1614 & ~i31),
  v1614 = (v617 & i32) | (v1615 & ~i32),
  v1615 = (v1000 & i33) | (v1611 & ~i33),
  v1616 = (v1620 & i11) | (v1617 & ~i11),
  v1617 = (v1620 & i12) | (v1618 & ~i12),
  v1618 = (v1620 & i13) | (v1619 & ~i13),
  v1619 = (v1843 & i14) | (v1620 & ~i14),
  v1620 = (v1732 & i15) | (v1621 & ~i15),
  v1621 = (v1677 & i16) | (v1622 & ~i16),
  v1622 = (v1654 & i17) | (v1623 & ~i17),
  v1623 = (v1639 & i19) | (v1624 & ~i19),
  v1624 = (v1632 & i20) | (v1625 & ~i20),
  v1625 = (v1626 & i21) | (v617 & ~i21),
  v1626 = (v1627 & i22) | (v617 & ~i22),
  v1627 = (v1628 & i29) | (v620 & ~i29),
  v1628 = (v617 & i30) | (v1629 & ~i30),
  v1629 = (v617 & i31) | (v1630 & ~i31),
  v1630 = (v617 & i32) | (v1631 & ~i32),
  v1631 = (v623 & i33) | (v617 & ~i33),
  v1632 = (v1633 & i21) | (v617 & ~i21),
  v1633 = (v1634 & i22) | (v617 & ~i22),
  v1634 = (v1635 & i29) | (v640 & ~i29),
  v1635 = (v617 & i30) | (v1636 & ~i30),
  v1636 = (v617 & i31) | (v1637 & ~i31),
  v1637 = (v617 & i32) | (v1638 & ~i32),
  v1638 = (v643 & i33) | (v617 & ~i33),
  v1639 = (v1647 & i20) | (v1640 & ~i20),
  v1640 = (v1641 & i21) | (v617 & ~i21),
  v1641 = (v1642 & i22) | (v617 & ~i22),
  v1642 = (v1643 & i29) | (v658 & ~i29),
  v1643 = (v617 & i30) | (v1644 & ~i30),
  v1644 = (v617 & i31) | (v1645 & ~i31),
  v1645 = (v617 & i32) | (v1646 & ~i32),
  v1646 = (v661 & i33) | (v617 & ~i33),
  v1647 = (v1648 & i21) | (v617 & ~i21),
  v1648 = (v1649 & i22) | (v617 & ~i22),
  v1649 = (v1650 & i29) | (v679 & ~i29),
  v1650 = (v617 & i30) | (v1651 & ~i30),
  v1651 = (v617 & i31) | (v1652 & ~i31),
  v1652 = (v617 & i32) | (v1653 & ~i32),
  v1653 = (v682 & i33) | (v617 & ~i33),
  v1654 = (v1670 & i19) | (v1655 & ~i19),
  v1655 = (v1663 & i20) | (v1656 & ~i20),
  v1656 = (v1657 & i21) | (v617 & ~i21),
  v1657 = (v1658 & i22) | (v617 & ~i22),
  v1658 = (v1659 & i29) | (v699 & ~i29),
  v1659 = (v617 & i30) | (v1660 & ~i30),
  v1660 = (v617 & i31) | (v1661 & ~i31),
  v1661 = (v617 & i32) | (v1662 & ~i32),
  v1662 = (v702 & i33) | (v617 & ~i33),
  v1663 = (v1664 & i21) | (v617 & ~i21),
  v1664 = (v1665 & i22) | (v617 & ~i22),
  v1665 = (v1666 & i29) | (v717 & ~i29),
  v1666 = (v617 & i30) | (v1667 & ~i30),
  v1667 = (v617 & i31) | (v1668 & ~i31),
  v1668 = (v617 & i32) | (v1669 & ~i32),
  v1669 = (v720 & i33) | (v617 & ~i33),
  v1670 = (v1671 & i21) | (v617 & ~i21),
  v1671 = (v1672 & i22) | (v617 & ~i22),
  v1672 = (v1673 & i29) | (v735 & ~i29),
  v1673 = (v617 & i30) | (v1674 & ~i30),
  v1674 = (v617 & i31) | (v1675 & ~i31),
  v1675 = (v617 & i32) | (v1676 & ~i32),
  v1676 = (v738 & i33) | (v617 & ~i33),
  v1677 = (v1709 & i17) | (v1678 & ~i17),
  v1678 = (v1694 & i19) | (v1679 & ~i19),
  v1679 = (v1687 & i20) | (v1680 & ~i20),
  v1680 = (v1681 & i21) | (v617 & ~i21),
  v1681 = (v1682 & i22) | (v617 & ~i22),
  v1682 = (v1683 & i29) | (v750 & ~i29),
  v1683 = (v617 & i30) | (v1684 & ~i30),
  v1684 = (v617 & i31) | (v1685 & ~i31),
  v1685 = (v617 & i32) | (v1686 & ~i32),
  v1686 = (v753 & i33) | (v617 & ~i33),
  v1687 = (v1688 & i21) | (v617 & ~i21),
  v1688 = (v1689 & i22) | (v617 & ~i22),
  v1689 = (v1690 & i29) | (v764 & ~i29),
  v1690 = (v617 & i30) | (v1691 & ~i30),
  v1691 = (v617 & i31) | (v1692 & ~i31),
  v1692 = (v617 & i32) | (v1693 & ~i32),
  v1693 = (v767 & i33) | (v617 & ~i33),
  v1694 = (v1702 & i20) | (v1695 & ~i20),
  v1695 = (v1696 & i21) | (v617 & ~i21),
  v1696 = (v1697 & i22) | (v617 & ~i22),
  v1697 = (v1698 & i29) | (v779 & ~i29),
  v1698 = (v617 & i30) | (v1699 & ~i30),
  v1699 = (v617 & i31) | (v1700 & ~i31),
  v1700 = (v617 & i32) | (v1701 & ~i32),
  v1701 = (v782 & i33) | (v617 & ~i33),
  v1702 = (v1703 & i21) | (v617 & ~i21),
  v1703 = (v1704 & i22) | (v617 & ~i22),
  v1704 = (v1705 & i29) | (v797 & ~i29),
  v1705 = (v617 & i30) | (v1706 & ~i30),
  v1706 = (v617 & i31) | (v1707 & ~i31),
  v1707 = (v617 & i32) | (v1708 & ~i32),
  v1708 = (v800 & i33) | (v617 & ~i33),
  v1709 = (v1725 & i19) | (v1710 & ~i19),
  \*clm_file_1_istate0  = ~v152,
  \*clm_file_1_istate1  = ~v64,
  v1710 = (v1718 & i20) | (v1711 & ~i20),
  v1711 = (v1712 & i21) | (v617 & ~i21),
  v1712 = (v1713 & i22) | (v617 & ~i22),
  v1713 = (v1714 & i29) | (v817 & ~i29),
  v1714 = (v617 & i30) | (v1715 & ~i30),
  v1715 = (v617 & i31) | (v1716 & ~i31),
  v1716 = (v617 & i32) | (v1717 & ~i32),
  v1717 = (v820 & i33) | (v617 & ~i33),
  v1718 = (v1719 & i21) | (v617 & ~i21),
  v1719 = (v1720 & i22) | (v617 & ~i22),
  v1720 = (v1721 & i29) | (v835 & ~i29),
  v1721 = (v617 & i30) | (v1722 & ~i30),
  v1722 = (v617 & i31) | (v1723 & ~i31),
  v1723 = (v617 & i32) | (v1724 & ~i32),
  v1724 = (v838 & i33) | (v617 & ~i33),
  v1725 = (v1726 & i21) | (v617 & ~i21),
  v1726 = (v1727 & i22) | (v617 & ~i22),
  v1727 = (v1728 & i29) | (v853 & ~i29),
  v1728 = (v617 & i30) | (v1729 & ~i30),
  v1729 = (v617 & i31) | (v1730 & ~i31),
  v1730 = (v617 & i32) | (v1731 & ~i32),
  v1731 = (v856 & i33) | (v617 & ~i33),
  v1732 = (v1788 & i16) | (v1733 & ~i16),
  v1733 = (v1765 & i17) | (v1734 & ~i17),
  v1734 = (v1750 & i19) | (v1735 & ~i19),
  v1735 = (v1743 & i20) | (v1736 & ~i20),
  v1736 = (v1737 & i21) | (v617 & ~i21),
  v1737 = (v1738 & i22) | (v617 & ~i22),
  v1738 = (v1739 & i29) | (v869 & ~i29),
  v1739 = (v617 & i30) | (v1740 & ~i30),
  v1740 = (v617 & i31) | (v1741 & ~i31),
  v1741 = (v617 & i32) | (v1742 & ~i32),
  v1742 = (v872 & i33) | (v617 & ~i33),
  v1743 = (v1744 & i21) | (v617 & ~i21),
  v1744 = (v1745 & i22) | (v617 & ~i22),
  v1745 = (v1746 & i29) | (v879 & ~i29),
  v1746 = (v617 & i30) | (v1747 & ~i30),
  v1747 = (v617 & i31) | (v1748 & ~i31),
  v1748 = (v617 & i32) | (v1749 & ~i32),
  v1749 = (v882 & i33) | (v617 & ~i33),
  v1750 = (v1758 & i20) | (v1751 & ~i20),
  v1751 = (v1752 & i21) | (v617 & ~i21),
  v1752 = (v1753 & i22) | (v617 & ~i22),
  v1753 = (v1754 & i29) | (v890 & ~i29),
  v1754 = (v617 & i30) | (v1755 & ~i30),
  v1755 = (v617 & i31) | (v1756 & ~i31),
  v1756 = (v617 & i32) | (v1757 & ~i32),
  v1757 = (v893 & i33) | (v617 & ~i33),
  v1758 = (v1759 & i21) | (v617 & ~i21),
  v1759 = (v1760 & i22) | (v617 & ~i22),
  v1760 = (v1761 & i29) | (v899 & ~i29),
  v1761 = (v617 & i30) | (v1762 & ~i30),
  v1762 = (v617 & i31) | (v1763 & ~i31),
  v1763 = (v617 & i32) | (v1764 & ~i32),
  v1764 = (v902 & i33) | (v617 & ~i33),
  v1765 = (v1781 & i19) | (v1766 & ~i19),
  v1766 = (v1774 & i20) | (v1767 & ~i20),
  v1767 = (v1768 & i21) | (v617 & ~i21),
  v1768 = (v1769 & i22) | (v617 & ~i22),
  v1769 = (v1770 & i29) | (v910 & ~i29),
  v1770 = (v617 & i30) | (v1771 & ~i30),
  v1771 = (v617 & i31) | (v1772 & ~i31),
  v1772 = (v617 & i32) | (v1773 & ~i32),
  v1773 = (v913 & i33) | (v617 & ~i33),
  v1774 = (v1775 & i21) | (v617 & ~i21),
  v1775 = (v1776 & i22) | (v617 & ~i22),
  v1776 = (v1777 & i29) | (v919 & ~i29),
  v1777 = (v617 & i30) | (v1778 & ~i30),
  v1778 = (v617 & i31) | (v1779 & ~i31),
  v1779 = (v617 & i32) | (v1780 & ~i32),
  v1780 = (v922 & i33) | (v617 & ~i33),
  v1781 = (v1782 & i21) | (v617 & ~i21),
  v1782 = (v1783 & i22) | (v617 & ~i22),
  v1783 = (v1784 & i29) | (v928 & ~i29),
  v1784 = (v617 & i30) | (v1785 & ~i30),
  v1785 = (v617 & i31) | (v1786 & ~i31),
  v1786 = (v617 & i32) | (v1787 & ~i32),
  v1787 = (v931 & i33) | (v617 & ~i33),
  v1788 = (v1820 & i17) | (v1789 & ~i17),
  v1789 = (v1805 & i19) | (v1790 & ~i19),
  v1790 = (v1798 & i20) | (v1791 & ~i20),
  v1791 = (v1792 & i21) | (v617 & ~i21),
  v1792 = (v1793 & i22) | (v617 & ~i22),
  v1793 = (v1794 & i29) | (v938 & ~i29),
  v1794 = (v617 & i30) | (v1795 & ~i30),
  v1795 = (v617 & i31) | (v1796 & ~i31),
  v1796 = (v617 & i32) | (v1797 & ~i32),
  v1797 = (v941 & i33) | (v617 & ~i33),
  v1798 = (v1799 & i21) | (v617 & ~i21),
  v1799 = (v1800 & i22) | (v617 & ~i22),
  v1800 = (v1801 & i29) | (v948 & ~i29),
  v1801 = (v617 & i30) | (v1802 & ~i30),
  v1802 = (v617 & i31) | (v1803 & ~i31),
  v1803 = (v617 & i32) | (v1804 & ~i32),
  v1804 = (v951 & i33) | (v617 & ~i33),
  v1805 = (v1813 & i20) | (v1806 & ~i20),
  v1806 = (v1807 & i21) | (v617 & ~i21),
  v1807 = (v1808 & i22) | (v617 & ~i22),
  v1808 = (v1809 & i29) | (v959 & ~i29),
  v1809 = (v617 & i30) | (v1810 & ~i30),
  v1810 = (v617 & i31) | (v1811 & ~i31),
  v1811 = (v617 & i32) | (v1812 & ~i32),
  v1812 = (v962 & i33) | (v617 & ~i33),
  v1813 = (v1814 & i21) | (v617 & ~i21),
  v1814 = (v1815 & i22) | (v617 & ~i22),
  v1815 = (v1816 & i29) | (v968 & ~i29),
  v1816 = (v617 & i30) | (v1817 & ~i30),
  v1817 = (v617 & i31) | (v1818 & ~i31),
  v1818 = (v617 & i32) | (v1819 & ~i32),
  v1819 = (v971 & i33) | (v617 & ~i33),
  v1820 = (v1836 & i19) | (v1821 & ~i19),
  v1821 = (v1829 & i20) | (v1822 & ~i20),
  v1822 = (v1823 & i21) | (v617 & ~i21),
  v1823 = (v1824 & i22) | (v617 & ~i22),
  v1824 = (v1825 & i29) | (v979 & ~i29),
  v1825 = (v617 & i30) | (v1826 & ~i30),
  v1826 = (v617 & i31) | (v1827 & ~i31),
  v1827 = (v617 & i32) | (v1828 & ~i32),
  v1828 = (v982 & i33) | (v617 & ~i33),
  v1829 = (v1830 & i21) | (v617 & ~i21),
  v1830 = (v1831 & i22) | (v617 & ~i22),
  v1831 = (v1832 & i29) | (v988 & ~i29),
  v1832 = (v617 & i30) | (v1833 & ~i30),
  v1833 = (v617 & i31) | (v1834 & ~i31),
  v1834 = (v617 & i32) | (v1835 & ~i32),
  v1835 = (v991 & i33) | (v617 & ~i33),
  v1836 = (v1837 & i21) | (v617 & ~i21),
  v1837 = (v1838 & i22) | (v617 & ~i22),
  v1838 = (v1839 & i29) | (v997 & ~i29),
  v1839 = (v617 & i30) | (v1840 & ~i30),
  v1840 = (v617 & i31) | (v1841 & ~i31),
  v1841 = (v617 & i32) | (v1842 & ~i32),
  v1842 = (v1000 & i33) | (v617 & ~i33),
  v1843 = (v1955 & i15) | (v1844 & ~i15),
  v1844 = (v1900 & i16) | (v1845 & ~i16),
  v1845 = (v1877 & i17) | (v1846 & ~i17),
  v1846 = (v1862 & i19) | (v1847 & ~i19),
  v1847 = (v1855 & i20) | (v1848 & ~i20),
  v1848 = (v1849 & i21) | (v617 & ~i21),
  v1849 = (v1850 & i22) | (v617 & ~i22),
  v1850 = (v1851 & i29) | (v1019 & ~i29),
  v1851 = (v617 & i30) | (v1852 & ~i30),
  v1852 = (v617 & i31) | (v1853 & ~i31),
  v1853 = (v617 & i32) | (v1854 & ~i32),
  v1854 = (v623 & i33) | (v1013 & ~i33),
  v1855 = (v1856 & i21) | (v617 & ~i21),
  v1856 = (v1857 & i22) | (v617 & ~i22),
  v1857 = (v1858 & i29) | (v1040 & ~i29),
  v1858 = (v617 & i30) | (v1859 & ~i30),
  v1859 = (v617 & i31) | (v1860 & ~i31),
  v1860 = (v617 & i32) | (v1861 & ~i32),
  v1861 = (v643 & i33) | (v1034 & ~i33),
  v1862 = (v1870 & i20) | (v1863 & ~i20),
  v1863 = (v1864 & i21) | (v617 & ~i21),
  v1864 = (v1865 & i22) | (v617 & ~i22),
  v1865 = (v1866 & i29) | (v1062 & ~i29),
  v1866 = (v617 & i30) | (v1867 & ~i30),
  v1867 = (v617 & i31) | (v1868 & ~i31),
  v1868 = (v617 & i32) | (v1869 & ~i32),
  v1869 = (v661 & i33) | (v1056 & ~i33),
  v1870 = (v1871 & i21) | (v617 & ~i21),
  v1871 = (v1872 & i22) | (v617 & ~i22),
  v1872 = (v1873 & i29) | (v1083 & ~i29),
  v1873 = (v617 & i30) | (v1874 & ~i30),
  v1874 = (v617 & i31) | (v1875 & ~i31),
  v1875 = (v617 & i32) | (v1876 & ~i32),
  v1876 = (v682 & i33) | (v1077 & ~i33),
  v1877 = (v1893 & i19) | (v1878 & ~i19),
  v1878 = (v1886 & i20) | (v1879 & ~i20),
  v1879 = (v1880 & i21) | (v617 & ~i21),
  v1880 = (v1881 & i22) | (v617 & ~i22),
  v1881 = (v1882 & i29) | (v1106 & ~i29),
  v1882 = (v617 & i30) | (v1883 & ~i30),
  v1883 = (v617 & i31) | (v1884 & ~i31),
  v1884 = (v617 & i32) | (v1885 & ~i32),
  v1885 = (v702 & i33) | (v1100 & ~i33),
  v1886 = (v1887 & i21) | (v617 & ~i21),
  v1887 = (v1888 & i22) | (v617 & ~i22),
  v1888 = (v1889 & i29) | (v1127 & ~i29),
  v1889 = (v617 & i30) | (v1890 & ~i30),
  v1890 = (v617 & i31) | (v1891 & ~i31),
  v1891 = (v617 & i32) | (v1892 & ~i32),
  v1892 = (v720 & i33) | (v1121 & ~i33),
  v1893 = (v1894 & i21) | (v617 & ~i21),
  v1894 = (v1895 & i22) | (v617 & ~i22),
  v1895 = (v1896 & i29) | (v1148 & ~i29),
  v1896 = (v617 & i30) | (v1897 & ~i30),
  v1897 = (v617 & i31) | (v1898 & ~i31),
  v1898 = (v617 & i32) | (v1899 & ~i32),
  v1899 = (v738 & i33) | (v1142 & ~i33),
  v1900 = (v1932 & i17) | (v1901 & ~i17),
  v1901 = (v1917 & i19) | (v1902 & ~i19),
  v1902 = (v1910 & i20) | (v1903 & ~i20),
  v1903 = (v1904 & i21) | (v617 & ~i21),
  v1904 = (v1905 & i22) | (v617 & ~i22),
  v1905 = (v1906 & i29) | (v1172 & ~i29),
  v1906 = (v617 & i30) | (v1907 & ~i30),
  v1907 = (v617 & i31) | (v1908 & ~i31),
  v1908 = (v617 & i32) | (v1909 & ~i32),
  v1909 = (v753 & i33) | (v1166 & ~i33),
  v1910 = (v1911 & i21) | (v617 & ~i21),
  v1911 = (v1912 & i22) | (v617 & ~i22),
  v1912 = (v1913 & i29) | (v1193 & ~i29),
  v1913 = (v617 & i30) | (v1914 & ~i30),
  v1914 = (v617 & i31) | (v1915 & ~i31),
  v1915 = (v617 & i32) | (v1916 & ~i32),
  v1916 = (v767 & i33) | (v1187 & ~i33),
  v1917 = (v1925 & i20) | (v1918 & ~i20),
  v1918 = (v1919 & i21) | (v617 & ~i21),
  v1919 = (v1920 & i22) | (v617 & ~i22),
  v1920 = (v1921 & i29) | (v1215 & ~i29),
  v1921 = (v617 & i30) | (v1922 & ~i30),
  v1922 = (v617 & i31) | (v1923 & ~i31),
  v1923 = (v617 & i32) | (v1924 & ~i32),
  v1924 = (v782 & i33) | (v1209 & ~i33),
  v1925 = (v1926 & i21) | (v617 & ~i21),
  v1926 = (v1927 & i22) | (v617 & ~i22),
  v1927 = (v1928 & i29) | (v1236 & ~i29),
  v1928 = (v617 & i30) | (v1929 & ~i30),
  v1929 = (v617 & i31) | (v1930 & ~i31),
  v1930 = (v617 & i32) | (v1931 & ~i32),
  v1931 = (v800 & i33) | (v1230 & ~i33),
  v1932 = (v1948 & i19) | (v1933 & ~i19),
  v1933 = (v1941 & i20) | (v1934 & ~i20),
  v1934 = (v1935 & i21) | (v617 & ~i21),
  v1935 = (v1936 & i22) | (v617 & ~i22),
  v1936 = (v1937 & i29) | (v1259 & ~i29),
  v1937 = (v617 & i30) | (v1938 & ~i30),
  v1938 = (v617 & i31) | (v1939 & ~i31),
  v1939 = (v617 & i32) | (v1940 & ~i32),
  v1940 = (v820 & i33) | (v1253 & ~i33),
  v1941 = (v1942 & i21) | (v617 & ~i21),
  v1942 = (v1943 & i22) | (v617 & ~i22),
  v1943 = (v1944 & i29) | (v1280 & ~i29),
  v1944 = (v617 & i30) | (v1945 & ~i30),
  v1945 = (v617 & i31) | (v1946 & ~i31),
  v1946 = (v617 & i32) | (v1947 & ~i32),
  v1947 = (v838 & i33) | (v1274 & ~i33),
  v1948 = (v1949 & i21) | (v617 & ~i21),
  v1949 = (v1950 & i22) | (v617 & ~i22),
  v1950 = (v1951 & i29) | (v1301 & ~i29),
  v1951 = (v617 & i30) | (v1952 & ~i30),
  v1952 = (v617 & i31) | (v1953 & ~i31),
  v1953 = (v617 & i32) | (v1954 & ~i32),
  v1954 = (v856 & i33) | (v1295 & ~i33),
  v1955 = (v2011 & i16) | (v1956 & ~i16),
  v1956 = (v1988 & i17) | (v1957 & ~i17),
  v1957 = (v1973 & i19) | (v1958 & ~i19),
  v1958 = (v1966 & i20) | (v1959 & ~i20),
  v1959 = (v1960 & i21) | (v617 & ~i21),
  v1960 = (v1961 & i22) | (v617 & ~i22),
  v1961 = (v1962 & i29) | (v1326 & ~i29),
  v1962 = (v617 & i30) | (v1963 & ~i30),
  v1963 = (v617 & i31) | (v1964 & ~i31),
  v1964 = (v617 & i32) | (v1965 & ~i32),
  v1965 = (v872 & i33) | (v1320 & ~i33),
  v1966 = (v1967 & i21) | (v617 & ~i21),
  v1967 = (v1968 & i22) | (v617 & ~i22),
  v1968 = (v1969 & i29) | (v1347 & ~i29),
  v1969 = (v617 & i30) | (v1970 & ~i30),
  v1970 = (v617 & i31) | (v1971 & ~i31),
  v1971 = (v617 & i32) | (v1972 & ~i32),
  v1972 = (v882 & i33) | (v1341 & ~i33),
  v1973 = (v1981 & i20) | (v1974 & ~i20),
  v1974 = (v1975 & i21) | (v617 & ~i21),
  v1975 = (v1976 & i22) | (v617 & ~i22),
  v1976 = (v1977 & i29) | (v1369 & ~i29),
  v1977 = (v617 & i30) | (v1978 & ~i30),
  v1978 = (v617 & i31) | (v1979 & ~i31),
  v1979 = (v617 & i32) | (v1980 & ~i32),
  v1980 = (v893 & i33) | (v1363 & ~i33),
  v1981 = (v1982 & i21) | (v617 & ~i21),
  v1982 = (v1983 & i22) | (v617 & ~i22),
  v1983 = (v1984 & i29) | (v1390 & ~i29),
  v1984 = (v617 & i30) | (v1985 & ~i30),
  v1985 = (v617 & i31) | (v1986 & ~i31),
  v1986 = (v617 & i32) | (v1987 & ~i32),
  v1987 = (v902 & i33) | (v1384 & ~i33),
  v1988 = (v2004 & i19) | (v1989 & ~i19),
  v1989 = (v1997 & i20) | (v1990 & ~i20),
  v1990 = (v1991 & i21) | (v617 & ~i21),
  v1991 = (v1992 & i22) | (v617 & ~i22),
  v1992 = (v1993 & i29) | (v1413 & ~i29),
  v1993 = (v617 & i30) | (v1994 & ~i30),
  v1994 = (v617 & i31) | (v1995 & ~i31),
  v1995 = (v617 & i32) | (v1996 & ~i32),
  v1996 = (v913 & i33) | (v1407 & ~i33),
  v1997 = (v1998 & i21) | (v617 & ~i21),
  v1998 = (v1999 & i22) | (v617 & ~i22),
  v1999 = (v2000 & i29) | (v1434 & ~i29),
  v2000 = (v617 & i30) | (v2001 & ~i30),
  v2001 = (v617 & i31) | (v2002 & ~i31),
  v2002 = (v617 & i32) | (v2003 & ~i32),
  v2003 = (v922 & i33) | (v1428 & ~i33),
  v2004 = (v2005 & i21) | (v617 & ~i21),
  v2005 = (v2006 & i22) | (v617 & ~i22),
  v2006 = (v2007 & i29) | (v1455 & ~i29),
  v2007 = (v617 & i30) | (v2008 & ~i30),
  v2008 = (v617 & i31) | (v2009 & ~i31),
  v2009 = (v617 & i32) | (v2010 & ~i32),
  v2010 = (v931 & i33) | (v1449 & ~i33),
  v2011 = (v2043 & i17) | (v2012 & ~i17),
  v2012 = (v2028 & i19) | (v2013 & ~i19),
  v2013 = (v2021 & i20) | (v2014 & ~i20),
  v2014 = (v2015 & i21) | (v617 & ~i21),
  v2015 = (v2016 & i22) | (v617 & ~i22),
  v2016 = (v2017 & i29) | (v1479 & ~i29),
  v2017 = (v617 & i30) | (v2018 & ~i30),
  v2018 = (v617 & i31) | (v2019 & ~i31),
  v2019 = (v617 & i32) | (v2020 & ~i32),
  v2020 = (v941 & i33) | (v1473 & ~i33),
  v2021 = (v2022 & i21) | (v617 & ~i21),
  v2022 = (v2023 & i22) | (v617 & ~i22),
  v2023 = (v2024 & i29) | (v1500 & ~i29),
  v2024 = (v617 & i30) | (v2025 & ~i30),
  v2025 = (v617 & i31) | (v2026 & ~i31),
  v2026 = (v617 & i32) | (v2027 & ~i32),
  v2027 = (v951 & i33) | (v1494 & ~i33),
  v2028 = (v2036 & i20) | (v2029 & ~i20),
  v2029 = (v2030 & i21) | (v617 & ~i21),
  v2030 = (v2031 & i22) | (v617 & ~i22),
  v2031 = (v2032 & i29) | (v1522 & ~i29),
  v2032 = (v617 & i30) | (v2033 & ~i30),
  v2033 = (v617 & i31) | (v2034 & ~i31),
  v2034 = (v617 & i32) | (v2035 & ~i32),
  v2035 = (v962 & i33) | (v1516 & ~i33),
  v2036 = (v2037 & i21) | (v617 & ~i21),
  v2037 = (v2038 & i22) | (v617 & ~i22),
  v2038 = (v2039 & i29) | (v1543 & ~i29),
  v2039 = (v617 & i30) | (v2040 & ~i30),
  v2040 = (v617 & i31) | (v2041 & ~i31),
  v2041 = (v617 & i32) | (v2042 & ~i32),
  v2042 = (v971 & i33) | (v1537 & ~i33),
  v2043 = (v2059 & i19) | (v2044 & ~i19),
  v2044 = (v2052 & i20) | (v2045 & ~i20),
  v2045 = (v2046 & i21) | (v617 & ~i21),
  v2046 = (v2047 & i22) | (v617 & ~i22),
  v2047 = (v2048 & i29) | (v1566 & ~i29),
  v2048 = (v617 & i30) | (v2049 & ~i30),
  v2049 = (v617 & i31) | (v2050 & ~i31),
  v2050 = (v617 & i32) | (v2051 & ~i32),
  v2051 = (v982 & i33) | (v1560 & ~i33),
  v2052 = (v2053 & i21) | (v617 & ~i21),
  v2053 = (v2054 & i22) | (v617 & ~i22),
  v2054 = (v2055 & i29) | (v1587 & ~i29),
  v2055 = (v617 & i30) | (v2056 & ~i30),
  v2056 = (v617 & i31) | (v2057 & ~i31),
  v2057 = (v617 & i32) | (v2058 & ~i32),
  v2058 = (v991 & i33) | (v1581 & ~i33),
  v2059 = (v2060 & i21) | (v617 & ~i21),
  v2060 = (v2061 & i22) | (v617 & ~i22),
  v2061 = (v2062 & i29) | (v1608 & ~i29),
  v2062 = (v617 & i30) | (v2063 & ~i30),
  v2063 = (v617 & i31) | (v2064 & ~i31),
  v2064 = (v617 & i32) | (v2065 & ~i32),
  v2065 = (v1000 & i33) | (v1602 & ~i33),
  v2066 = (v617 & i11) | (v2067 & ~i11),
  v2067 = (v617 & i12) | (v2068 & ~i12),
  v2068 = (v617 & i13) | (v2069 & ~i13),
  v2069 = (v2070 & i14) | (v617 & ~i14),
  v2070 = (v2112 & i15) | (v2071 & ~i15),
  v2071 = (v2092 & i16) | (v2072 & ~i16),
  v2072 = (v2084 & i17) | (v2073 & ~i17),
  v2073 = (v2079 & i19) | (v2074 & ~i19),
  v2074 = (v2077 & i20) | (v2075 & ~i20),
  v2075 = (v2076 & i21) | (v617 & ~i21),
  v2076 = (v1009 & i22) | (v617 & ~i22),
  v2077 = (v2078 & i21) | (v617 & ~i21),
  v2078 = (v1030 & i22) | (v617 & ~i22),
  v2079 = (v2082 & i20) | (v2080 & ~i20),
  v2080 = (v2081 & i21) | (v617 & ~i21),
  v2081 = (v1052 & i22) | (v617 & ~i22),
  v2082 = (v2083 & i21) | (v617 & ~i21),
  v2083 = (v1073 & i22) | (v617 & ~i22),
  v2084 = (v2090 & i19) | (v2085 & ~i19),
  v2085 = (v2088 & i20) | (v2086 & ~i20),
  v2086 = (v2087 & i21) | (v617 & ~i21),
  v2087 = (v1096 & i22) | (v617 & ~i22),
  v2088 = (v2089 & i21) | (v617 & ~i21),
  v2089 = (v1117 & i22) | (v617 & ~i22),
  v2090 = (v2091 & i21) | (v617 & ~i21),
  v2091 = (v1138 & i22) | (v617 & ~i22),
  v2092 = (v2104 & i17) | (v2093 & ~i17),
  v2093 = (v2099 & i19) | (v2094 & ~i19),
  v2094 = (v2097 & i20) | (v2095 & ~i20),
  v2095 = (v2096 & i21) | (v617 & ~i21),
  v2096 = (v1162 & i22) | (v617 & ~i22),
  v2097 = (v2098 & i21) | (v617 & ~i21),
  v2098 = (v1183 & i22) | (v617 & ~i22),
  v2099 = (v2102 & i20) | (v2100 & ~i20),
  v2100 = (v2101 & i21) | (v617 & ~i21),
  v2101 = (v1205 & i22) | (v617 & ~i22),
  v2102 = (v2103 & i21) | (v617 & ~i21),
  v2103 = (v1226 & i22) | (v617 & ~i22),
  v2104 = (v2110 & i19) | (v2105 & ~i19),
  v2105 = (v2108 & i20) | (v2106 & ~i20),
  v2106 = (v2107 & i21) | (v617 & ~i21),
  v2107 = (v1249 & i22) | (v617 & ~i22),
  v2108 = (v2109 & i21) | (v617 & ~i21),
  v2109 = (v1270 & i22) | (v617 & ~i22),
  v2110 = (v2111 & i21) | (v617 & ~i21),
  v2111 = (v1291 & i22) | (v617 & ~i22),
  v2112 = (v2133 & i16) | (v2113 & ~i16),
  v2113 = (v2125 & i17) | (v2114 & ~i17),
  v2114 = (v2120 & i19) | (v2115 & ~i19),
  v2115 = (v2118 & i20) | (v2116 & ~i20),
  v2116 = (v2117 & i21) | (v617 & ~i21),
  v2117 = (v1316 & i22) | (v617 & ~i22),
  v2118 = (v2119 & i21) | (v617 & ~i21),
  v2119 = (v1337 & i22) | (v617 & ~i22),
  v2120 = (v2123 & i20) | (v2121 & ~i20),
  v2121 = (v2122 & i21) | (v617 & ~i21),
  v2122 = (v1359 & i22) | (v617 & ~i22),
  v2123 = (v2124 & i21) | (v617 & ~i21),
  v2124 = (v1380 & i22) | (v617 & ~i22),
  v2125 = (v2131 & i19) | (v2126 & ~i19),
  v2126 = (v2129 & i20) | (v2127 & ~i20),
  v2127 = (v2128 & i21) | (v617 & ~i21),
  v2128 = (v1403 & i22) | (v617 & ~i22),
  v2129 = (v2130 & i21) | (v617 & ~i21),
  v2130 = (v1424 & i22) | (v617 & ~i22),
  v2131 = (v2132 & i21) | (v617 & ~i21),
  v2132 = (v1445 & i22) | (v617 & ~i22),
  v2133 = (v2145 & i17) | (v2134 & ~i17),
  v2134 = (v2140 & i19) | (v2135 & ~i19),
  v2135 = (v2138 & i20) | (v2136 & ~i20),
  v2136 = (v2137 & i21) | (v617 & ~i21),
  v2137 = (v1469 & i22) | (v617 & ~i22),
  v2138 = (v2139 & i21) | (v617 & ~i21),
  v2139 = (v1490 & i22) | (v617 & ~i22),
  v2140 = (v2143 & i20) | (v2141 & ~i20),
  v2141 = (v2142 & i21) | (v617 & ~i21),
  v2142 = (v1512 & i22) | (v617 & ~i22),
  v2143 = (v2144 & i21) | (v617 & ~i21),
  v2144 = (v1533 & i22) | (v617 & ~i22),
  v2145 = (v2151 & i19) | (v2146 & ~i19),
  v2146 = (v2149 & i20) | (v2147 & ~i20),
  v2147 = (v2148 & i21) | (v617 & ~i21),
  v2148 = (v1556 & i22) | (v617 & ~i22),
  v2149 = (v2150 & i21) | (v617 & ~i21),
  v2150 = (v1577 & i22) | (v617 & ~i22),
  v2151 = (v2152 & i21) | (v617 & ~i21),
  v2152 = (v1598 & i22) | (v617 & ~i22),
  v2153 = (v63 & i2) | (v2154 & ~i2),
  v2154 = (v63 & i3) | (v2155 & ~i3),
  v2155 = (v3672 & i7) | (v2156 & ~i7),
  v2156 = (v3672 & i8) | (v2157 & ~i8),
  v2157 = (v3672 & i9) | (v2158 & ~i9),
  v2158 = (v3383 & i10) | (v2159 & ~i10),
  v2159 = (v3148 & i11) | (v2160 & ~i11),
  v2160 = (v3148 & i12) | (v2161 & ~i12),
  v2161 = (v3148 & i13) | (v2162 & ~i13),
  v2162 = (v2586 & i14) | (v2163 & ~i14),
  v2163 = (v2441 & i15) | (v2164 & ~i15),
  v2164 = (v2320 & i16) | (v2165 & ~i16),
  v2165 = (v2267 & i17) | (v2166 & ~i17),
  v2166 = (v2227 & i19) | (v2167 & ~i19),
  v2167 = (v2207 & i20) | (v2168 & ~i20),
  v2168 = (v2172 & i21) | (v2169 & ~i21),
  v2169 = (v63 & i30) | (v2170 & ~i30),
  v2170 = (v63 & i31) | (v2171 & ~i31),
  v2171 = (v63 & i32) | (v35 & ~i32),
  v2172 = (v2177 & i22) | (v2173 & ~i22),
  v2173 = (v63 & i30) | (v2174 & ~i30),
  v2174 = (v63 & i31) | (v2175 & ~i31),
  v2175 = (v63 & i32) | (v2176 & ~i32),
  v2176 = (v36 & i45) | (v6 & ~i45),
  v2177 = (v2193 & i25) | (v2178 & ~i25),
  v2178 = (v63 & i30) | (v2179 & ~i30),
  v2179 = (v63 & i31) | (v2180 & ~i31),
  v2180 = (v63 & i32) | (v2181 & ~i32),
  v2181 = (v2189 & i33) | (v2182 & ~i33),
  v2182 = (v2187 & i37) | (v2183 & ~i37),
  v2183 = (v2184 & i42) | (v2176 & ~i42),
  v2184 = (v2176 & i43) | (v2185 & ~i43),
  v2185 = (v2186 & i44) | (v2176 & ~i44),
  v2186 = (v36 & i45) | (v12 & ~i45),
  v2187 = (v2183 & i38) | (v2188 & ~i38),
  v2188 = (v2186 & i39) | (v2176 & ~i39),
  v2189 = (v2192 & i37) | (v2190 & ~i37),
  v2190 = (v2191 & i42) | (v2186 & ~i42),
  v2191 = (v2186 & i43) | (v2185 & ~i43),
  v2192 = (v2190 & i38) | (v2188 & ~i38),
  v2193 = (v63 & i30) | (v2194 & ~i30),
  v2194 = (v63 & i31) | (v2195 & ~i31),
  v2195 = (v63 & i32) | (v2196 & ~i32),
  v2196 = (v2197 & i33) | (v2182 & ~i33),
  v2197 = (v2206 & i36) | (v2198 & ~i36),
  v2198 = (v2205 & i37) | (v2199 & ~i37),
  v2199 = (v2201 & i38) | (v2200 & ~i38),
  v2200 = (v2183 & i39) | (v2201 & ~i39),
  v2201 = (v2190 & i41) | (v2202 & ~i41),
  v2202 = (v2191 & i42) | (v2203 & ~i42),
  v2203 = (v2186 & i43) | (v2204 & ~i43),
  v2204 = (v2176 & i44) | (v2186 & ~i44),
  v2205 = (v2201 & i38) | (v2188 & ~i38),
  v2206 = (v2205 & i37) | (v2201 & ~i37),
  v2207 = (v2211 & i21) | (v2208 & ~i21),
  v2208 = (v63 & i30) | (v2209 & ~i30),
  v2209 = (v63 & i31) | (v2210 & ~i31),
  v2210 = (v63 & i32) | (v41 & ~i32),
  v2211 = (v2215 & i22) | (v2212 & ~i22),
  v2212 = (v63 & i30) | (v2213 & ~i30),
  v2213 = (v63 & i31) | (v2214 & ~i31),
  v2214 = (v63 & i32) | (v2186 & ~i32),
  v2215 = (v2216 & i25) | (v2178 & ~i25),
  v2216 = (v63 & i30) | (v2217 & ~i30),
  v2217 = (v63 & i31) | (v2218 & ~i31),
  v2218 = (v63 & i32) | (v2219 & ~i32),
  v2219 = (v2220 & i33) | (v2182 & ~i33),
  v2220 = (v2226 & i36) | (v2221 & ~i36),
  v2221 = (v2225 & i37) | (v2222 & ~i37),
  v2222 = (v2224 & i38) | (v2223 & ~i38),
  v2223 = (v2224 & i39) | (v2183 & ~i39),
  v2224 = (v2190 & i41) | (v2191 & ~i41),
  v2225 = (v2224 & i38) | (v2188 & ~i38),
  v2226 = (v2225 & i37) | (v2224 & ~i37),
  v2227 = (v2249 & i20) | (v2228 & ~i20),
  v2228 = (v2229 & i21) | (v2169 & ~i21),
  v2229 = (v2230 & i22) | (v2173 & ~i22),
  v2230 = (v2231 & i25) | (v2178 & ~i25),
  v2231 = (v63 & i30) | (v2232 & ~i30),
  v2232 = (v63 & i31) | (v2233 & ~i31),
  v2233 = (v63 & i32) | (v2234 & ~i32),
  v2234 = (v2235 & i33) | (v2182 & ~i33),
  v2235 = (v2245 & i35) | (v2236 & ~i35),
  v2236 = (v2244 & i36) | (v2237 & ~i36),
  v2237 = (v2243 & i37) | (v2238 & ~i37),
  v2238 = (v2239 & i38) | (v2183 & ~i38),
  v2239 = (v2201 & i40) | (v2240 & ~i40),
  v2240 = (v2190 & i41) | (v2241 & ~i41),
  v2241 = (v2191 & i42) | (v2242 & ~i42),
  v2242 = (v2186 & i43) | (v2176 & ~i43),
  v2243 = (v2239 & i38) | (v2188 & ~i38),
  v2244 = (v2243 & i37) | (v2239 & ~i37),
  v2245 = (v2244 & i36) | (v2246 & ~i36),
  v2246 = (v2243 & i37) | (v2247 & ~i37),
  v2247 = (v2239 & i38) | (v2248 & ~i38),
  v2248 = (v2183 & i39) | (v2239 & ~i39),
  v2249 = (v2250 & i21) | (v2208 & ~i21),
  v2250 = (v2251 & i22) | (v2212 & ~i22),
  v2251 = (v2252 & i25) | (v2178 & ~i25),
  v2252 = (v63 & i30) | (v2253 & ~i30),
  v2253 = (v63 & i31) | (v2254 & ~i31),
  v2254 = (v63 & i32) | (v2255 & ~i32),
  v2255 = (v2256 & i33) | (v2182 & ~i33),
  v2256 = (v2263 & i35) | (v2257 & ~i35),
  v2257 = (v2262 & i36) | (v2258 & ~i36),
  v2258 = (v2261 & i37) | (v2259 & ~i37),
  v2259 = (v2260 & i38) | (v2183 & ~i38),
  v2260 = (v2224 & i40) | (v2240 & ~i40),
  v2261 = (v2260 & i38) | (v2188 & ~i38),
  v2262 = (v2261 & i37) | (v2260 & ~i37),
  v2263 = (v2262 & i36) | (v2264 & ~i36),
  v2264 = (v2261 & i37) | (v2265 & ~i37),
  v2265 = (v2260 & i38) | (v2266 & ~i38),
  v2266 = (v2260 & i39) | (v2183 & ~i39),
  v2267 = (v2305 & i19) | (v2268 & ~i19),
  v2268 = (v2287 & i20) | (v2269 & ~i20),
  v2269 = (v2270 & i21) | (v2169 & ~i21),
  v2270 = (v2271 & i22) | (v2173 & ~i22),
  v2271 = (v2272 & i25) | (v2178 & ~i25),
  v2272 = (v63 & i30) | (v2273 & ~i30),
  v2273 = (v63 & i31) | (v2274 & ~i31),
  v2274 = (v63 & i32) | (v2275 & ~i32),
  v2275 = (v2276 & i33) | (v2182 & ~i33),
  v2276 = (v2284 & i35) | (v2277 & ~i35),
  v2277 = (v2283 & i36) | (v2278 & ~i36),
  v2278 = (v2282 & i37) | (v2279 & ~i37),
  v2279 = (v2281 & i38) | (v2280 & ~i38),
  v2280 = (v2183 & i39) | (v2281 & ~i39),
  v2281 = (v2240 & i40) | (v2201 & ~i40),
  v2282 = (v2281 & i38) | (v2188 & ~i38),
  v2283 = (v2282 & i37) | (v2281 & ~i37),
  v2284 = (v2283 & i36) | (v2285 & ~i36),
  v2285 = (v2282 & i37) | (v2286 & ~i37),
  v2286 = (v2281 & i38) | (v2183 & ~i38),
  v2287 = (v2288 & i21) | (v2208 & ~i21),
  v2288 = (v2289 & i22) | (v2212 & ~i22),
  v2289 = (v2290 & i25) | (v2178 & ~i25),
  v2290 = (v63 & i30) | (v2291 & ~i30),
  v2291 = (v63 & i31) | (v2292 & ~i31),
  v2292 = (v63 & i32) | (v2293 & ~i32),
  v2293 = (v2294 & i33) | (v2182 & ~i33),
  v2294 = (v2302 & i35) | (v2295 & ~i35),
  v2295 = (v2301 & i36) | (v2296 & ~i36),
  v2296 = (v2300 & i37) | (v2297 & ~i37),
  v2297 = (v2299 & i38) | (v2298 & ~i38),
  v2298 = (v2299 & i39) | (v2183 & ~i39),
  v2299 = (v2240 & i40) | (v2224 & ~i40),
  v2300 = (v2299 & i38) | (v2188 & ~i38),
  v2301 = (v2300 & i37) | (v2299 & ~i37),
  v2302 = (v2301 & i36) | (v2303 & ~i36),
  v2303 = (v2300 & i37) | (v2304 & ~i37),
  v2304 = (v2299 & i38) | (v2183 & ~i38),
  v2305 = (v2318 & i20) | (v2306 & ~i20),
  v2306 = (v2307 & i21) | (v2169 & ~i21),
  v2307 = (v2308 & i22) | (v2173 & ~i22),
  v2308 = (v2309 & i25) | (v2178 & ~i25),
  v2309 = (v63 & i30) | (v2310 & ~i30),
  v2310 = (v63 & i31) | (v2311 & ~i31),
  v2311 = (v63 & i32) | (v2312 & ~i32),
  v2312 = (v2313 & i33) | (v2182 & ~i33),
  v2313 = (v2317 & i36) | (v2314 & ~i36),
  v2314 = (v2316 & i37) | (v2315 & ~i37),
  v2315 = (v2240 & i38) | (v2183 & ~i38),
  v2316 = (v2240 & i38) | (v2188 & ~i38),
  v2317 = (v2316 & i37) | (v2240 & ~i37),
  v2318 = (v2319 & i21) | (v2208 & ~i21),
  v2319 = (v2308 & i22) | (v2212 & ~i22),
  v2320 = (v2388 & i17) | (v2321 & ~i17),
  v2321 = (v2351 & i19) | (v2322 & ~i19),
  v2322 = (v2337 & i20) | (v2323 & ~i20),
  v2323 = (v2324 & i21) | (v2169 & ~i21),
  v2324 = (v2325 & i22) | (v2173 & ~i22),
  v2325 = (v2326 & i25) | (v2178 & ~i25),
  v2326 = (v63 & i30) | (v2327 & ~i30),
  v2327 = (v63 & i31) | (v2328 & ~i31),
  v2328 = (v63 & i32) | (v2329 & ~i32),
  v2329 = (v2330 & i33) | (v2182 & ~i33),
  v2330 = (v2336 & i36) | (v2331 & ~i36),
  v2331 = (v2335 & i37) | (v2332 & ~i37),
  v2332 = (v2334 & i38) | (v2333 & ~i38),
  v2333 = (v2183 & i39) | (v2334 & ~i39),
  v2334 = (v2241 & i41) | (v2202 & ~i41),
  v2335 = (v2334 & i38) | (v2188 & ~i38),
  v2336 = (v2335 & i37) | (v2334 & ~i37),
  v2337 = (v2338 & i21) | (v2208 & ~i21),
  v2338 = (v2339 & i22) | (v2212 & ~i22),
  v2339 = (v2340 & i25) | (v2178 & ~i25),
  v2340 = (v63 & i30) | (v2341 & ~i30),
  v2341 = (v63 & i31) | (v2342 & ~i31),
  v2342 = (v63 & i32) | (v2343 & ~i32),
  v2343 = (v2344 & i33) | (v2182 & ~i33),
  v2344 = (v2350 & i36) | (v2345 & ~i36),
  v2345 = (v2349 & i37) | (v2346 & ~i37),
  v2346 = (v2348 & i38) | (v2347 & ~i38),
  v2347 = (v2348 & i39) | (v2183 & ~i39),
  v2348 = (v2241 & i41) | (v2191 & ~i41),
  v2349 = (v2348 & i38) | (v2188 & ~i38),
  v2350 = (v2349 & i37) | (v2348 & ~i37),
  v2351 = (v2370 & i20) | (v2352 & ~i20),
  v2352 = (v2353 & i21) | (v2169 & ~i21),
  v2353 = (v2354 & i22) | (v2173 & ~i22),
  v2354 = (v2355 & i25) | (v2178 & ~i25),
  v2355 = (v63 & i30) | (v2356 & ~i30),
  v2356 = (v63 & i31) | (v2357 & ~i31),
  v2357 = (v63 & i32) | (v2358 & ~i32),
  v2358 = (v2359 & i33) | (v2182 & ~i33),
  v2359 = (v2366 & i35) | (v2360 & ~i35),
  v2360 = (v2365 & i36) | (v2361 & ~i36),
  v2361 = (v2364 & i37) | (v2362 & ~i37),
  v2362 = (v2363 & i38) | (v2183 & ~i38),
  v2363 = (v2334 & i40) | (v2241 & ~i40),
  v2364 = (v2363 & i38) | (v2188 & ~i38),
  v2365 = (v2364 & i37) | (v2363 & ~i37),
  v2366 = (v2365 & i36) | (v2367 & ~i36),
  v2367 = (v2364 & i37) | (v2368 & ~i37),
  v2368 = (v2363 & i38) | (v2369 & ~i38),
  v2369 = (v2183 & i39) | (v2363 & ~i39),
  v2370 = (v2371 & i21) | (v2208 & ~i21),
  v2371 = (v2372 & i22) | (v2212 & ~i22),
  v2372 = (v2373 & i25) | (v2178 & ~i25),
  v2373 = (v63 & i30) | (v2374 & ~i30),
  v2374 = (v63 & i31) | (v2375 & ~i31),
  v2375 = (v63 & i32) | (v2376 & ~i32),
  v2376 = (v2377 & i33) | (v2182 & ~i33),
  v2377 = (v2384 & i35) | (v2378 & ~i35),
  v2378 = (v2383 & i36) | (v2379 & ~i36),
  v2379 = (v2382 & i37) | (v2380 & ~i37),
  v2380 = (v2381 & i38) | (v2183 & ~i38),
  v2381 = (v2348 & i40) | (v2241 & ~i40),
  v2382 = (v2381 & i38) | (v2188 & ~i38),
  v2383 = (v2382 & i37) | (v2381 & ~i37),
  v2384 = (v2383 & i36) | (v2385 & ~i36),
  v2385 = (v2382 & i37) | (v2386 & ~i37),
  v2386 = (v2381 & i38) | (v2387 & ~i38),
  v2387 = (v2381 & i39) | (v2183 & ~i39),
  v2388 = (v2426 & i19) | (v2389 & ~i19),
  v2389 = (v2408 & i20) | (v2390 & ~i20),
  v2390 = (v2391 & i21) | (v2169 & ~i21),
  v2391 = (v2392 & i22) | (v2173 & ~i22),
  v2392 = (v2393 & i25) | (v2178 & ~i25),
  v2393 = (v63 & i30) | (v2394 & ~i30),
  v2394 = (v63 & i31) | (v2395 & ~i31),
  v2395 = (v63 & i32) | (v2396 & ~i32),
  v2396 = (v2397 & i33) | (v2182 & ~i33),
  v2397 = (v2405 & i35) | (v2398 & ~i35),
  v2398 = (v2404 & i36) | (v2399 & ~i36),
  v2399 = (v2403 & i37) | (v2400 & ~i37),
  v2400 = (v2402 & i38) | (v2401 & ~i38),
  v2401 = (v2183 & i39) | (v2402 & ~i39),
  v2402 = (v2241 & i40) | (v2334 & ~i40),
  v2403 = (v2402 & i38) | (v2188 & ~i38),
  v2404 = (v2403 & i37) | (v2402 & ~i37),
  v2405 = (v2404 & i36) | (v2406 & ~i36),
  v2406 = (v2403 & i37) | (v2407 & ~i37),
  v2407 = (v2402 & i38) | (v2183 & ~i38),
  v2408 = (v2409 & i21) | (v2208 & ~i21),
  v2409 = (v2410 & i22) | (v2212 & ~i22),
  v2410 = (v2411 & i25) | (v2178 & ~i25),
  v2411 = (v63 & i30) | (v2412 & ~i30),
  v2412 = (v63 & i31) | (v2413 & ~i31),
  v2413 = (v63 & i32) | (v2414 & ~i32),
  v2414 = (v2415 & i33) | (v2182 & ~i33),
  v2415 = (v2423 & i35) | (v2416 & ~i35),
  v2416 = (v2422 & i36) | (v2417 & ~i36),
  v2417 = (v2421 & i37) | (v2418 & ~i37),
  v2418 = (v2420 & i38) | (v2419 & ~i38),
  v2419 = (v2420 & i39) | (v2183 & ~i39),
  v2420 = (v2241 & i40) | (v2348 & ~i40),
  v2421 = (v2420 & i38) | (v2188 & ~i38),
  v2422 = (v2421 & i37) | (v2420 & ~i37),
  v2423 = (v2422 & i36) | (v2424 & ~i36),
  v2424 = (v2421 & i37) | (v2425 & ~i37),
  v2425 = (v2420 & i38) | (v2183 & ~i38),
  v2426 = (v2439 & i20) | (v2427 & ~i20),
  v2427 = (v2428 & i21) | (v2169 & ~i21),
  v2428 = (v2429 & i22) | (v2173 & ~i22),
  v2429 = (v2430 & i25) | (v2178 & ~i25),
  v2430 = (v63 & i30) | (v2431 & ~i30),
  v2431 = (v63 & i31) | (v2432 & ~i31),
  v2432 = (v63 & i32) | (v2433 & ~i32),
  v2433 = (v2434 & i33) | (v2182 & ~i33),
  v2434 = (v2438 & i36) | (v2435 & ~i36),
  v2435 = (v2437 & i37) | (v2436 & ~i37),
  v2436 = (v2241 & i38) | (v2183 & ~i38),
  v2437 = (v2241 & i38) | (v2188 & ~i38),
  v2438 = (v2437 & i37) | (v2241 & ~i37),
  v2439 = (v2440 & i21) | (v2208 & ~i21),
  v2440 = (v2429 & i22) | (v2212 & ~i22),
  v2441 = (v2514 & i16) | (v2442 & ~i16),
  v2442 = (v2484 & i17) | (v2443 & ~i17),
  v2443 = (v2465 & i19) | (v2444 & ~i19),
  v2444 = (v2455 & i20) | (v2445 & ~i20),
  v2445 = (v2446 & i21) | (v2169 & ~i21),
  v2446 = (v2447 & i22) | (v2173 & ~i22),
  v2447 = (v2448 & i25) | (v2178 & ~i25),
  v2448 = (v63 & i30) | (v2449 & ~i30),
  v2449 = (v63 & i31) | (v2450 & ~i31),
  v2450 = (v63 & i32) | (v2451 & ~i32),
  v2451 = (v2452 & i33) | (v2182 & ~i33),
  v2452 = (v2453 & i36) | (v2198 & ~i36),
  v2453 = (v2205 & i37) | (v2454 & ~i37),
  v2454 = (v2201 & i38) | (v2183 & ~i38),
  v2455 = (v2456 & i21) | (v2208 & ~i21),
  v2456 = (v2457 & i22) | (v2212 & ~i22),
  v2457 = (v2458 & i25) | (v2178 & ~i25),
  v2458 = (v63 & i30) | (v2459 & ~i30),
  v2459 = (v63 & i31) | (v2460 & ~i31),
  v2460 = (v63 & i32) | (v2461 & ~i32),
  v2461 = (v2462 & i33) | (v2182 & ~i33),
  v2462 = (v2463 & i36) | (v2221 & ~i36),
  v2463 = (v2225 & i37) | (v2464 & ~i37),
  v2464 = (v2224 & i38) | (v2183 & ~i38),
  v2465 = (v2475 & i20) | (v2466 & ~i20),
  v2466 = (v2467 & i21) | (v2169 & ~i21),
  v2467 = (v2468 & i22) | (v2173 & ~i22),
  v2468 = (v2469 & i25) | (v2178 & ~i25),
  v2469 = (v63 & i30) | (v2470 & ~i30),
  v2470 = (v63 & i31) | (v2471 & ~i31),
  v2471 = (v63 & i32) | (v2472 & ~i32),
  v2472 = (v2473 & i33) | (v2182 & ~i33),
  v2473 = (v2474 & i35) | (v2237 & ~i35),
  v2474 = (v2237 & i36) | (v2246 & ~i36),
  v2475 = (v2476 & i21) | (v2208 & ~i21),
  v2476 = (v2477 & i22) | (v2212 & ~i22),
  v2477 = (v2478 & i25) | (v2178 & ~i25),
  v2478 = (v63 & i30) | (v2479 & ~i30),
  v2479 = (v63 & i31) | (v2480 & ~i31),
  v2480 = (v63 & i32) | (v2481 & ~i32),
  v2481 = (v2482 & i33) | (v2182 & ~i33),
  v2482 = (v2483 & i35) | (v2258 & ~i35),
  v2483 = (v2258 & i36) | (v2264 & ~i36),
  v2484 = (v2504 & i19) | (v2485 & ~i19),
  v2485 = (v2495 & i20) | (v2486 & ~i20),
  v2486 = (v2487 & i21) | (v2169 & ~i21),
  v2487 = (v2488 & i22) | (v2173 & ~i22),
  v2488 = (v2489 & i25) | (v2178 & ~i25),
  v2489 = (v63 & i30) | (v2490 & ~i30),
  v2490 = (v63 & i31) | (v2491 & ~i31),
  v2491 = (v63 & i32) | (v2492 & ~i32),
  v2492 = (v2493 & i33) | (v2182 & ~i33),
  v2493 = (v2285 & i35) | (v2494 & ~i35),
  v2494 = (v2285 & i36) | (v2278 & ~i36),
  v2495 = (v2496 & i21) | (v2208 & ~i21),
  v2496 = (v2497 & i22) | (v2212 & ~i22),
  v2497 = (v2498 & i25) | (v2178 & ~i25),
  v2498 = (v63 & i30) | (v2499 & ~i30),
  v2499 = (v63 & i31) | (v2500 & ~i31),
  v2500 = (v63 & i32) | (v2501 & ~i32),
  v2501 = (v2502 & i33) | (v2182 & ~i33),
  v2502 = (v2303 & i35) | (v2503 & ~i35),
  v2503 = (v2303 & i36) | (v2296 & ~i36),
  v2504 = (v2512 & i20) | (v2505 & ~i20),
  v2505 = (v2506 & i21) | (v2169 & ~i21),
  v2506 = (v2507 & i22) | (v2173 & ~i22),
  v2507 = (v2508 & i25) | (v2178 & ~i25),
  v2508 = (v63 & i30) | (v2509 & ~i30),
  v2509 = (v63 & i31) | (v2510 & ~i31),
  v2510 = (v63 & i32) | (v2511 & ~i32),
  v2511 = (v2314 & i33) | (v2182 & ~i33),
  v2512 = (v2513 & i21) | (v2208 & ~i21),
  v2513 = (v2507 & i22) | (v2212 & ~i22),
  v2514 = (v2556 & i17) | (v2515 & ~i17),
  v2515 = (v2537 & i19) | (v2516 & ~i19),
  v2516 = (v2527 & i20) | (v2517 & ~i20),
  v2517 = (v2518 & i21) | (v2169 & ~i21),
  v2518 = (v2519 & i22) | (v2173 & ~i22),
  v2519 = (v2520 & i25) | (v2178 & ~i25),
  v2520 = (v63 & i30) | (v2521 & ~i30),
  v2521 = (v63 & i31) | (v2522 & ~i31),
  v2522 = (v63 & i32) | (v2523 & ~i32),
  v2523 = (v2524 & i33) | (v2182 & ~i33),
  v2524 = (v2525 & i36) | (v2331 & ~i36),
  v2525 = (v2335 & i37) | (v2526 & ~i37),
  v2526 = (v2334 & i38) | (v2183 & ~i38),
  v2527 = (v2528 & i21) | (v2208 & ~i21),
  v2528 = (v2529 & i22) | (v2212 & ~i22),
  v2529 = (v2530 & i25) | (v2178 & ~i25),
  v2530 = (v63 & i30) | (v2531 & ~i30),
  v2531 = (v63 & i31) | (v2532 & ~i31),
  v2532 = (v63 & i32) | (v2533 & ~i32),
  v2533 = (v2534 & i33) | (v2182 & ~i33),
  v2534 = (v2535 & i36) | (v2345 & ~i36),
  v2535 = (v2349 & i37) | (v2536 & ~i37),
  v2536 = (v2348 & i38) | (v2183 & ~i38),
  v2537 = (v2547 & i20) | (v2538 & ~i20),
  v2538 = (v2539 & i21) | (v2169 & ~i21),
  v2539 = (v2540 & i22) | (v2173 & ~i22),
  v2540 = (v2541 & i25) | (v2178 & ~i25),
  v2541 = (v63 & i30) | (v2542 & ~i30),
  v2542 = (v63 & i31) | (v2543 & ~i31),
  v2543 = (v63 & i32) | (v2544 & ~i32),
  v2544 = (v2545 & i33) | (v2182 & ~i33),
  v2545 = (v2546 & i35) | (v2361 & ~i35),
  v2546 = (v2361 & i36) | (v2367 & ~i36),
  v2547 = (v2548 & i21) | (v2208 & ~i21),
  v2548 = (v2549 & i22) | (v2212 & ~i22),
  v2549 = (v2550 & i25) | (v2178 & ~i25),
  v2550 = (v63 & i30) | (v2551 & ~i30),
  v2551 = (v63 & i31) | (v2552 & ~i31),
  v2552 = (v63 & i32) | (v2553 & ~i32),
  v2553 = (v2554 & i33) | (v2182 & ~i33),
  v2554 = (v2555 & i35) | (v2379 & ~i35),
  v2555 = (v2379 & i36) | (v2385 & ~i36),
  v2556 = (v2576 & i19) | (v2557 & ~i19),
  v2557 = (v2567 & i20) | (v2558 & ~i20),
  v2558 = (v2559 & i21) | (v2169 & ~i21),
  v2559 = (v2560 & i22) | (v2173 & ~i22),
  v2560 = (v2561 & i25) | (v2178 & ~i25),
  v2561 = (v63 & i30) | (v2562 & ~i30),
  v2562 = (v63 & i31) | (v2563 & ~i31),
  v2563 = (v63 & i32) | (v2564 & ~i32),
  v2564 = (v2565 & i33) | (v2182 & ~i33),
  v2565 = (v2406 & i35) | (v2566 & ~i35),
  v2566 = (v2406 & i36) | (v2399 & ~i36),
  v2567 = (v2568 & i21) | (v2208 & ~i21),
  v2568 = (v2569 & i22) | (v2212 & ~i22),
  v2569 = (v2570 & i25) | (v2178 & ~i25),
  v2570 = (v63 & i30) | (v2571 & ~i30),
  v2571 = (v63 & i31) | (v2572 & ~i31),
  v2572 = (v63 & i32) | (v2573 & ~i32),
  v2573 = (v2574 & i33) | (v2182 & ~i33),
  v2574 = (v2424 & i35) | (v2575 & ~i35),
  v2575 = (v2424 & i36) | (v2417 & ~i36),
  v2576 = (v2584 & i20) | (v2577 & ~i20),
  v2577 = (v2578 & i21) | (v2169 & ~i21),
  v2578 = (v2579 & i22) | (v2173 & ~i22),
  v2579 = (v2580 & i25) | (v2178 & ~i25),
  v2580 = (v63 & i30) | (v2581 & ~i30),
  v2581 = (v63 & i31) | (v2582 & ~i31),
  v2582 = (v63 & i32) | (v2583 & ~i32),
  v2583 = (v2435 & i33) | (v2182 & ~i33),
  v2584 = (v2585 & i21) | (v2208 & ~i21),
  v2585 = (v2579 & i22) | (v2212 & ~i22),
  v2586 = (v2919 & i15) | (v2587 & ~i15),
  v2587 = (v2756 & i16) | (v2588 & ~i16),
  v2588 = (v2685 & i17) | (v2589 & ~i17),
  v2589 = (v2633 & i19) | (v2590 & ~i19),
  v2590 = (v2611 & i20) | (v2591 & ~i20),
  v2591 = (v2592 & i21) | (v2169 & ~i21),
  v2592 = (v2593 & i22) | (v2173 & ~i22),
  v2593 = (v2605 & i25) | (v2594 & ~i25),
  v2594 = (v63 & i30) | (v2595 & ~i30),
  v2595 = (v63 & i31) | (v2596 & ~i31),
  v2596 = (v63 & i32) | (v2597 & ~i32),
  v2597 = (v2189 & i33) | (v2598 & ~i33),
  v2598 = (v2604 & i36) | (v2599 & ~i36),
  v2599 = (v2603 & i37) | (v2600 & ~i37),
  v2600 = (v2602 & i38) | (v2601 & ~i38),
  v2601 = (v2190 & i39) | (v2602 & ~i39),
  v2602 = (v2183 & i41) | (v2184 & ~i41),
  v2603 = (v2602 & i38) | (v2188 & ~i38),
  v2604 = (v2603 & i37) | (v2602 & ~i37),
  v2605 = (v63 & i30) | (v2606 & ~i30),
  v2606 = (v63 & i31) | (v2607 & ~i31),
  v2607 = (v63 & i32) | (v2608 & ~i32),
  v2608 = (v2610 & i33) | (v2609 & ~i33),
  v2609 = (v2598 & i34) | (v2182 & ~i34),
  v2610 = (v2189 & i34) | (v2197 & ~i34),
  v2611 = (v2612 & i21) | (v2208 & ~i21),
  v2612 = (v2613 & i22) | (v2212 & ~i22),
  v2613 = (v2627 & i25) | (v2614 & ~i25),
  v2614 = (v63 & i30) | (v2615 & ~i30),
  v2615 = (v63 & i31) | (v2616 & ~i31),
  v2616 = (v63 & i32) | (v2617 & ~i32),
  v2617 = (v2189 & i33) | (v2618 & ~i33),
  v2618 = (v2626 & i36) | (v2619 & ~i36),
  v2619 = (v2625 & i37) | (v2620 & ~i37),
  v2620 = (v2622 & i38) | (v2621 & ~i38),
  v2621 = (v2622 & i39) | (v2190 & ~i39),
  v2622 = (v2183 & i41) | (v2623 & ~i41),
  v2623 = (v2184 & i42) | (v2624 & ~i42),
  v2624 = (v2176 & i43) | (v2204 & ~i43),
  v2625 = (v2622 & i38) | (v2188 & ~i38),
  v2626 = (v2625 & i37) | (v2622 & ~i37),
  v2627 = (v63 & i30) | (v2628 & ~i30),
  v2628 = (v63 & i31) | (v2629 & ~i31),
  v2629 = (v63 & i32) | (v2630 & ~i32),
  v2630 = (v2632 & i33) | (v2631 & ~i33),
  v2631 = (v2618 & i34) | (v2182 & ~i34),
  v2632 = (v2189 & i34) | (v2220 & ~i34),
  v2633 = (v2661 & i20) | (v2634 & ~i20),
  v2634 = (v2635 & i21) | (v2169 & ~i21),
  v2635 = (v2636 & i22) | (v2173 & ~i22),
  v2636 = (v2655 & i25) | (v2637 & ~i25),
  v2637 = (v63 & i30) | (v2638 & ~i30),
  v2638 = (v63 & i31) | (v2639 & ~i31),
  v2639 = (v63 & i32) | (v2640 & ~i32),
  v2640 = (v2189 & i33) | (v2641 & ~i33),
  v2641 = (v2651 & i35) | (v2642 & ~i35),
  v2642 = (v2650 & i36) | (v2643 & ~i36),
  v2643 = (v2649 & i37) | (v2644 & ~i37),
  v2644 = (v2645 & i38) | (v2190 & ~i38),
  v2645 = (v2602 & i40) | (v2646 & ~i40),
  v2646 = (v2183 & i41) | (v2647 & ~i41),
  v2647 = (v2184 & i42) | (v2648 & ~i42),
  v2648 = (v2176 & i43) | (v2186 & ~i43),
  v2649 = (v2645 & i38) | (v2188 & ~i38),
  v2650 = (v2649 & i37) | (v2645 & ~i37),
  v2651 = (v2650 & i36) | (v2652 & ~i36),
  v2652 = (v2649 & i37) | (v2653 & ~i37),
  v2653 = (v2645 & i38) | (v2654 & ~i38),
  v2654 = (v2190 & i39) | (v2645 & ~i39),
  v2655 = (v63 & i30) | (v2656 & ~i30),
  v2656 = (v63 & i31) | (v2657 & ~i31),
  v2657 = (v63 & i32) | (v2658 & ~i32),
  v2658 = (v2660 & i33) | (v2659 & ~i33),
  v2659 = (v2641 & i34) | (v2182 & ~i34),
  v2660 = (v2189 & i34) | (v2235 & ~i34),
  v2661 = (v2662 & i21) | (v2208 & ~i21),
  v2662 = (v2663 & i22) | (v2212 & ~i22),
  v2663 = (v2679 & i25) | (v2664 & ~i25),
  v2664 = (v63 & i30) | (v2665 & ~i30),
  v2665 = (v63 & i31) | (v2666 & ~i31),
  v2666 = (v63 & i32) | (v2667 & ~i32),
  v2667 = (v2189 & i33) | (v2668 & ~i33),
  v2668 = (v2675 & i35) | (v2669 & ~i35),
  v2669 = (v2674 & i36) | (v2670 & ~i36),
  v2670 = (v2673 & i37) | (v2671 & ~i37),
  v2671 = (v2672 & i38) | (v2190 & ~i38),
  v2672 = (v2622 & i40) | (v2646 & ~i40),
  v2673 = (v2672 & i38) | (v2188 & ~i38),
  v2674 = (v2673 & i37) | (v2672 & ~i37),
  v2675 = (v2674 & i36) | (v2676 & ~i36),
  v2676 = (v2673 & i37) | (v2677 & ~i37),
  v2677 = (v2672 & i38) | (v2678 & ~i38),
  v2678 = (v2672 & i39) | (v2190 & ~i39),
  v2679 = (v63 & i30) | (v2680 & ~i30),
  v2680 = (v63 & i31) | (v2681 & ~i31),
  v2681 = (v63 & i32) | (v2682 & ~i32),
  v2682 = (v2684 & i33) | (v2683 & ~i33),
  v2683 = (v2668 & i34) | (v2182 & ~i34),
  v2684 = (v2189 & i34) | (v2256 & ~i34),
  v2685 = (v2735 & i19) | (v2686 & ~i19),
  v2686 = (v2711 & i20) | (v2687 & ~i20),
  v2687 = (v2688 & i21) | (v2169 & ~i21),
  v2688 = (v2689 & i22) | (v2173 & ~i22),
  v2689 = (v2705 & i25) | (v2690 & ~i25),
  v2690 = (v63 & i30) | (v2691 & ~i30),
  v2691 = (v63 & i31) | (v2692 & ~i31),
  v2692 = (v63 & i32) | (v2693 & ~i32),
  v2693 = (v2189 & i33) | (v2694 & ~i33),
  v2694 = (v2702 & i35) | (v2695 & ~i35),
  v2695 = (v2701 & i36) | (v2696 & ~i36),
  v2696 = (v2700 & i37) | (v2697 & ~i37),
  v2697 = (v2699 & i38) | (v2698 & ~i38),
  v2698 = (v2190 & i39) | (v2699 & ~i39),
  v2699 = (v2646 & i40) | (v2602 & ~i40),
  v2700 = (v2699 & i38) | (v2188 & ~i38),
  v2701 = (v2700 & i37) | (v2699 & ~i37),
  v2702 = (v2701 & i36) | (v2703 & ~i36),
  v2703 = (v2700 & i37) | (v2704 & ~i37),
  v2704 = (v2699 & i38) | (v2190 & ~i38),
  v2705 = (v63 & i30) | (v2706 & ~i30),
  v2706 = (v63 & i31) | (v2707 & ~i31),
  v2707 = (v63 & i32) | (v2708 & ~i32),
  v2708 = (v2710 & i33) | (v2709 & ~i33),
  v2709 = (v2694 & i34) | (v2182 & ~i34),
  v2710 = (v2189 & i34) | (v2276 & ~i34),
  v2711 = (v2712 & i21) | (v2208 & ~i21),
  v2712 = (v2713 & i22) | (v2212 & ~i22),
  v2713 = (v2729 & i25) | (v2714 & ~i25),
  v2714 = (v63 & i30) | (v2715 & ~i30),
  v2715 = (v63 & i31) | (v2716 & ~i31),
  v2716 = (v63 & i32) | (v2717 & ~i32),
  v2717 = (v2189 & i33) | (v2718 & ~i33),
  v2718 = (v2726 & i35) | (v2719 & ~i35),
  v2719 = (v2725 & i36) | (v2720 & ~i36),
  v2720 = (v2724 & i37) | (v2721 & ~i37),
  v2721 = (v2723 & i38) | (v2722 & ~i38),
  v2722 = (v2723 & i39) | (v2190 & ~i39),
  v2723 = (v2646 & i40) | (v2622 & ~i40),
  v2724 = (v2723 & i38) | (v2188 & ~i38),
  v2725 = (v2724 & i37) | (v2723 & ~i37),
  v2726 = (v2725 & i36) | (v2727 & ~i36),
  v2727 = (v2724 & i37) | (v2728 & ~i37),
  v2728 = (v2723 & i38) | (v2190 & ~i38),
  v2729 = (v63 & i30) | (v2730 & ~i30),
  v2730 = (v63 & i31) | (v2731 & ~i31),
  v2731 = (v63 & i32) | (v2732 & ~i32),
  v2732 = (v2734 & i33) | (v2733 & ~i33),
  v2733 = (v2718 & i34) | (v2182 & ~i34),
  v2734 = (v2189 & i34) | (v2294 & ~i34),
  v2735 = (v2754 & i20) | (v2736 & ~i20),
  v2736 = (v2737 & i21) | (v2169 & ~i21),
  v2737 = (v2738 & i22) | (v2173 & ~i22),
  v2738 = (v2748 & i25) | (v2739 & ~i25),
  v2739 = (v63 & i30) | (v2740 & ~i30),
  v2740 = (v63 & i31) | (v2741 & ~i31),
  v2741 = (v63 & i32) | (v2742 & ~i32),
  v2742 = (v2189 & i33) | (v2743 & ~i33),
  v2743 = (v2747 & i36) | (v2744 & ~i36),
  v2744 = (v2746 & i37) | (v2745 & ~i37),
  v2745 = (v2646 & i38) | (v2190 & ~i38),
  v2746 = (v2646 & i38) | (v2188 & ~i38),
  v2747 = (v2746 & i37) | (v2646 & ~i37),
  v2748 = (v63 & i30) | (v2749 & ~i30),
  v2749 = (v63 & i31) | (v2750 & ~i31),
  v2750 = (v63 & i32) | (v2751 & ~i32),
  v2751 = (v2753 & i33) | (v2752 & ~i33),
  v2752 = (v2743 & i34) | (v2182 & ~i34),
  v2753 = (v2189 & i34) | (v2313 & ~i34),
  v2754 = (v2755 & i21) | (v2208 & ~i21),
  v2755 = (v2738 & i22) | (v2212 & ~i22),
  v2756 = (v2848 & i17) | (v2757 & ~i17),
  v2757 = (v2799 & i19) | (v2758 & ~i19),
  v2758 = (v2779 & i20) | (v2759 & ~i20),
  v2759 = (v2760 & i21) | (v2169 & ~i21),
  v2760 = (v2761 & i22) | (v2173 & ~i22),
  v2761 = (v2773 & i25) | (v2762 & ~i25),
  v2762 = (v63 & i30) | (v2763 & ~i30),
  v2763 = (v63 & i31) | (v2764 & ~i31),
  v2764 = (v63 & i32) | (v2765 & ~i32),
  v2765 = (v2189 & i33) | (v2766 & ~i33),
  v2766 = (v2772 & i36) | (v2767 & ~i36),
  v2767 = (v2771 & i37) | (v2768 & ~i37),
  v2768 = (v2770 & i38) | (v2769 & ~i38),
  v2769 = (v2190 & i39) | (v2770 & ~i39),
  v2770 = (v2647 & i41) | (v2184 & ~i41),
  v2771 = (v2770 & i38) | (v2188 & ~i38),
  v2772 = (v2771 & i37) | (v2770 & ~i37),
  v2773 = (v63 & i30) | (v2774 & ~i30),
  v2774 = (v63 & i31) | (v2775 & ~i31),
  v2775 = (v63 & i32) | (v2776 & ~i32),
  v2776 = (v2778 & i33) | (v2777 & ~i33),
  v2777 = (v2766 & i34) | (v2182 & ~i34),
  v2778 = (v2189 & i34) | (v2330 & ~i34),
  v2779 = (v2780 & i21) | (v2208 & ~i21),
  v2780 = (v2781 & i22) | (v2212 & ~i22),
  v2781 = (v2793 & i25) | (v2782 & ~i25),
  v2782 = (v63 & i30) | (v2783 & ~i30),
  v2783 = (v63 & i31) | (v2784 & ~i31),
  v2784 = (v63 & i32) | (v2785 & ~i32),
  v2785 = (v2189 & i33) | (v2786 & ~i33),
  v2786 = (v2792 & i36) | (v2787 & ~i36),
  v2787 = (v2791 & i37) | (v2788 & ~i37),
  v2788 = (v2790 & i38) | (v2789 & ~i38),
  v2789 = (v2790 & i39) | (v2190 & ~i39),
  v2790 = (v2647 & i41) | (v2623 & ~i41),
  v2791 = (v2790 & i38) | (v2188 & ~i38),
  v2792 = (v2791 & i37) | (v2790 & ~i37),
  v2793 = (v63 & i30) | (v2794 & ~i30),
  v2794 = (v63 & i31) | (v2795 & ~i31),
  v2795 = (v63 & i32) | (v2796 & ~i32),
  v2796 = (v2798 & i33) | (v2797 & ~i33),
  v2797 = (v2786 & i34) | (v2182 & ~i34),
  v2798 = (v2189 & i34) | (v2344 & ~i34),
  v2799 = (v2824 & i20) | (v2800 & ~i20),
  v2800 = (v2801 & i21) | (v2169 & ~i21),
  v2801 = (v2802 & i22) | (v2173 & ~i22),
  v2802 = (v2818 & i25) | (v2803 & ~i25),
  v2803 = (v63 & i30) | (v2804 & ~i30),
  v2804 = (v63 & i31) | (v2805 & ~i31),
  v2805 = (v63 & i32) | (v2806 & ~i32),
  v2806 = (v2189 & i33) | (v2807 & ~i33),
  v2807 = (v2814 & i35) | (v2808 & ~i35),
  v2808 = (v2813 & i36) | (v2809 & ~i36),
  v2809 = (v2812 & i37) | (v2810 & ~i37),
  v2810 = (v2811 & i38) | (v2190 & ~i38),
  v2811 = (v2770 & i40) | (v2647 & ~i40),
  v2812 = (v2811 & i38) | (v2188 & ~i38),
  v2813 = (v2812 & i37) | (v2811 & ~i37),
  v2814 = (v2813 & i36) | (v2815 & ~i36),
  v2815 = (v2812 & i37) | (v2816 & ~i37),
  v2816 = (v2811 & i38) | (v2817 & ~i38),
  v2817 = (v2190 & i39) | (v2811 & ~i39),
  v2818 = (v63 & i30) | (v2819 & ~i30),
  v2819 = (v63 & i31) | (v2820 & ~i31),
  v2820 = (v63 & i32) | (v2821 & ~i32),
  v2821 = (v2823 & i33) | (v2822 & ~i33),
  v2822 = (v2807 & i34) | (v2182 & ~i34),
  v2823 = (v2189 & i34) | (v2359 & ~i34),
  v2824 = (v2825 & i21) | (v2208 & ~i21),
  v2825 = (v2826 & i22) | (v2212 & ~i22),
  v2826 = (v2842 & i25) | (v2827 & ~i25),
  v2827 = (v63 & i30) | (v2828 & ~i30),
  v2828 = (v63 & i31) | (v2829 & ~i31),
  v2829 = (v63 & i32) | (v2830 & ~i32),
  v2830 = (v2189 & i33) | (v2831 & ~i33),
  v2831 = (v2838 & i35) | (v2832 & ~i35),
  v2832 = (v2837 & i36) | (v2833 & ~i36),
  v2833 = (v2836 & i37) | (v2834 & ~i37),
  v2834 = (v2835 & i38) | (v2190 & ~i38),
  v2835 = (v2790 & i40) | (v2647 & ~i40),
  v2836 = (v2835 & i38) | (v2188 & ~i38),
  v2837 = (v2836 & i37) | (v2835 & ~i37),
  v2838 = (v2837 & i36) | (v2839 & ~i36),
  v2839 = (v2836 & i37) | (v2840 & ~i37),
  v2840 = (v2835 & i38) | (v2841 & ~i38),
  v2841 = (v2835 & i39) | (v2190 & ~i39),
  v2842 = (v63 & i30) | (v2843 & ~i30),
  v2843 = (v63 & i31) | (v2844 & ~i31),
  v2844 = (v63 & i32) | (v2845 & ~i32),
  v2845 = (v2847 & i33) | (v2846 & ~i33),
  v2846 = (v2831 & i34) | (v2182 & ~i34),
  v2847 = (v2189 & i34) | (v2377 & ~i34),
  v2848 = (v2898 & i19) | (v2849 & ~i19),
  v2849 = (v2874 & i20) | (v2850 & ~i20),
  v2850 = (v2851 & i21) | (v2169 & ~i21),
  v2851 = (v2852 & i22) | (v2173 & ~i22),
  v2852 = (v2868 & i25) | (v2853 & ~i25),
  v2853 = (v63 & i30) | (v2854 & ~i30),
  v2854 = (v63 & i31) | (v2855 & ~i31),
  v2855 = (v63 & i32) | (v2856 & ~i32),
  v2856 = (v2189 & i33) | (v2857 & ~i33),
  v2857 = (v2865 & i35) | (v2858 & ~i35),
  v2858 = (v2864 & i36) | (v2859 & ~i36),
  v2859 = (v2863 & i37) | (v2860 & ~i37),
  v2860 = (v2862 & i38) | (v2861 & ~i38),
  v2861 = (v2190 & i39) | (v2862 & ~i39),
  v2862 = (v2647 & i40) | (v2770 & ~i40),
  v2863 = (v2862 & i38) | (v2188 & ~i38),
  v2864 = (v2863 & i37) | (v2862 & ~i37),
  v2865 = (v2864 & i36) | (v2866 & ~i36),
  v2866 = (v2863 & i37) | (v2867 & ~i37),
  v2867 = (v2862 & i38) | (v2190 & ~i38),
  v2868 = (v63 & i30) | (v2869 & ~i30),
  v2869 = (v63 & i31) | (v2870 & ~i31),
  v2870 = (v63 & i32) | (v2871 & ~i32),
  v2871 = (v2873 & i33) | (v2872 & ~i33),
  v2872 = (v2857 & i34) | (v2182 & ~i34),
  v2873 = (v2189 & i34) | (v2397 & ~i34),
  v2874 = (v2875 & i21) | (v2208 & ~i21),
  v2875 = (v2876 & i22) | (v2212 & ~i22),
  v2876 = (v2892 & i25) | (v2877 & ~i25),
  v2877 = (v63 & i30) | (v2878 & ~i30),
  v2878 = (v63 & i31) | (v2879 & ~i31),
  v2879 = (v63 & i32) | (v2880 & ~i32),
  v2880 = (v2189 & i33) | (v2881 & ~i33),
  v2881 = (v2889 & i35) | (v2882 & ~i35),
  v2882 = (v2888 & i36) | (v2883 & ~i36),
  v2883 = (v2887 & i37) | (v2884 & ~i37),
  v2884 = (v2886 & i38) | (v2885 & ~i38),
  v2885 = (v2886 & i39) | (v2190 & ~i39),
  v2886 = (v2647 & i40) | (v2790 & ~i40),
  v2887 = (v2886 & i38) | (v2188 & ~i38),
  v2888 = (v2887 & i37) | (v2886 & ~i37),
  v2889 = (v2888 & i36) | (v2890 & ~i36),
  v2890 = (v2887 & i37) | (v2891 & ~i37),
  v2891 = (v2886 & i38) | (v2190 & ~i38),
  v2892 = (v63 & i30) | (v2893 & ~i30),
  v2893 = (v63 & i31) | (v2894 & ~i31),
  v2894 = (v63 & i32) | (v2895 & ~i32),
  v2895 = (v2897 & i33) | (v2896 & ~i33),
  v2896 = (v2881 & i34) | (v2182 & ~i34),
  v2897 = (v2189 & i34) | (v2415 & ~i34),
  v2898 = (v2917 & i20) | (v2899 & ~i20),
  v2899 = (v2900 & i21) | (v2169 & ~i21),
  v2900 = (v2901 & i22) | (v2173 & ~i22),
  v2901 = (v2911 & i25) | (v2902 & ~i25),
  v2902 = (v63 & i30) | (v2903 & ~i30),
  v2903 = (v63 & i31) | (v2904 & ~i31),
  v2904 = (v63 & i32) | (v2905 & ~i32),
  v2905 = (v2189 & i33) | (v2906 & ~i33),
  v2906 = (v2910 & i36) | (v2907 & ~i36),
  v2907 = (v2909 & i37) | (v2908 & ~i37),
  v2908 = (v2647 & i38) | (v2190 & ~i38),
  v2909 = (v2647 & i38) | (v2188 & ~i38),
  v2910 = (v2909 & i37) | (v2647 & ~i37),
  v2911 = (v63 & i30) | (v2912 & ~i30),
  v2912 = (v63 & i31) | (v2913 & ~i31),
  v2913 = (v63 & i32) | (v2914 & ~i32),
  v2914 = (v2916 & i33) | (v2915 & ~i33),
  v2915 = (v2906 & i34) | (v2182 & ~i34),
  v2916 = (v2189 & i34) | (v2434 & ~i34),
  v2917 = (v2918 & i21) | (v2208 & ~i21),
  v2918 = (v2901 & i22) | (v2212 & ~i22),
  v2919 = (v3034 & i16) | (v2920 & ~i16),
  v2920 = (v2986 & i17) | (v2921 & ~i17),
  v2921 = (v2955 & i19) | (v2922 & ~i19),
  v2922 = (v2939 & i20) | (v2923 & ~i20),
  v2923 = (v2924 & i21) | (v2169 & ~i21),
  v2924 = (v2925 & i22) | (v2173 & ~i22),
  v2925 = (v2933 & i25) | (v2926 & ~i25),
  v2926 = (v63 & i30) | (v2927 & ~i30),
  v2927 = (v63 & i31) | (v2928 & ~i31),
  v2928 = (v63 & i32) | (v2929 & ~i32),
  v2929 = (v2189 & i33) | (v2930 & ~i33),
  v2930 = (v2931 & i36) | (v2599 & ~i36),
  v2931 = (v2603 & i37) | (v2932 & ~i37),
  v2932 = (v2602 & i38) | (v2190 & ~i38),
  v2933 = (v63 & i30) | (v2934 & ~i30),
  v2934 = (v63 & i31) | (v2935 & ~i31),
  v2935 = (v63 & i32) | (v2936 & ~i32),
  v2936 = (v2938 & i33) | (v2937 & ~i33),
  v2937 = (v2930 & i34) | (v2182 & ~i34),
  v2938 = (v2189 & i34) | (v2452 & ~i34),
  v2939 = (v2940 & i21) | (v2208 & ~i21),
  v2940 = (v2941 & i22) | (v2212 & ~i22),
  v2941 = (v2949 & i25) | (v2942 & ~i25),
  v2942 = (v63 & i30) | (v2943 & ~i30),
  v2943 = (v63 & i31) | (v2944 & ~i31),
  v2944 = (v63 & i32) | (v2945 & ~i32),
  v2945 = (v2189 & i33) | (v2946 & ~i33),
  v2946 = (v2947 & i36) | (v2619 & ~i36),
  v2947 = (v2625 & i37) | (v2948 & ~i37),
  v2948 = (v2622 & i38) | (v2190 & ~i38),
  v2949 = (v63 & i30) | (v2950 & ~i30),
  v2950 = (v63 & i31) | (v2951 & ~i31),
  v2951 = (v63 & i32) | (v2952 & ~i32),
  v2952 = (v2954 & i33) | (v2953 & ~i33),
  v2953 = (v2946 & i34) | (v2182 & ~i34),
  v2954 = (v2189 & i34) | (v2462 & ~i34),
  v2955 = (v2971 & i20) | (v2956 & ~i20),
  v2956 = (v2957 & i21) | (v2169 & ~i21),
  v2957 = (v2958 & i22) | (v2173 & ~i22),
  v2958 = (v2965 & i25) | (v2959 & ~i25),
  v2959 = (v63 & i30) | (v2960 & ~i30),
  v2960 = (v63 & i31) | (v2961 & ~i31),
  v2961 = (v63 & i32) | (v2962 & ~i32),
  v2962 = (v2189 & i33) | (v2963 & ~i33),
  v2963 = (v2964 & i35) | (v2643 & ~i35),
  v2964 = (v2643 & i36) | (v2652 & ~i36),
  v2965 = (v63 & i30) | (v2966 & ~i30),
  v2966 = (v63 & i31) | (v2967 & ~i31),
  v2967 = (v63 & i32) | (v2968 & ~i32),
  v2968 = (v2970 & i33) | (v2969 & ~i33),
  v2969 = (v2963 & i34) | (v2182 & ~i34),
  v2970 = (v2189 & i34) | (v2473 & ~i34),
  v2971 = (v2972 & i21) | (v2208 & ~i21),
  v2972 = (v2973 & i22) | (v2212 & ~i22),
  v2973 = (v2980 & i25) | (v2974 & ~i25),
  v2974 = (v63 & i30) | (v2975 & ~i30),
  v2975 = (v63 & i31) | (v2976 & ~i31),
  v2976 = (v63 & i32) | (v2977 & ~i32),
  v2977 = (v2189 & i33) | (v2978 & ~i33),
  v2978 = (v2979 & i35) | (v2670 & ~i35),
  v2979 = (v2670 & i36) | (v2676 & ~i36),
  v2980 = (v63 & i30) | (v2981 & ~i30),
  v2981 = (v63 & i31) | (v2982 & ~i31),
  v2982 = (v63 & i32) | (v2983 & ~i32),
  v2983 = (v2985 & i33) | (v2984 & ~i33),
  v2984 = (v2978 & i34) | (v2182 & ~i34),
  v2985 = (v2189 & i34) | (v2482 & ~i34),
  v2986 = (v3018 & i19) | (v2987 & ~i19),
  v2987 = (v3003 & i20) | (v2988 & ~i20),
  v2988 = (v2989 & i21) | (v2169 & ~i21),
  v2989 = (v2990 & i22) | (v2173 & ~i22),
  v2990 = (v2997 & i25) | (v2991 & ~i25),
  v2991 = (v63 & i30) | (v2992 & ~i30),
  v2992 = (v63 & i31) | (v2993 & ~i31),
  v2993 = (v63 & i32) | (v2994 & ~i32),
  v2994 = (v2189 & i33) | (v2995 & ~i33),
  v2995 = (v2703 & i35) | (v2996 & ~i35),
  v2996 = (v2703 & i36) | (v2696 & ~i36),
  v2997 = (v63 & i30) | (v2998 & ~i30),
  v2998 = (v63 & i31) | (v2999 & ~i31),
  v2999 = (v63 & i32) | (v3000 & ~i32),
  v3000 = (v3002 & i33) | (v3001 & ~i33),
  v3001 = (v2995 & i34) | (v2182 & ~i34),
  v3002 = (v2189 & i34) | (v2493 & ~i34),
  v3003 = (v3004 & i21) | (v2208 & ~i21),
  v3004 = (v3005 & i22) | (v2212 & ~i22),
  v3005 = (v3012 & i25) | (v3006 & ~i25),
  v3006 = (v63 & i30) | (v3007 & ~i30),
  v3007 = (v63 & i31) | (v3008 & ~i31),
  v3008 = (v63 & i32) | (v3009 & ~i32),
  v3009 = (v2189 & i33) | (v3010 & ~i33),
  v3010 = (v2727 & i35) | (v3011 & ~i35),
  v3011 = (v2727 & i36) | (v2720 & ~i36),
  v3012 = (v63 & i30) | (v3013 & ~i30),
  v3013 = (v63 & i31) | (v3014 & ~i31),
  v3014 = (v63 & i32) | (v3015 & ~i32),
  v3015 = (v3017 & i33) | (v3016 & ~i33),
  v3016 = (v3010 & i34) | (v2182 & ~i34),
  v3017 = (v2189 & i34) | (v2502 & ~i34),
  v3018 = (v3032 & i20) | (v3019 & ~i20),
  v3019 = (v3020 & i21) | (v2169 & ~i21),
  v3020 = (v3021 & i22) | (v2173 & ~i22),
  v3021 = (v3026 & i25) | (v3022 & ~i25),
  v3022 = (v63 & i30) | (v3023 & ~i30),
  v3023 = (v63 & i31) | (v3024 & ~i31),
  v3024 = (v63 & i32) | (v3025 & ~i32),
  v3025 = (v2189 & i33) | (v2744 & ~i33),
  v3026 = (v63 & i30) | (v3027 & ~i30),
  v3027 = (v63 & i31) | (v3028 & ~i31),
  v3028 = (v63 & i32) | (v3029 & ~i32),
  v3029 = (v3031 & i33) | (v3030 & ~i33),
  v3030 = (v2744 & i34) | (v2182 & ~i34),
  v3031 = (v2189 & i34) | (v2314 & ~i34),
  v3032 = (v3033 & i21) | (v2208 & ~i21),
  v3033 = (v3021 & i22) | (v2212 & ~i22),
  v3034 = (v3100 & i17) | (v3035 & ~i17),
  v3035 = (v3069 & i19) | (v3036 & ~i19),
  v3036 = (v3053 & i20) | (v3037 & ~i20),
  v3037 = (v3038 & i21) | (v2169 & ~i21),
  v3038 = (v3039 & i22) | (v2173 & ~i22),
  v3039 = (v3047 & i25) | (v3040 & ~i25),
  v3040 = (v63 & i30) | (v3041 & ~i30),
  v3041 = (v63 & i31) | (v3042 & ~i31),
  v3042 = (v63 & i32) | (v3043 & ~i32),
  v3043 = (v2189 & i33) | (v3044 & ~i33),
  v3044 = (v3045 & i36) | (v2767 & ~i36),
  v3045 = (v2771 & i37) | (v3046 & ~i37),
  v3046 = (v2770 & i38) | (v2190 & ~i38),
  v3047 = (v63 & i30) | (v3048 & ~i30),
  v3048 = (v63 & i31) | (v3049 & ~i31),
  v3049 = (v63 & i32) | (v3050 & ~i32),
  v3050 = (v3052 & i33) | (v3051 & ~i33),
  v3051 = (v3044 & i34) | (v2182 & ~i34),
  v3052 = (v2189 & i34) | (v2524 & ~i34),
  v3053 = (v3054 & i21) | (v2208 & ~i21),
  v3054 = (v3055 & i22) | (v2212 & ~i22),
  v3055 = (v3063 & i25) | (v3056 & ~i25),
  v3056 = (v63 & i30) | (v3057 & ~i30),
  v3057 = (v63 & i31) | (v3058 & ~i31),
  v3058 = (v63 & i32) | (v3059 & ~i32),
  v3059 = (v2189 & i33) | (v3060 & ~i33),
  v3060 = (v3061 & i36) | (v2787 & ~i36),
  v3061 = (v2791 & i37) | (v3062 & ~i37),
  v3062 = (v2790 & i38) | (v2190 & ~i38),
  v3063 = (v63 & i30) | (v3064 & ~i30),
  v3064 = (v63 & i31) | (v3065 & ~i31),
  v3065 = (v63 & i32) | (v3066 & ~i32),
  v3066 = (v3068 & i33) | (v3067 & ~i33),
  v3067 = (v3060 & i34) | (v2182 & ~i34),
  v3068 = (v2189 & i34) | (v2534 & ~i34),
  v3069 = (v3085 & i20) | (v3070 & ~i20),
  v3070 = (v3071 & i21) | (v2169 & ~i21),
  v3071 = (v3072 & i22) | (v2173 & ~i22),
  v3072 = (v3079 & i25) | (v3073 & ~i25),
  v3073 = (v63 & i30) | (v3074 & ~i30),
  v3074 = (v63 & i31) | (v3075 & ~i31),
  v3075 = (v63 & i32) | (v3076 & ~i32),
  v3076 = (v2189 & i33) | (v3077 & ~i33),
  v3077 = (v3078 & i35) | (v2809 & ~i35),
  v3078 = (v2809 & i36) | (v2815 & ~i36),
  v3079 = (v63 & i30) | (v3080 & ~i30),
  v3080 = (v63 & i31) | (v3081 & ~i31),
  v3081 = (v63 & i32) | (v3082 & ~i32),
  v3082 = (v3084 & i33) | (v3083 & ~i33),
  v3083 = (v3077 & i34) | (v2182 & ~i34),
  v3084 = (v2189 & i34) | (v2545 & ~i34),
  v3085 = (v3086 & i21) | (v2208 & ~i21),
  v3086 = (v3087 & i22) | (v2212 & ~i22),
  v3087 = (v3094 & i25) | (v3088 & ~i25),
  v3088 = (v63 & i30) | (v3089 & ~i30),
  v3089 = (v63 & i31) | (v3090 & ~i31),
  v3090 = (v63 & i32) | (v3091 & ~i32),
  v3091 = (v2189 & i33) | (v3092 & ~i33),
  v3092 = (v3093 & i35) | (v2833 & ~i35),
  v3093 = (v2833 & i36) | (v2839 & ~i36),
  v3094 = (v63 & i30) | (v3095 & ~i30),
  v3095 = (v63 & i31) | (v3096 & ~i31),
  v3096 = (v63 & i32) | (v3097 & ~i32),
  v3097 = (v3099 & i33) | (v3098 & ~i33),
  v3098 = (v3092 & i34) | (v2182 & ~i34),
  v3099 = (v2189 & i34) | (v2554 & ~i34),
  v3100 = (v3132 & i19) | (v3101 & ~i19),
  v3101 = (v3117 & i20) | (v3102 & ~i20),
  v3102 = (v3103 & i21) | (v2169 & ~i21),
  v3103 = (v3104 & i22) | (v2173 & ~i22),
  v3104 = (v3111 & i25) | (v3105 & ~i25),
  v3105 = (v63 & i30) | (v3106 & ~i30),
  v3106 = (v63 & i31) | (v3107 & ~i31),
  v3107 = (v63 & i32) | (v3108 & ~i32),
  v3108 = (v2189 & i33) | (v3109 & ~i33),
  v3109 = (v2866 & i35) | (v3110 & ~i35),
  v3110 = (v2866 & i36) | (v2859 & ~i36),
  v3111 = (v63 & i30) | (v3112 & ~i30),
  v3112 = (v63 & i31) | (v3113 & ~i31),
  v3113 = (v63 & i32) | (v3114 & ~i32),
  v3114 = (v3116 & i33) | (v3115 & ~i33),
  v3115 = (v3109 & i34) | (v2182 & ~i34),
  v3116 = (v2189 & i34) | (v2565 & ~i34),
  v3117 = (v3118 & i21) | (v2208 & ~i21),
  v3118 = (v3119 & i22) | (v2212 & ~i22),
  v3119 = (v3126 & i25) | (v3120 & ~i25),
  v3120 = (v63 & i30) | (v3121 & ~i30),
  v3121 = (v63 & i31) | (v3122 & ~i31),
  v3122 = (v63 & i32) | (v3123 & ~i32),
  v3123 = (v2189 & i33) | (v3124 & ~i33),
  v3124 = (v2890 & i35) | (v3125 & ~i35),
  v3125 = (v2890 & i36) | (v2883 & ~i36),
  v3126 = (v63 & i30) | (v3127 & ~i30),
  v3127 = (v63 & i31) | (v3128 & ~i31),
  v3128 = (v63 & i32) | (v3129 & ~i32),
  v3129 = (v3131 & i33) | (v3130 & ~i33),
  v3130 = (v3124 & i34) | (v2182 & ~i34),
  v3131 = (v2189 & i34) | (v2574 & ~i34),
  v3132 = (v3146 & i20) | (v3133 & ~i20),
  v3133 = (v3134 & i21) | (v2169 & ~i21),
  v3134 = (v3135 & i22) | (v2173 & ~i22),
  v3135 = (v3140 & i25) | (v3136 & ~i25),
  v3136 = (v63 & i30) | (v3137 & ~i30),
  v3137 = (v63 & i31) | (v3138 & ~i31),
  v3138 = (v63 & i32) | (v3139 & ~i32),
  v3139 = (v2189 & i33) | (v2907 & ~i33),
  v3140 = (v63 & i30) | (v3141 & ~i30),
  v3141 = (v63 & i31) | (v3142 & ~i31),
  v3142 = (v63 & i32) | (v3143 & ~i32),
  v3143 = (v3145 & i33) | (v3144 & ~i33),
  v3144 = (v2907 & i34) | (v2182 & ~i34),
  v3145 = (v2189 & i34) | (v2435 & ~i34),
  v3146 = (v3147 & i21) | (v2208 & ~i21),
  v3147 = (v3135 & i22) | (v2212 & ~i22),
  v3148 = (v3266 & i15) | (v3149 & ~i15),
  v3149 = (v3208 & i16) | (v3150 & ~i16),
  v3150 = (v3182 & i17) | (v3151 & ~i17),
  v3151 = (v3167 & i19) | (v3152 & ~i19),
  v3152 = (v3160 & i20) | (v3153 & ~i20),
  v3153 = (v3154 & i21) | (v2169 & ~i21),
  v3154 = (v3155 & i22) | (v2173 & ~i22),
  v3155 = (v3156 & i25) | (v2178 & ~i25),
  v3156 = (v63 & i30) | (v3157 & ~i30),
  v3157 = (v63 & i31) | (v3158 & ~i31),
  v3158 = (v63 & i32) | (v3159 & ~i32),
  v3159 = (v2610 & i33) | (v2182 & ~i33),
  v3160 = (v3161 & i21) | (v2208 & ~i21),
  v3161 = (v3162 & i22) | (v2212 & ~i22),
  v3162 = (v3163 & i25) | (v2178 & ~i25),
  v3163 = (v63 & i30) | (v3164 & ~i30),
  v3164 = (v63 & i31) | (v3165 & ~i31),
  v3165 = (v63 & i32) | (v3166 & ~i32),
  v3166 = (v2632 & i33) | (v2182 & ~i33),
  v3167 = (v3175 & i20) | (v3168 & ~i20),
  v3168 = (v3169 & i21) | (v2169 & ~i21),
  v3169 = (v3170 & i22) | (v2173 & ~i22),
  v3170 = (v3171 & i25) | (v2178 & ~i25),
  v3171 = (v63 & i30) | (v3172 & ~i30),
  v3172 = (v63 & i31) | (v3173 & ~i31),
  v3173 = (v63 & i32) | (v3174 & ~i32),
  v3174 = (v2660 & i33) | (v2182 & ~i33),
  v3175 = (v3176 & i21) | (v2208 & ~i21),
  v3176 = (v3177 & i22) | (v2212 & ~i22),
  v3177 = (v3178 & i25) | (v2178 & ~i25),
  v3178 = (v63 & i30) | (v3179 & ~i30),
  v3179 = (v63 & i31) | (v3180 & ~i31),
  v3180 = (v63 & i32) | (v3181 & ~i32),
  v3181 = (v2684 & i33) | (v2182 & ~i33),
  v3182 = (v3198 & i19) | (v3183 & ~i19),
  v3183 = (v3191 & i20) | (v3184 & ~i20),
  v3184 = (v3185 & i21) | (v2169 & ~i21),
  v3185 = (v3186 & i22) | (v2173 & ~i22),
  v3186 = (v3187 & i25) | (v2178 & ~i25),
  v3187 = (v63 & i30) | (v3188 & ~i30),
  v3188 = (v63 & i31) | (v3189 & ~i31),
  v3189 = (v63 & i32) | (v3190 & ~i32),
  v3190 = (v2710 & i33) | (v2182 & ~i33),
  v3191 = (v3192 & i21) | (v2208 & ~i21),
  v3192 = (v3193 & i22) | (v2212 & ~i22),
  v3193 = (v3194 & i25) | (v2178 & ~i25),
  v3194 = (v63 & i30) | (v3195 & ~i30),
  v3195 = (v63 & i31) | (v3196 & ~i31),
  v3196 = (v63 & i32) | (v3197 & ~i32),
  v3197 = (v2734 & i33) | (v2182 & ~i33),
  v3198 = (v3206 & i20) | (v3199 & ~i20),
  v3199 = (v3200 & i21) | (v2169 & ~i21),
  v3200 = (v3201 & i22) | (v2173 & ~i22),
  v3201 = (v3202 & i25) | (v2178 & ~i25),
  v3202 = (v63 & i30) | (v3203 & ~i30),
  v3203 = (v63 & i31) | (v3204 & ~i31),
  v3204 = (v63 & i32) | (v3205 & ~i32),
  v3205 = (v2753 & i33) | (v2182 & ~i33),
  v3206 = (v3207 & i21) | (v2208 & ~i21),
  v3207 = (v3201 & i22) | (v2212 & ~i22),
  v3208 = (v3240 & i17) | (v3209 & ~i17),
  v3209 = (v3225 & i19) | (v3210 & ~i19),
  v3210 = (v3218 & i20) | (v3211 & ~i20),
  v3211 = (v3212 & i21) | (v2169 & ~i21),
  v3212 = (v3213 & i22) | (v2173 & ~i22),
  v3213 = (v3214 & i25) | (v2178 & ~i25),
  v3214 = (v63 & i30) | (v3215 & ~i30),
  v3215 = (v63 & i31) | (v3216 & ~i31),
  v3216 = (v63 & i32) | (v3217 & ~i32),
  v3217 = (v2778 & i33) | (v2182 & ~i33),
  v3218 = (v3219 & i21) | (v2208 & ~i21),
  v3219 = (v3220 & i22) | (v2212 & ~i22),
  v3220 = (v3221 & i25) | (v2178 & ~i25),
  v3221 = (v63 & i30) | (v3222 & ~i30),
  v3222 = (v63 & i31) | (v3223 & ~i31),
  v3223 = (v63 & i32) | (v3224 & ~i32),
  v3224 = (v2798 & i33) | (v2182 & ~i33),
  v3225 = (v3233 & i20) | (v3226 & ~i20),
  v3226 = (v3227 & i21) | (v2169 & ~i21),
  v3227 = (v3228 & i22) | (v2173 & ~i22),
  v3228 = (v3229 & i25) | (v2178 & ~i25),
  v3229 = (v63 & i30) | (v3230 & ~i30),
  v3230 = (v63 & i31) | (v3231 & ~i31),
  v3231 = (v63 & i32) | (v3232 & ~i32),
  v3232 = (v2823 & i33) | (v2182 & ~i33),
  v3233 = (v3234 & i21) | (v2208 & ~i21),
  v3234 = (v3235 & i22) | (v2212 & ~i22),
  v3235 = (v3236 & i25) | (v2178 & ~i25),
  v3236 = (v63 & i30) | (v3237 & ~i30),
  v3237 = (v63 & i31) | (v3238 & ~i31),
  v3238 = (v63 & i32) | (v3239 & ~i32),
  v3239 = (v2847 & i33) | (v2182 & ~i33),
  v3240 = (v3256 & i19) | (v3241 & ~i19),
  v3241 = (v3249 & i20) | (v3242 & ~i20),
  v3242 = (v3243 & i21) | (v2169 & ~i21),
  v3243 = (v3244 & i22) | (v2173 & ~i22),
  v3244 = (v3245 & i25) | (v2178 & ~i25),
  v3245 = (v63 & i30) | (v3246 & ~i30),
  v3246 = (v63 & i31) | (v3247 & ~i31),
  v3247 = (v63 & i32) | (v3248 & ~i32),
  v3248 = (v2873 & i33) | (v2182 & ~i33),
  v3249 = (v3250 & i21) | (v2208 & ~i21),
  v3250 = (v3251 & i22) | (v2212 & ~i22),
  v3251 = (v3252 & i25) | (v2178 & ~i25),
  v3252 = (v63 & i30) | (v3253 & ~i30),
  v3253 = (v63 & i31) | (v3254 & ~i31),
  v3254 = (v63 & i32) | (v3255 & ~i32),
  v3255 = (v2897 & i33) | (v2182 & ~i33),
  v3256 = (v3264 & i20) | (v3257 & ~i20),
  v3257 = (v3258 & i21) | (v2169 & ~i21),
  v3258 = (v3259 & i22) | (v2173 & ~i22),
  v3259 = (v3260 & i25) | (v2178 & ~i25),
  v3260 = (v63 & i30) | (v3261 & ~i30),
  v3261 = (v63 & i31) | (v3262 & ~i31),
  v3262 = (v63 & i32) | (v3263 & ~i32),
  v3263 = (v2916 & i33) | (v2182 & ~i33),
  v3264 = (v3265 & i21) | (v2208 & ~i21),
  v3265 = (v3259 & i22) | (v2212 & ~i22),
  v3266 = (v3325 & i16) | (v3267 & ~i16),
  v3267 = (v3299 & i17) | (v3268 & ~i17),
  v3268 = (v3284 & i19) | (v3269 & ~i19),
  v3269 = (v3277 & i20) | (v3270 & ~i20),
  v3270 = (v3271 & i21) | (v2169 & ~i21),
  v3271 = (v3272 & i22) | (v2173 & ~i22),
  v3272 = (v3273 & i25) | (v2178 & ~i25),
  v3273 = (v63 & i30) | (v3274 & ~i30),
  v3274 = (v63 & i31) | (v3275 & ~i31),
  v3275 = (v63 & i32) | (v3276 & ~i32),
  v3276 = (v2938 & i33) | (v2182 & ~i33),
  v3277 = (v3278 & i21) | (v2208 & ~i21),
  v3278 = (v3279 & i22) | (v2212 & ~i22),
  v3279 = (v3280 & i25) | (v2178 & ~i25),
  v3280 = (v63 & i30) | (v3281 & ~i30),
  v3281 = (v63 & i31) | (v3282 & ~i31),
  v3282 = (v63 & i32) | (v3283 & ~i32),
  v3283 = (v2954 & i33) | (v2182 & ~i33),
  v3284 = (v3292 & i20) | (v3285 & ~i20),
  v3285 = (v3286 & i21) | (v2169 & ~i21),
  v3286 = (v3287 & i22) | (v2173 & ~i22),
  v3287 = (v3288 & i25) | (v2178 & ~i25),
  v3288 = (v63 & i30) | (v3289 & ~i30),
  v3289 = (v63 & i31) | (v3290 & ~i31),
  v3290 = (v63 & i32) | (v3291 & ~i32),
  v3291 = (v2970 & i33) | (v2182 & ~i33),
  v3292 = (v3293 & i21) | (v2208 & ~i21),
  v3293 = (v3294 & i22) | (v2212 & ~i22),
  v3294 = (v3295 & i25) | (v2178 & ~i25),
  v3295 = (v63 & i30) | (v3296 & ~i30),
  v3296 = (v63 & i31) | (v3297 & ~i31),
  v3297 = (v63 & i32) | (v3298 & ~i32),
  v3298 = (v2985 & i33) | (v2182 & ~i33),
  v3299 = (v3315 & i19) | (v3300 & ~i19),
  v3300 = (v3308 & i20) | (v3301 & ~i20),
  v3301 = (v3302 & i21) | (v2169 & ~i21),
  v3302 = (v3303 & i22) | (v2173 & ~i22),
  v3303 = (v3304 & i25) | (v2178 & ~i25),
  v3304 = (v63 & i30) | (v3305 & ~i30),
  v3305 = (v63 & i31) | (v3306 & ~i31),
  v3306 = (v63 & i32) | (v3307 & ~i32),
  v3307 = (v3002 & i33) | (v2182 & ~i33),
  v3308 = (v3309 & i21) | (v2208 & ~i21),
  v3309 = (v3310 & i22) | (v2212 & ~i22),
  v3310 = (v3311 & i25) | (v2178 & ~i25),
  v3311 = (v63 & i30) | (v3312 & ~i30),
  v3312 = (v63 & i31) | (v3313 & ~i31),
  v3313 = (v63 & i32) | (v3314 & ~i32),
  v3314 = (v3017 & i33) | (v2182 & ~i33),
  v3315 = (v3323 & i20) | (v3316 & ~i20),
  v3316 = (v3317 & i21) | (v2169 & ~i21),
  v3317 = (v3318 & i22) | (v2173 & ~i22),
  v3318 = (v3319 & i25) | (v2178 & ~i25),
  v3319 = (v63 & i30) | (v3320 & ~i30),
  v3320 = (v63 & i31) | (v3321 & ~i31),
  v3321 = (v63 & i32) | (v3322 & ~i32),
  v3322 = (v3031 & i33) | (v2182 & ~i33),
  v3323 = (v3324 & i21) | (v2208 & ~i21),
  v3324 = (v3318 & i22) | (v2212 & ~i22),
  v3325 = (v3357 & i17) | (v3326 & ~i17),
  v3326 = (v3342 & i19) | (v3327 & ~i19),
  v3327 = (v3335 & i20) | (v3328 & ~i20),
  v3328 = (v3329 & i21) | (v2169 & ~i21),
  v3329 = (v3330 & i22) | (v2173 & ~i22),
  v3330 = (v3331 & i25) | (v2178 & ~i25),
  v3331 = (v63 & i30) | (v3332 & ~i30),
  v3332 = (v63 & i31) | (v3333 & ~i31),
  v3333 = (v63 & i32) | (v3334 & ~i32),
  v3334 = (v3052 & i33) | (v2182 & ~i33),
  v3335 = (v3336 & i21) | (v2208 & ~i21),
  v3336 = (v3337 & i22) | (v2212 & ~i22),
  v3337 = (v3338 & i25) | (v2178 & ~i25),
  v3338 = (v63 & i30) | (v3339 & ~i30),
  v3339 = (v63 & i31) | (v3340 & ~i31),
  v3340 = (v63 & i32) | (v3341 & ~i32),
  v3341 = (v3068 & i33) | (v2182 & ~i33),
  v3342 = (v3350 & i20) | (v3343 & ~i20),
  v3343 = (v3344 & i21) | (v2169 & ~i21),
  v3344 = (v3345 & i22) | (v2173 & ~i22),
  v3345 = (v3346 & i25) | (v2178 & ~i25),
  v3346 = (v63 & i30) | (v3347 & ~i30),
  v3347 = (v63 & i31) | (v3348 & ~i31),
  v3348 = (v63 & i32) | (v3349 & ~i32),
  v3349 = (v3084 & i33) | (v2182 & ~i33),
  v3350 = (v3351 & i21) | (v2208 & ~i21),
  v3351 = (v3352 & i22) | (v2212 & ~i22),
  v3352 = (v3353 & i25) | (v2178 & ~i25),
  v3353 = (v63 & i30) | (v3354 & ~i30),
  v3354 = (v63 & i31) | (v3355 & ~i31),
  v3355 = (v63 & i32) | (v3356 & ~i32),
  v3356 = (v3099 & i33) | (v2182 & ~i33),
  v3357 = (v3373 & i19) | (v3358 & ~i19),
  v3358 = (v3366 & i20) | (v3359 & ~i20),
  v3359 = (v3360 & i21) | (v2169 & ~i21),
  v3360 = (v3361 & i22) | (v2173 & ~i22),
  v3361 = (v3362 & i25) | (v2178 & ~i25),
  v3362 = (v63 & i30) | (v3363 & ~i30),
  v3363 = (v63 & i31) | (v3364 & ~i31),
  v3364 = (v63 & i32) | (v3365 & ~i32),
  v3365 = (v3116 & i33) | (v2182 & ~i33),
  v3366 = (v3367 & i21) | (v2208 & ~i21),
  v3367 = (v3368 & i22) | (v2212 & ~i22),
  v3368 = (v3369 & i25) | (v2178 & ~i25),
  v3369 = (v63 & i30) | (v3370 & ~i30),
  v3370 = (v63 & i31) | (v3371 & ~i31),
  v3371 = (v63 & i32) | (v3372 & ~i32),
  v3372 = (v3131 & i33) | (v2182 & ~i33),
  v3373 = (v3381 & i20) | (v3374 & ~i20),
  v3374 = (v3375 & i21) | (v2169 & ~i21),
  v3375 = (v3376 & i22) | (v2173 & ~i22),
  v3376 = (v3377 & i25) | (v2178 & ~i25),
  v3377 = (v63 & i30) | (v3378 & ~i30),
  v3378 = (v63 & i31) | (v3379 & ~i31),
  v3379 = (v63 & i32) | (v3380 & ~i32),
  v3380 = (v3145 & i33) | (v2182 & ~i33),
  v3381 = (v3382 & i21) | (v2208 & ~i21),
  v3382 = (v3376 & i22) | (v2212 & ~i22),
  v3383 = (v3577 & i11) | (v3384 & ~i11),
  v3384 = (v3577 & i12) | (v3385 & ~i12),
  v3385 = (v3577 & i13) | (v3386 & ~i13),
  v3386 = (v3482 & i14) | (v3387 & ~i14),
  v3387 = (v3435 & i15) | (v3388 & ~i15),
  v3388 = (v3412 & i16) | (v3389 & ~i16),
  v3389 = (v3401 & i17) | (v3390 & ~i17),
  v3390 = (v3396 & i19) | (v3391 & ~i19),
  v3391 = (v3394 & i20) | (v3392 & ~i20),
  v3392 = (v3393 & i21) | (v2169 & ~i21),
  v3393 = (v2193 & i22) | (v2173 & ~i22),
  v3394 = (v3395 & i21) | (v2208 & ~i21),
  v3395 = (v2216 & i22) | (v2212 & ~i22),
  v3396 = (v3399 & i20) | (v3397 & ~i20),
  v3397 = (v3398 & i21) | (v2169 & ~i21),
  v3398 = (v2231 & i22) | (v2173 & ~i22),
  v3399 = (v3400 & i21) | (v2208 & ~i21),
  v3400 = (v2252 & i22) | (v2212 & ~i22),
  v3401 = (v3407 & i19) | (v3402 & ~i19),
  v3402 = (v3405 & i20) | (v3403 & ~i20),
  v3403 = (v3404 & i21) | (v2169 & ~i21),
  v3404 = (v2272 & i22) | (v2173 & ~i22),
  v3405 = (v3406 & i21) | (v2208 & ~i21),
  v3406 = (v2290 & i22) | (v2212 & ~i22),
  v3407 = (v3410 & i20) | (v3408 & ~i20),
  v3408 = (v3409 & i21) | (v2169 & ~i21),
  v3409 = (v2309 & i22) | (v2173 & ~i22),
  v3410 = (v3411 & i21) | (v2208 & ~i21),
  v3411 = (v2309 & i22) | (v2212 & ~i22),
  v3412 = (v3424 & i17) | (v3413 & ~i17),
  v3413 = (v3419 & i19) | (v3414 & ~i19),
  v3414 = (v3417 & i20) | (v3415 & ~i20),
  v3415 = (v3416 & i21) | (v2169 & ~i21),
  v3416 = (v2326 & i22) | (v2173 & ~i22),
  v3417 = (v3418 & i21) | (v2208 & ~i21),
  v3418 = (v2340 & i22) | (v2212 & ~i22),
  v3419 = (v3422 & i20) | (v3420 & ~i20),
  v3420 = (v3421 & i21) | (v2169 & ~i21),
  v3421 = (v2355 & i22) | (v2173 & ~i22),
  v3422 = (v3423 & i21) | (v2208 & ~i21),
  v3423 = (v2373 & i22) | (v2212 & ~i22),
  v3424 = (v3430 & i19) | (v3425 & ~i19),
  v3425 = (v3428 & i20) | (v3426 & ~i20),
  v3426 = (v3427 & i21) | (v2169 & ~i21),
  v3427 = (v2393 & i22) | (v2173 & ~i22),
  v3428 = (v3429 & i21) | (v2208 & ~i21),
  v3429 = (v2411 & i22) | (v2212 & ~i22),
  v3430 = (v3433 & i20) | (v3431 & ~i20),
  v3431 = (v3432 & i21) | (v2169 & ~i21),
  v3432 = (v2430 & i22) | (v2173 & ~i22),
  v3433 = (v3434 & i21) | (v2208 & ~i21),
  v3434 = (v2430 & i22) | (v2212 & ~i22),
  v3435 = (v3459 & i16) | (v3436 & ~i16),
  v3436 = (v3448 & i17) | (v3437 & ~i17),
  v3437 = (v3443 & i19) | (v3438 & ~i19),
  v3438 = (v3441 & i20) | (v3439 & ~i20),
  v3439 = (v3440 & i21) | (v2169 & ~i21),
  v3440 = (v2448 & i22) | (v2173 & ~i22),
  v3441 = (v3442 & i21) | (v2208 & ~i21),
  v3442 = (v2458 & i22) | (v2212 & ~i22),
  v3443 = (v3446 & i20) | (v3444 & ~i20),
  v3444 = (v3445 & i21) | (v2169 & ~i21),
  v3445 = (v2469 & i22) | (v2173 & ~i22),
  v3446 = (v3447 & i21) | (v2208 & ~i21),
  v3447 = (v2478 & i22) | (v2212 & ~i22),
  v3448 = (v3454 & i19) | (v3449 & ~i19),
  v3449 = (v3452 & i20) | (v3450 & ~i20),
  v3450 = (v3451 & i21) | (v2169 & ~i21),
  v3451 = (v2489 & i22) | (v2173 & ~i22),
  v3452 = (v3453 & i21) | (v2208 & ~i21),
  v3453 = (v2498 & i22) | (v2212 & ~i22),
  v3454 = (v3457 & i20) | (v3455 & ~i20),
  v3455 = (v3456 & i21) | (v2169 & ~i21),
  v3456 = (v2508 & i22) | (v2173 & ~i22),
  v3457 = (v3458 & i21) | (v2208 & ~i21),
  v3458 = (v2508 & i22) | (v2212 & ~i22),
  v3459 = (v3471 & i17) | (v3460 & ~i17),
  v3460 = (v3466 & i19) | (v3461 & ~i19),
  v3461 = (v3464 & i20) | (v3462 & ~i20),
  v3462 = (v3463 & i21) | (v2169 & ~i21),
  v3463 = (v2520 & i22) | (v2173 & ~i22),
  v3464 = (v3465 & i21) | (v2208 & ~i21),
  v3465 = (v2530 & i22) | (v2212 & ~i22),
  v3466 = (v3469 & i20) | (v3467 & ~i20),
  v3467 = (v3468 & i21) | (v2169 & ~i21),
  v3468 = (v2541 & i22) | (v2173 & ~i22),
  v3469 = (v3470 & i21) | (v2208 & ~i21),
  v3470 = (v2550 & i22) | (v2212 & ~i22),
  v3471 = (v3477 & i19) | (v3472 & ~i19),
  v3472 = (v3475 & i20) | (v3473 & ~i20),
  v3473 = (v3474 & i21) | (v2169 & ~i21),
  v3474 = (v2561 & i22) | (v2173 & ~i22),
  v3475 = (v3476 & i21) | (v2208 & ~i21),
  v3476 = (v2570 & i22) | (v2212 & ~i22),
  v3477 = (v3480 & i20) | (v3478 & ~i20),
  v3478 = (v3479 & i21) | (v2169 & ~i21),
  v3479 = (v2580 & i22) | (v2173 & ~i22),
  v3480 = (v3481 & i21) | (v2208 & ~i21),
  v3481 = (v2580 & i22) | (v2212 & ~i22),
  v3482 = (v3530 & i15) | (v3483 & ~i15),
  v3483 = (v3507 & i16) | (v3484 & ~i16),
  v3484 = (v3496 & i17) | (v3485 & ~i17),
  v3485 = (v3491 & i19) | (v3486 & ~i19),
  v3486 = (v3489 & i20) | (v3487 & ~i20),
  v3487 = (v3488 & i21) | (v2169 & ~i21),
  v3488 = (v2605 & i22) | (v2173 & ~i22),
  v3489 = (v3490 & i21) | (v2208 & ~i21),
  v3490 = (v2627 & i22) | (v2212 & ~i22),
  v3491 = (v3494 & i20) | (v3492 & ~i20),
  v3492 = (v3493 & i21) | (v2169 & ~i21),
  v3493 = (v2655 & i22) | (v2173 & ~i22),
  v3494 = (v3495 & i21) | (v2208 & ~i21),
  v3495 = (v2679 & i22) | (v2212 & ~i22),
  v3496 = (v3502 & i19) | (v3497 & ~i19),
  v3497 = (v3500 & i20) | (v3498 & ~i20),
  v3498 = (v3499 & i21) | (v2169 & ~i21),
  v3499 = (v2705 & i22) | (v2173 & ~i22),
  v3500 = (v3501 & i21) | (v2208 & ~i21),
  v3501 = (v2729 & i22) | (v2212 & ~i22),
  v3502 = (v3505 & i20) | (v3503 & ~i20),
  v3503 = (v3504 & i21) | (v2169 & ~i21),
  v3504 = (v2748 & i22) | (v2173 & ~i22),
  v3505 = (v3506 & i21) | (v2208 & ~i21),
  v3506 = (v2748 & i22) | (v2212 & ~i22),
  v3507 = (v3519 & i17) | (v3508 & ~i17),
  v3508 = (v3514 & i19) | (v3509 & ~i19),
  v3509 = (v3512 & i20) | (v3510 & ~i20),
  v3510 = (v3511 & i21) | (v2169 & ~i21),
  v3511 = (v2773 & i22) | (v2173 & ~i22),
  v3512 = (v3513 & i21) | (v2208 & ~i21),
  v3513 = (v2793 & i22) | (v2212 & ~i22),
  v3514 = (v3517 & i20) | (v3515 & ~i20),
  v3515 = (v3516 & i21) | (v2169 & ~i21),
  v3516 = (v2818 & i22) | (v2173 & ~i22),
  v3517 = (v3518 & i21) | (v2208 & ~i21),
  v3518 = (v2842 & i22) | (v2212 & ~i22),
  v3519 = (v3525 & i19) | (v3520 & ~i19),
  v3520 = (v3523 & i20) | (v3521 & ~i20),
  v3521 = (v3522 & i21) | (v2169 & ~i21),
  v3522 = (v2868 & i22) | (v2173 & ~i22),
  v3523 = (v3524 & i21) | (v2208 & ~i21),
  v3524 = (v2892 & i22) | (v2212 & ~i22),
  v3525 = (v3528 & i20) | (v3526 & ~i20),
  v3526 = (v3527 & i21) | (v2169 & ~i21),
  v3527 = (v2911 & i22) | (v2173 & ~i22),
  v3528 = (v3529 & i21) | (v2208 & ~i21),
  v3529 = (v2911 & i22) | (v2212 & ~i22),
  v3530 = (v3554 & i16) | (v3531 & ~i16),
  v3531 = (v3543 & i17) | (v3532 & ~i17),
  v3532 = (v3538 & i19) | (v3533 & ~i19),
  v3533 = (v3536 & i20) | (v3534 & ~i20),
  v3534 = (v3535 & i21) | (v2169 & ~i21),
  v3535 = (v2933 & i22) | (v2173 & ~i22),
  v3536 = (v3537 & i21) | (v2208 & ~i21),
  v3537 = (v2949 & i22) | (v2212 & ~i22),
  v3538 = (v3541 & i20) | (v3539 & ~i20),
  v3539 = (v3540 & i21) | (v2169 & ~i21),
  v3540 = (v2965 & i22) | (v2173 & ~i22),
  v3541 = (v3542 & i21) | (v2208 & ~i21),
  v3542 = (v2980 & i22) | (v2212 & ~i22),
  v3543 = (v3549 & i19) | (v3544 & ~i19),
  v3544 = (v3547 & i20) | (v3545 & ~i20),
  v3545 = (v3546 & i21) | (v2169 & ~i21),
  v3546 = (v2997 & i22) | (v2173 & ~i22),
  v3547 = (v3548 & i21) | (v2208 & ~i21),
  v3548 = (v3012 & i22) | (v2212 & ~i22),
  v3549 = (v3552 & i20) | (v3550 & ~i20),
  v3550 = (v3551 & i21) | (v2169 & ~i21),
  v3551 = (v3026 & i22) | (v2173 & ~i22),
  v3552 = (v3553 & i21) | (v2208 & ~i21),
  v3553 = (v3026 & i22) | (v2212 & ~i22),
  v3554 = (v3566 & i17) | (v3555 & ~i17),
  v3555 = (v3561 & i19) | (v3556 & ~i19),
  v3556 = (v3559 & i20) | (v3557 & ~i20),
  v3557 = (v3558 & i21) | (v2169 & ~i21),
  v3558 = (v3047 & i22) | (v2173 & ~i22),
  v3559 = (v3560 & i21) | (v2208 & ~i21),
  v3560 = (v3063 & i22) | (v2212 & ~i22),
  v3561 = (v3564 & i20) | (v3562 & ~i20),
  v3562 = (v3563 & i21) | (v2169 & ~i21),
  v3563 = (v3079 & i22) | (v2173 & ~i22),
  v3564 = (v3565 & i21) | (v2208 & ~i21),
  v3565 = (v3094 & i22) | (v2212 & ~i22),
  v3566 = (v3572 & i19) | (v3567 & ~i19),
  v3567 = (v3570 & i20) | (v3568 & ~i20),
  v3568 = (v3569 & i21) | (v2169 & ~i21),
  v3569 = (v3111 & i22) | (v2173 & ~i22),
  v3570 = (v3571 & i21) | (v2208 & ~i21),
  v3571 = (v3126 & i22) | (v2212 & ~i22),
  v3572 = (v3575 & i20) | (v3573 & ~i20),
  v3573 = (v3574 & i21) | (v2169 & ~i21),
  v3574 = (v3140 & i22) | (v2173 & ~i22),
  v3575 = (v3576 & i21) | (v2208 & ~i21),
  v3576 = (v3140 & i22) | (v2212 & ~i22),
  v3577 = (v3625 & i15) | (v3578 & ~i15),
  v3578 = (v3602 & i16) | (v3579 & ~i16),
  v3579 = (v3591 & i17) | (v3580 & ~i17),
  v3580 = (v3586 & i19) | (v3581 & ~i19),
  v3581 = (v3584 & i20) | (v3582 & ~i20),
  v3582 = (v3583 & i21) | (v2169 & ~i21),
  v3583 = (v3156 & i22) | (v2173 & ~i22),
  v3584 = (v3585 & i21) | (v2208 & ~i21),
  v3585 = (v3163 & i22) | (v2212 & ~i22),
  v3586 = (v3589 & i20) | (v3587 & ~i20),
  v3587 = (v3588 & i21) | (v2169 & ~i21),
  v3588 = (v3171 & i22) | (v2173 & ~i22),
  v3589 = (v3590 & i21) | (v2208 & ~i21),
  v3590 = (v3178 & i22) | (v2212 & ~i22),
  v3591 = (v3597 & i19) | (v3592 & ~i19),
  v3592 = (v3595 & i20) | (v3593 & ~i20),
  v3593 = (v3594 & i21) | (v2169 & ~i21),
  v3594 = (v3187 & i22) | (v2173 & ~i22),
  v3595 = (v3596 & i21) | (v2208 & ~i21),
  v3596 = (v3194 & i22) | (v2212 & ~i22),
  v3597 = (v3600 & i20) | (v3598 & ~i20),
  v3598 = (v3599 & i21) | (v2169 & ~i21),
  v3599 = (v3202 & i22) | (v2173 & ~i22),
  v3600 = (v3601 & i21) | (v2208 & ~i21),
  v3601 = (v3202 & i22) | (v2212 & ~i22),
  v3602 = (v3614 & i17) | (v3603 & ~i17),
  v3603 = (v3609 & i19) | (v3604 & ~i19),
  v3604 = (v3607 & i20) | (v3605 & ~i20),
  v3605 = (v3606 & i21) | (v2169 & ~i21),
  v3606 = (v3214 & i22) | (v2173 & ~i22),
  v3607 = (v3608 & i21) | (v2208 & ~i21),
  v3608 = (v3221 & i22) | (v2212 & ~i22),
  v3609 = (v3612 & i20) | (v3610 & ~i20),
  v3610 = (v3611 & i21) | (v2169 & ~i21),
  v3611 = (v3229 & i22) | (v2173 & ~i22),
  v3612 = (v3613 & i21) | (v2208 & ~i21),
  v3613 = (v3236 & i22) | (v2212 & ~i22),
  v3614 = (v3620 & i19) | (v3615 & ~i19),
  v3615 = (v3618 & i20) | (v3616 & ~i20),
  v3616 = (v3617 & i21) | (v2169 & ~i21),
  v3617 = (v3245 & i22) | (v2173 & ~i22),
  v3618 = (v3619 & i21) | (v2208 & ~i21),
  v3619 = (v3252 & i22) | (v2212 & ~i22),
  v3620 = (v3623 & i20) | (v3621 & ~i20),
  v3621 = (v3622 & i21) | (v2169 & ~i21),
  v3622 = (v3260 & i22) | (v2173 & ~i22),
  v3623 = (v3624 & i21) | (v2208 & ~i21),
  v3624 = (v3260 & i22) | (v2212 & ~i22),
  v3625 = (v3649 & i16) | (v3626 & ~i16),
  v3626 = (v3638 & i17) | (v3627 & ~i17),
  v3627 = (v3633 & i19) | (v3628 & ~i19),
  v3628 = (v3631 & i20) | (v3629 & ~i20),
  v3629 = (v3630 & i21) | (v2169 & ~i21),
  v3630 = (v3273 & i22) | (v2173 & ~i22),
  v3631 = (v3632 & i21) | (v2208 & ~i21),
  v3632 = (v3280 & i22) | (v2212 & ~i22),
  v3633 = (v3636 & i20) | (v3634 & ~i20),
  v3634 = (v3635 & i21) | (v2169 & ~i21),
  v3635 = (v3288 & i22) | (v2173 & ~i22),
  v3636 = (v3637 & i21) | (v2208 & ~i21),
  v3637 = (v3295 & i22) | (v2212 & ~i22),
  v3638 = (v3644 & i19) | (v3639 & ~i19),
  v3639 = (v3642 & i20) | (v3640 & ~i20),
  v3640 = (v3641 & i21) | (v2169 & ~i21),
  v3641 = (v3304 & i22) | (v2173 & ~i22),
  v3642 = (v3643 & i21) | (v2208 & ~i21),
  v3643 = (v3311 & i22) | (v2212 & ~i22),
  v3644 = (v3647 & i20) | (v3645 & ~i20),
  v3645 = (v3646 & i21) | (v2169 & ~i21),
  v3646 = (v3319 & i22) | (v2173 & ~i22),
  v3647 = (v3648 & i21) | (v2208 & ~i21),
  v3648 = (v3319 & i22) | (v2212 & ~i22),
  v3649 = (v3661 & i17) | (v3650 & ~i17),
  v3650 = (v3656 & i19) | (v3651 & ~i19),
  v3651 = (v3654 & i20) | (v3652 & ~i20),
  v3652 = (v3653 & i21) | (v2169 & ~i21),
  v3653 = (v3331 & i22) | (v2173 & ~i22),
  v3654 = (v3655 & i21) | (v2208 & ~i21),
  v3655 = (v3338 & i22) | (v2212 & ~i22),
  v3656 = (v3659 & i20) | (v3657 & ~i20),
  v3657 = (v3658 & i21) | (v2169 & ~i21),
  v3658 = (v3346 & i22) | (v2173 & ~i22),
  v3659 = (v3660 & i21) | (v2208 & ~i21),
  v3660 = (v3353 & i22) | (v2212 & ~i22),
  v3661 = (v3667 & i19) | (v3662 & ~i19),
  v3662 = (v3665 & i20) | (v3663 & ~i20),
  v3663 = (v3664 & i21) | (v2169 & ~i21),
  v3664 = (v3362 & i22) | (v2173 & ~i22),
  v3665 = (v3666 & i21) | (v2208 & ~i21),
  v3666 = (v3369 & i22) | (v2212 & ~i22),
  v3667 = (v3670 & i20) | (v3668 & ~i20),
  v3668 = (v3669 & i21) | (v2169 & ~i21),
  v3669 = (v3377 & i22) | (v2173 & ~i22),
  v3670 = (v3671 & i21) | (v2208 & ~i21),
  v3671 = (v3377 & i22) | (v2212 & ~i22),
  v3672 = (v3676 & i11) | (v3673 & ~i11),
  v3673 = (v3676 & i12) | (v3674 & ~i12),
  v3674 = (v3676 & i13) | (v3675 & ~i13),
  v3675 = (v3681 & i14) | (v3676 & ~i14),
  v3676 = (v3679 & i20) | (v3677 & ~i20),
  v3677 = (v3678 & i21) | (v2169 & ~i21),
  v3678 = (v2178 & i22) | (v2173 & ~i22),
  v3679 = (v3680 & i21) | (v2208 & ~i21),
  v3680 = (v2178 & i22) | (v2212 & ~i22),
  v3681 = (v3785 & i15) | (v3682 & ~i15),
  v3682 = (v3734 & i16) | (v3683 & ~i16),
  v3683 = (v3711 & i17) | (v3684 & ~i17),
  v3684 = (v3698 & i19) | (v3685 & ~i19),
  v3685 = (v3692 & i20) | (v3686 & ~i20),
  v3686 = (v3687 & i21) | (v2169 & ~i21),
  v3687 = (v3688 & i22) | (v2173 & ~i22),
  v3688 = (v63 & i30) | (v3689 & ~i30),
  v3689 = (v63 & i31) | (v3690 & ~i31),
  v3690 = (v63 & i32) | (v3691 & ~i32),
  v3691 = (v2189 & i33) | (v2609 & ~i33),
  v3692 = (v3693 & i21) | (v2208 & ~i21),
  v3693 = (v3694 & i22) | (v2212 & ~i22),
  v3694 = (v63 & i30) | (v3695 & ~i30),
  v3695 = (v63 & i31) | (v3696 & ~i31),
  v3696 = (v63 & i32) | (v3697 & ~i32),
  v3697 = (v2189 & i33) | (v2631 & ~i33),
  v3698 = (v3705 & i20) | (v3699 & ~i20),
  v3699 = (v3700 & i21) | (v2169 & ~i21),
  v3700 = (v3701 & i22) | (v2173 & ~i22),
  v3701 = (v63 & i30) | (v3702 & ~i30),
  v3702 = (v63 & i31) | (v3703 & ~i31),
  v3703 = (v63 & i32) | (v3704 & ~i32),
  v3704 = (v2189 & i33) | (v2659 & ~i33),
  v3705 = (v3706 & i21) | (v2208 & ~i21),
  v3706 = (v3707 & i22) | (v2212 & ~i22),
  v3707 = (v63 & i30) | (v3708 & ~i30),
  v3708 = (v63 & i31) | (v3709 & ~i31),
  v3709 = (v63 & i32) | (v3710 & ~i32),
  v3710 = (v2189 & i33) | (v2683 & ~i33),
  v3711 = (v3725 & i19) | (v3712 & ~i19),
  v3712 = (v3719 & i20) | (v3713 & ~i20),
  v3713 = (v3714 & i21) | (v2169 & ~i21),
  v3714 = (v3715 & i22) | (v2173 & ~i22),
  v3715 = (v63 & i30) | (v3716 & ~i30),
  v3716 = (v63 & i31) | (v3717 & ~i31),
  v3717 = (v63 & i32) | (v3718 & ~i32),
  v3718 = (v2189 & i33) | (v2709 & ~i33),
  v3719 = (v3720 & i21) | (v2208 & ~i21),
  v3720 = (v3721 & i22) | (v2212 & ~i22),
  v3721 = (v63 & i30) | (v3722 & ~i30),
  v3722 = (v63 & i31) | (v3723 & ~i31),
  v3723 = (v63 & i32) | (v3724 & ~i32),
  v3724 = (v2189 & i33) | (v2733 & ~i33),
  v3725 = (v3732 & i20) | (v3726 & ~i20),
  v3726 = (v3727 & i21) | (v2169 & ~i21),
  v3727 = (v3728 & i22) | (v2173 & ~i22),
  v3728 = (v63 & i30) | (v3729 & ~i30),
  v3729 = (v63 & i31) | (v3730 & ~i31),
  v3730 = (v63 & i32) | (v3731 & ~i32),
  v3731 = (v2189 & i33) | (v2752 & ~i33),
  v3732 = (v3733 & i21) | (v2208 & ~i21),
  v3733 = (v3728 & i22) | (v2212 & ~i22),
  v3734 = (v3762 & i17) | (v3735 & ~i17),
  v3735 = (v3749 & i19) | (v3736 & ~i19),
  v3736 = (v3743 & i20) | (v3737 & ~i20),
  v3737 = (v3738 & i21) | (v2169 & ~i21),
  v3738 = (v3739 & i22) | (v2173 & ~i22),
  v3739 = (v63 & i30) | (v3740 & ~i30),
  v3740 = (v63 & i31) | (v3741 & ~i31),
  v3741 = (v63 & i32) | (v3742 & ~i32),
  v3742 = (v2189 & i33) | (v2777 & ~i33),
  v3743 = (v3744 & i21) | (v2208 & ~i21),
  v3744 = (v3745 & i22) | (v2212 & ~i22),
  v3745 = (v63 & i30) | (v3746 & ~i30),
  v3746 = (v63 & i31) | (v3747 & ~i31),
  v3747 = (v63 & i32) | (v3748 & ~i32),
  v3748 = (v2189 & i33) | (v2797 & ~i33),
  v3749 = (v3756 & i20) | (v3750 & ~i20),
  v3750 = (v3751 & i21) | (v2169 & ~i21),
  v3751 = (v3752 & i22) | (v2173 & ~i22),
  v3752 = (v63 & i30) | (v3753 & ~i30),
  v3753 = (v63 & i31) | (v3754 & ~i31),
  v3754 = (v63 & i32) | (v3755 & ~i32),
  v3755 = (v2189 & i33) | (v2822 & ~i33),
  v3756 = (v3757 & i21) | (v2208 & ~i21),
  v3757 = (v3758 & i22) | (v2212 & ~i22),
  v3758 = (v63 & i30) | (v3759 & ~i30),
  v3759 = (v63 & i31) | (v3760 & ~i31),
  v3760 = (v63 & i32) | (v3761 & ~i32),
  v3761 = (v2189 & i33) | (v2846 & ~i33),
  v3762 = (v3776 & i19) | (v3763 & ~i19),
  v3763 = (v3770 & i20) | (v3764 & ~i20),
  v3764 = (v3765 & i21) | (v2169 & ~i21),
  v3765 = (v3766 & i22) | (v2173 & ~i22),
  v3766 = (v63 & i30) | (v3767 & ~i30),
  v3767 = (v63 & i31) | (v3768 & ~i31),
  v3768 = (v63 & i32) | (v3769 & ~i32),
  v3769 = (v2189 & i33) | (v2872 & ~i33),
  v10000 = (v9301 & i22) | (v9289 & ~i22),
  v10001 = (v10004 & i20) | (v10002 & ~i20),
  v10002 = (v10003 & i21) | (v9312 & ~i21),
  v3770 = (v3771 & i21) | (v2208 & ~i21),
  v10003 = (v9345 & i22) | (v9329 & ~i22),
  v3771 = (v3772 & i22) | (v2212 & ~i22),
  v10004 = (v10005 & i21) | (v9355 & ~i21),
  v3772 = (v63 & i30) | (v3773 & ~i30),
  v10005 = (v9388 & i22) | (v9372 & ~i22),
  v3773 = (v63 & i31) | (v3774 & ~i31),
  v10006 = (v10012 & i19) | (v10007 & ~i19),
  v3774 = (v63 & i32) | (v3775 & ~i32),
  v10007 = (v10010 & i20) | (v10008 & ~i20),
  v3775 = (v2189 & i33) | (v2896 & ~i33),
  v10008 = (v10009 & i21) | (v9400 & ~i21),
  v3776 = (v3783 & i20) | (v3777 & ~i20),
  v10009 = (v9433 & i22) | (v9417 & ~i22),
  v3777 = (v3778 & i21) | (v2169 & ~i21),
  v3778 = (v3779 & i22) | (v2173 & ~i22),
  v3779 = (v63 & i30) | (v3780 & ~i30),
  v10010 = (v10011 & i21) | (v9443 & ~i21),
  v10011 = (v9476 & i22) | (v9460 & ~i22),
  v10012 = (v10013 & i21) | (v9486 & ~i21),
  v3780 = (v63 & i31) | (v3781 & ~i31),
  v10013 = (v9507 & i22) | (v9497 & ~i22),
  v3781 = (v63 & i32) | (v3782 & ~i32),
  v10014 = (v10035 & i16) | (v10015 & ~i16),
  v3782 = (v2189 & i33) | (v2915 & ~i33),
  v10015 = (v10027 & i17) | (v10016 & ~i17),
  v3783 = (v3784 & i21) | (v2208 & ~i21),
  v10016 = (v10022 & i19) | (v10017 & ~i19),
  v3784 = (v3779 & i22) | (v2212 & ~i22),
  v10017 = (v10020 & i20) | (v10018 & ~i20),
  v3785 = (v3837 & i16) | (v3786 & ~i16),
  v10018 = (v10019 & i21) | (v9521 & ~i21),
  v3786 = (v3814 & i17) | (v3787 & ~i17),
  v10019 = (v9538 & i22) | (v9530 & ~i22),
  v3787 = (v3801 & i19) | (v3788 & ~i19),
  v3788 = (v3795 & i20) | (v3789 & ~i20),
  v3789 = (v3790 & i21) | (v2169 & ~i21),
  v10020 = (v10021 & i21) | (v9549 & ~i21),
  v10021 = (v9566 & i22) | (v9558 & ~i22),
  v10022 = (v10025 & i20) | (v10023 & ~i20),
  v3790 = (v3791 & i22) | (v2173 & ~i22),
  v10023 = (v10024 & i21) | (v9578 & ~i21),
  v3791 = (v63 & i30) | (v3792 & ~i30),
  v10024 = (v9593 & i22) | (v9586 & ~i22),
  v3792 = (v63 & i31) | (v3793 & ~i31),
  v10025 = (v10026 & i21) | (v9604 & ~i21),
  v3793 = (v63 & i32) | (v3794 & ~i32),
  v10026 = (v9619 & i22) | (v9612 & ~i22),
  v3794 = (v2189 & i33) | (v2937 & ~i33),
  v10027 = (v10033 & i19) | (v10028 & ~i19),
  v3795 = (v3796 & i21) | (v2208 & ~i21),
  v10028 = (v10031 & i20) | (v10029 & ~i20),
  v3796 = (v3797 & i22) | (v2212 & ~i22),
  v10029 = (v10030 & i21) | (v9632 & ~i21),
  v3797 = (v63 & i30) | (v3798 & ~i30),
  v3798 = (v63 & i31) | (v3799 & ~i31),
  v3799 = (v63 & i32) | (v3800 & ~i32),
  v10030 = (v9647 & i22) | (v9640 & ~i22),
  v10031 = (v10032 & i21) | (v9658 & ~i21),
  v10032 = (v9673 & i22) | (v9666 & ~i22),
  v10033 = (v10034 & i21) | (v9684 & ~i21),
  v10034 = (v9695 & i22) | (v9690 & ~i22),
  v10035 = (v10047 & i17) | (v10036 & ~i17),
  v10036 = (v10042 & i19) | (v10037 & ~i19),
  v10037 = (v10040 & i20) | (v10038 & ~i20),
  v10038 = (v10039 & i21) | (v9708 & ~i21),
  v10039 = (v9725 & i22) | (v9717 & ~i22),
  v10040 = (v10041 & i21) | (v9735 & ~i21),
  v10041 = (v9752 & i22) | (v9744 & ~i22),
  v10042 = (v10045 & i20) | (v10043 & ~i20),
  v10043 = (v10044 & i21) | (v9763 & ~i21),
  v10044 = (v9778 & i22) | (v9771 & ~i22),
  v10045 = (v10046 & i21) | (v9788 & ~i21),
  v10046 = (v9803 & i22) | (v9796 & ~i22),
  v10047 = (v10053 & i19) | (v10048 & ~i19),
  v10048 = (v10051 & i20) | (v10049 & ~i20),
  v10049 = (v10050 & i21) | (v9815 & ~i21),
  v10050 = (v9830 & i22) | (v9823 & ~i22),
  v10051 = (v10052 & i21) | (v9840 & ~i21),
  v10052 = (v9855 & i22) | (v9848 & ~i22),
  v10053 = (v10054 & i21) | (v9865 & ~i21),
  v10054 = (v9876 & i22) | (v9871 & ~i22),
  v10055 = i29,
  v10056 = (v10063 & i2) | (v10057 & ~i2),
  v10057 = (v10063 & i3) | (~v10058 & ~i3),
  v10058 = (v10063 & i11) | (v10059 & ~i11),
  v10059 = (v10064 & i12) | (v10060 & ~i12),
  v10060 = (v10063 & i13) | (v10061 & ~i13),
  v10061 = (v10062 & i14) | ~i14,
  v10062 = v63 & i29,
  v10063 = i14,
  v10064 = (v10063 & i13) | (v10065 & ~i13),
  v10065 = (~v10066 & ~i14) | i14,
  v10066 = (v10067 & ~i26) | i26,
  v10067 = i27,
  v10068 = (v10081 & i2) | (v10069 & ~i2),
  v10069 = (v10081 & i3) | (~v10070 & ~i3),
  v10070 = (v10076 & i11) | (v10071 & ~i11),
  v10071 = (v10074 & i12) | (v10072 & ~i12),
  v10072 = (v10063 & i13) | (~v10073 & ~i13),
  v10073 = v10062 & i14,
  v10074 = (v10063 & i13) | (v10075 & ~i13),
  v10075 = (v10067 & i14) | ~i14,
  v10076 = (v10080 & i12) | (v10077 & ~i12),
  v10077 = (v10063 & i13) | (~v10078 & ~i13),
  v10078 = v10079 & i14,
  v10079 = (v10067 & i26) | ~i26,
  v10080 = (~v10063 & ~i13) | (v10063 & i13),
  v10081 = i13,
  v10082 = (v10090 & i2) | (v10083 & ~i2),
  v10083 = (v10090 & i3) | (~v10084 & ~i3),
  v10084 = (v10089 & i11) | (v10085 & ~i11),
  v10085 = (v10087 & i12) | (~v10086 & ~i12),
  v10086 = v10063 & i13,
  v10087 = (v10063 & i13) | (v10088 & ~i13),
  v10088 = (v10067 & i14) | (~v10066 & ~i14),
  v10089 = (~v10086 & ~i12) | (v10086 & i12),
  v10090 = i12,
  v10091 = (v10098 & i2) | (v10092 & ~i2),
  v10092 = (v10098 & i3) | (~v10093 & ~i3),
  v3800 = (v2189 & i33) | (v2953 & ~i33),
  v10093 = (v10095 & i11) | (~v10094 & ~i11),
  v3801 = (v3808 & i20) | (v3802 & ~i20),
  v10094 = v10086 & i12,
  v3802 = (v3803 & i21) | (v2169 & ~i21),
  v10095 = (v10086 & i12) | (~v10096 & ~i12),
  v3803 = (v3804 & i22) | (v2173 & ~i22),
  v10096 = (v10097 & ~i13) | i13,
  v3804 = (v63 & i30) | (v3805 & ~i30),
  v10097 = (v10079 & i14) | ~i14,
  v3805 = (v63 & i31) | (v3806 & ~i31),
  v10098 = i11,
  v3806 = (v63 & i32) | (v3807 & ~i32),
  v10099 = (v10107 & i2) | (v10100 & ~i2),
  v3807 = (v2189 & i33) | (v2969 & ~i33),
  v3808 = (v3809 & i21) | (v2208 & ~i21),
  v3809 = (v3810 & i22) | (v2212 & ~i22),
  v3810 = (v63 & i30) | (v3811 & ~i30),
  v3811 = (v63 & i31) | (v3812 & ~i31),
  v3812 = (v63 & i32) | (v3813 & ~i32),
  v3813 = (v2189 & i33) | (v2984 & ~i33),
  v3814 = (v3828 & i19) | (v3815 & ~i19),
  v3815 = (v3822 & i20) | (v3816 & ~i20),
  v3816 = (v3817 & i21) | (v2169 & ~i21),
  v3817 = (v3818 & i22) | (v2173 & ~i22),
  v3818 = (v63 & i30) | (v3819 & ~i30),
  v3819 = (v63 & i31) | (v3820 & ~i31),
  v3820 = (v63 & i32) | (v3821 & ~i32),
  v3821 = (v2189 & i33) | (v3001 & ~i33),
  v3822 = (v3823 & i21) | (v2208 & ~i21),
  v3823 = (v3824 & i22) | (v2212 & ~i22),
  v3824 = (v63 & i30) | (v3825 & ~i30),
  v3825 = (v63 & i31) | (v3826 & ~i31),
  v3826 = (v63 & i32) | (v3827 & ~i32),
  v3827 = (v2189 & i33) | (v3016 & ~i33),
  v3828 = (v3835 & i20) | (v3829 & ~i20),
  v3829 = (v3830 & i21) | (v2169 & ~i21),
  v3830 = (v3831 & i22) | (v2173 & ~i22),
  v3831 = (v63 & i30) | (v3832 & ~i30),
  v3832 = (v63 & i31) | (v3833 & ~i31),
  v3833 = (v63 & i32) | (v3834 & ~i32),
  v3834 = (v2189 & i33) | (v3030 & ~i33),
  v3835 = (v3836 & i21) | (v2208 & ~i21),
  v3836 = (v3831 & i22) | (v2212 & ~i22),
  v3837 = (v3865 & i17) | (v3838 & ~i17),
  v3838 = (v3852 & i19) | (v3839 & ~i19),
  v3839 = (v3846 & i20) | (v3840 & ~i20),
  v3840 = (v3841 & i21) | (v2169 & ~i21),
  v3841 = (v3842 & i22) | (v2173 & ~i22),
  v3842 = (v63 & i30) | (v3843 & ~i30),
  v3843 = (v63 & i31) | (v3844 & ~i31),
  v3844 = (v63 & i32) | (v3845 & ~i32),
  v3845 = (v2189 & i33) | (v3051 & ~i33),
  v3846 = (v3847 & i21) | (v2208 & ~i21),
  v3847 = (v3848 & i22) | (v2212 & ~i22),
  v3848 = (v63 & i30) | (v3849 & ~i30),
  v3849 = (v63 & i31) | (v3850 & ~i31),
  v3850 = (v63 & i32) | (v3851 & ~i32),
  v3851 = (v2189 & i33) | (v3067 & ~i33),
  v3852 = (v3859 & i20) | (v3853 & ~i20),
  v3853 = (v3854 & i21) | (v2169 & ~i21),
  v3854 = (v3855 & i22) | (v2173 & ~i22),
  v3855 = (v63 & i30) | (v3856 & ~i30),
  v3856 = (v63 & i31) | (v3857 & ~i31),
  v3857 = (v63 & i32) | (v3858 & ~i32),
  v3858 = (v2189 & i33) | (v3083 & ~i33),
  v3859 = (v3860 & i21) | (v2208 & ~i21),
  v3860 = (v3861 & i22) | (v2212 & ~i22),
  v3861 = (v63 & i30) | (v3862 & ~i30),
  v3862 = (v63 & i31) | (v3863 & ~i31),
  v3863 = (v63 & i32) | (v3864 & ~i32),
  v3864 = (v2189 & i33) | (v3098 & ~i33),
  v3865 = (v3879 & i19) | (v3866 & ~i19),
  v3866 = (v3873 & i20) | (v3867 & ~i20),
  v3867 = (v3868 & i21) | (v2169 & ~i21),
  v3868 = (v3869 & i22) | (v2173 & ~i22),
  v3869 = (v63 & i30) | (v3870 & ~i30),
  v10100 = (v10107 & i3) | (~v10101 & ~i3),
  v10101 = (v10107 & i7) | (v10102 & ~i7),
  v10102 = (v10108 & i8) | (v10103 & ~i8),
  v3870 = (v63 & i31) | (v3871 & ~i31),
  v10103 = (v10107 & i9) | (~v10104 & ~i9),
  v3871 = (v63 & i32) | (v3872 & ~i32),
  v10104 = (v10106 & i10) | (v10105 & ~i10),
  v3872 = (v2189 & i33) | (v3115 & ~i33),
  v10105 = i25,
  v3873 = (v3874 & i21) | (v2208 & ~i21),
  v10106 = (v63 & i29) | ~i29,
  v3874 = (v3875 & i22) | (v2212 & ~i22),
  v10107 = i10,
  v3875 = (v63 & i30) | (v3876 & ~i30),
  v10108 = (v10107 & i9) | (v10109 & ~i9),
  v3876 = (v63 & i31) | (v3877 & ~i31),
  v10109 = (~v10110 & ~i10) | i10,
  v3877 = (v63 & i32) | (v3878 & ~i32),
  v3878 = (v2189 & i33) | (v3130 & ~i33),
  v3879 = (v3886 & i20) | (v3880 & ~i20),
  v10110 = (v10111 & ~i23) | i23,
  v10111 = i24,
  v10112 = (v10125 & i2) | (v10113 & ~i2),
  v3880 = (v3881 & i21) | (v2169 & ~i21),
  v10113 = (v10125 & i3) | (~v10114 & ~i3),
  v3881 = (v3882 & i22) | (v2173 & ~i22),
  v10114 = (v10120 & i7) | (v10115 & ~i7),
  v3882 = (v63 & i30) | (v3883 & ~i30),
  v10115 = (v10118 & i8) | (v10116 & ~i8),
  v3883 = (v63 & i31) | (v3884 & ~i31),
  v10116 = (v10107 & i9) | (v10117 & ~i9),
  v3884 = (v63 & i32) | (v3885 & ~i32),
  v10117 = (v10106 & i10) | ~i10,
  v3885 = (v2189 & i33) | (v3144 & ~i33),
  v10118 = (v10107 & i9) | (v10119 & ~i9),
  v3886 = (v3887 & i21) | (v2208 & ~i21),
  v10119 = (v10111 & i10) | ~i10,
  v3887 = (v3882 & i22) | (v2212 & ~i22),
  v3888 = (v27 & i2) | (v3889 & ~i2),
  v3889 = (v27 & i3) | (v3890 & ~i3),
  v10120 = (v10124 & i8) | (v10121 & ~i8),
  v10121 = (v10107 & i9) | (~v10122 & ~i9),
  v10122 = v10123 & i10,
  v3890 = (v4918 & i4) | (v3891 & ~i4),
  v10123 = (v10111 & i23) | ~i23,
  v3891 = (v4918 & i5) | (v3892 & ~i5),
  v10124 = (~v10107 & ~i9) | (v10107 & i9),
  v3892 = (v4918 & i6) | (v3893 & ~i6),
  v10125 = i9,
  v3893 = (v4829 & i7) | (v3894 & ~i7),
  v10126 = (v10134 & i2) | (v10127 & ~i2),
  v3894 = (v4829 & i8) | (v3895 & ~i8),
  v10127 = (v10134 & i3) | (~v10128 & ~i3),
  v3895 = (v4829 & i9) | (v3896 & ~i9),
  v10128 = (v10133 & i7) | (v10129 & ~i7),
  v3896 = (v4519 & i10) | (v3897 & ~i10),
  v10129 = (v10131 & i8) | (~v10130 & ~i8),
  v3897 = (v3901 & i11) | (v3898 & ~i11),
  v3898 = (v3901 & i12) | (v3899 & ~i12),
  v3899 = (v3901 & i13) | (v3900 & ~i13),
  v10130 = v10107 & i9,
  v10131 = (v10107 & i9) | (v10132 & ~i9),
  v10132 = (v10111 & i10) | (~v10110 & ~i10),
  v10133 = (~v10130 & ~i8) | (v10130 & i8),
  v10134 = i8,
  v10135 = (v10142 & i2) | (v10136 & ~i2),
  v10136 = (v10142 & i3) | (~v10137 & ~i3),
  v10137 = (v10139 & i7) | (~v10138 & ~i7),
  v10138 = v10130 & i8,
  v10139 = (v10130 & i8) | (~v10140 & ~i8),
  v10140 = (v10141 & ~i9) | i9,
  v10141 = (v10123 & i10) | ~i10,
  v10142 = i7,
  v10143 = (v10246 & i2) | (~v10144 & ~i2),
  v10144 = (v10239 & i3) | (~v10145 & ~i3),
  v10145 = (v10231 & i6) | (~v10146 & ~i6),
  v10146 = (v10214 & i7) | (v10147 & ~i7),
  v10147 = (v10179 & i8) | (v10148 & ~i8),
  v10148 = (v10163 & i9) | (v10149 & ~i9),
  v10149 = (v10159 & i11) | (v10150 & ~i11),
  v10150 = (v10154 & i12) | (v10151 & ~i12),
  v10151 = (v10152 & i13) | ~i13,
  v10152 = (v10153 & i14) | ~i14,
  v10153 = (v7448 & i30) | ~i30,
  v10154 = (v10153 & i13) | (v10155 & ~i13),
  v10155 = (v10158 & i14) | (v10156 & ~i14),
  v10156 = (v10153 & i26) | (v10157 & ~i26),
  v10157 = (v10153 & i27) | ~i27,
  v10158 = (v10153 & ~i27) | i27,
  v10159 = (v10153 & i12) | (v10160 & ~i12),
  v10160 = (v10153 & i13) | (v10161 & ~i13),
  v10161 = (v10162 & i14) | (v10153 & ~i14),
  v10162 = (v10157 & i26) | (v10153 & ~i26),
  v10163 = (v10164 & i10) | (v10149 & ~i10),
  v10164 = (v10175 & i11) | (v10165 & ~i11),
  v10165 = (v10170 & i12) | (v10166 & ~i12),
  v10166 = (v10168 & i13) | (v10167 & ~i13),
  v10167 = (v8373 & i30) | ~i30,
  v10168 = (v10169 & i14) | (v10167 & ~i14),
  v10169 = (v6430 & i30) | ~i30,
  v10170 = (v10169 & i13) | (v10171 & ~i13),
  v10171 = (v10174 & i14) | (v10172 & ~i14),
  v10172 = (v10169 & i26) | (v10173 & ~i26),
  v10173 = (v10169 & i27) | (v10167 & ~i27),
  v10174 = (v10167 & i27) | (v10169 & ~i27),
  v10175 = (v10169 & i12) | (v10176 & ~i12),
  v10176 = (v10169 & i13) | (v10177 & ~i13),
  v10177 = (v10178 & i14) | (v10169 & ~i14),
  v10178 = (v10173 & i26) | (v10169 & ~i26),
  v10179 = (v10164 & i9) | (v10180 & ~i9),
  v10180 = (v10200 & i10) | (v10181 & ~i10),
  v10181 = (v10195 & i11) | (v10182 & ~i11),
  v10182 = (v10189 & i12) | (v10183 & ~i12),
  v10183 = (v10186 & i13) | (v10184 & ~i13),
  v10184 = (v10167 & i23) | (v10185 & ~i23),
  v10185 = (v10167 & i24) | ~i24,
  v10186 = (v10187 & i14) | (v10184 & ~i14),
  v10187 = (v10169 & i23) | (v10188 & ~i23),
  v10188 = (v10169 & i24) | (v10153 & ~i24),
  v10189 = (v10187 & i13) | (v10190 & ~i13),
  v10190 = (v10193 & i14) | (v10191 & ~i14),
  v10191 = (v10172 & i23) | (v10192 & ~i23),
  v10192 = (v10172 & i24) | (v10156 & ~i24),
  v3900 = (v4268 & i14) | (v3901 & ~i14),
  v10193 = (v10174 & i23) | (v10194 & ~i23),
  v3901 = (v4143 & i15) | (v3902 & ~i15),
  v10194 = (v10174 & i24) | (v10158 & ~i24),
  v3902 = (v4032 & i16) | (v3903 & ~i16),
  v10195 = (v10187 & i12) | (v10196 & ~i12),
  v3903 = (v3985 & i17) | (v3904 & ~i17),
  v10196 = (v10187 & i13) | (v10197 & ~i13),
  v3904 = (v3949 & i19) | (v3905 & ~i19),
  v10197 = (v10198 & i14) | (v10187 & ~i14),
  v3905 = (v3933 & i20) | (v3906 & ~i20),
  v10198 = (v10178 & i23) | (v10199 & ~i23),
  v3906 = (v3907 & i21) | (v27 & ~i21),
  v10199 = (v10178 & i24) | (v10162 & ~i24),
  v3907 = (v3911 & i22) | (v3908 & ~i22),
  v3908 = (v27 & i30) | (v3909 & ~i30),
  v3909 = (v27 & i31) | (v3910 & ~i31),
  v3910 = (~v49 & ~i32) | i32,
  v3911 = (v3920 & i25) | (v3912 & ~i25),
  v3912 = (v27 & i30) | (v3913 & ~i30),
  v3913 = (v27 & i31) | (v3914 & ~i31),
  v3914 = (~v3915 & ~i32) | i32,
  v3915 = (v3919 & i37) | (v3916 & ~i37),
  v3916 = (v3918 & i42) | (v3917 & ~i42),
  v3917 = (~v20 & ~i45) | i45,
  v3918 = (v3917 & i43) | (v49 & ~i43),
  v3919 = (v3916 & i38) | (v3917 & ~i38),
  v3920 = (v27 & i30) | (v3921 & ~i30),
  v3921 = (v27 & i31) | (v3922 & ~i31),
  v3922 = (~v3923 & ~i32) | i32,
  v3923 = (v3932 & i36) | (v3924 & ~i36),
  v3924 = (v3931 & i37) | (v3925 & ~i37),
  v3925 = (v3927 & i38) | (v3926 & ~i38),
  v3926 = (v3916 & i39) | (v3927 & ~i39),
  v3927 = (v3916 & i41) | (v3928 & ~i41),
  v3928 = (v3918 & i42) | (v3929 & ~i42),
  v3929 = (v3917 & i43) | (v3930 & ~i43),
  v3930 = (v49 & i44) | (v3917 & ~i44),
  v3931 = (v3927 & i38) | (v3917 & ~i38),
  v3932 = (v3931 & i37) | (v3927 & ~i37),
  v3933 = (v3934 & i21) | (v27 & ~i21),
  v3934 = (v3935 & i22) | (v3908 & ~i22),
  v3935 = (v3936 & i25) | (v3912 & ~i25),
  v3936 = (v27 & i30) | (v3937 & ~i30),
  v3937 = (v27 & i31) | (v3938 & ~i31),
  v3938 = (~v3939 & ~i32) | i32,
  v3939 = (v3948 & i36) | (v3940 & ~i36),
  v3940 = (v3947 & i37) | (v3941 & ~i37),
  v3941 = (v3943 & i38) | (v3942 & ~i38),
  v3942 = (v3943 & i39) | (v3916 & ~i39),
  v3943 = (v3916 & i41) | (v3944 & ~i41),
  v3944 = (v3918 & i42) | (v3945 & ~i42),
  v3945 = (v3917 & i43) | (v3946 & ~i43),
  v3946 = (v3917 & i44) | (v49 & ~i44),
  v3947 = (v3943 & i38) | (v3917 & ~i38),
  v3948 = (v3947 & i37) | (v3943 & ~i37),
  v3949 = (v3968 & i20) | (v3950 & ~i20),
  v3950 = (v3951 & i21) | (v27 & ~i21),
  v3951 = (v3952 & i22) | (v3908 & ~i22),
  v3952 = (v3953 & i25) | (v3912 & ~i25),
  v3953 = (v27 & i30) | (v3954 & ~i30),
  v3954 = (v27 & i31) | (v3955 & ~i31),
  v3955 = (~v3956 & ~i32) | i32,
  v3956 = (v3964 & i35) | (v3957 & ~i35),
  v3957 = (v3963 & i36) | (v3958 & ~i36),
  v3958 = (v3962 & i37) | (v3959 & ~i37),
  v3959 = (v3960 & i38) | (v3916 & ~i38),
  v3960 = (v3927 & i40) | (v3961 & ~i40),
  v3961 = (v3916 & i41) | (v3918 & ~i41),
  v3962 = (v3960 & i38) | (v3917 & ~i38),
  v3963 = (v3962 & i37) | (v3960 & ~i37),
  v3964 = (v3963 & i36) | (v3965 & ~i36),
  v3965 = (v3962 & i37) | (v3966 & ~i37),
  v3966 = (v3960 & i38) | (v3967 & ~i38),
  v3967 = (v3916 & i39) | (v3960 & ~i39),
  v3968 = (v3969 & i21) | (v27 & ~i21),
  v3969 = (v3970 & i22) | (v3908 & ~i22),
  v10200 = (v10210 & i11) | (v10201 & ~i11),
  v10201 = (v10206 & i12) | (v10202 & ~i12),
  v10202 = (v10204 & i13) | (v10203 & ~i13),
  v3970 = (v3971 & i25) | (v3912 & ~i25),
  v10203 = (v10167 & ~i24) | i24,
  v3971 = (v27 & i30) | (v3972 & ~i30),
  v10204 = (v10205 & i14) | (v10203 & ~i14),
  v3972 = (v27 & i31) | (v3973 & ~i31),
  v10205 = (v10153 & i24) | (v10169 & ~i24),
  v3973 = (~v3974 & ~i32) | i32,
  v10206 = (v10205 & i13) | (v10207 & ~i13),
  v3974 = (v3981 & i35) | (v3975 & ~i35),
  v10207 = (v10209 & i14) | (v10208 & ~i14),
  v3975 = (v3980 & i36) | (v3976 & ~i36),
  v10208 = (v10156 & i24) | (v10172 & ~i24),
  v3976 = (v3979 & i37) | (v3977 & ~i37),
  v10209 = (v10158 & i24) | (v10174 & ~i24),
  v3977 = (v3978 & i38) | (v3916 & ~i38),
  v3978 = (v3943 & i40) | (v3961 & ~i40),
  v3979 = (v3978 & i38) | (v3917 & ~i38),
  v10210 = (v10205 & i12) | (v10211 & ~i12),
  v10211 = (v10205 & i13) | (v10212 & ~i13),
  v10212 = (v10213 & i14) | (v10205 & ~i14),
  v3980 = (v3979 & i37) | (v3978 & ~i37),
  v10213 = (v10162 & i24) | (v10178 & ~i24),
  v3981 = (v3980 & i36) | (v3982 & ~i36),
  v10214 = (v10164 & i8) | (v10215 & ~i8),
  v3982 = (v3979 & i37) | (v3983 & ~i37),
  v10215 = (v10164 & i9) | (v10216 & ~i9),
  v3983 = (v3978 & i38) | (v3984 & ~i38),
  v10216 = (v10217 & i10) | (v10164 & ~i10),
  v3984 = (v3978 & i39) | (v3916 & ~i39),
  v10217 = (v10227 & i11) | (v10218 & ~i11),
  v3985 = (v4021 & i19) | (v3986 & ~i19),
  v10218 = (v10223 & i12) | (v10219 & ~i12),
  v3986 = (v4004 & i20) | (v3987 & ~i20),
  v10219 = (v10221 & i13) | (v10220 & ~i13),
  v3987 = (v3988 & i21) | (v27 & ~i21),
  v3988 = (v3989 & i22) | (v3908 & ~i22),
  v3989 = (v3990 & i25) | (v3912 & ~i25),
  v10220 = (v10185 & i23) | (v10167 & ~i23),
  v10221 = (v10222 & i14) | (v10220 & ~i14),
  v10222 = (v10188 & i23) | (v10169 & ~i23),
  v3990 = (v27 & i30) | (v3991 & ~i30),
  v10223 = (v10222 & i13) | (v10224 & ~i13),
  v3991 = (v27 & i31) | (v3992 & ~i31),
  v10224 = (v10226 & i14) | (v10225 & ~i14),
  v3992 = (~v3993 & ~i32) | i32,
  v10225 = (v10192 & i23) | (v10172 & ~i23),
  v3993 = (v4001 & i35) | (v3994 & ~i35),
  v10226 = (v10194 & i23) | (v10174 & ~i23),
  v3994 = (v4000 & i36) | (v3995 & ~i36),
  v10227 = (v10222 & i12) | (v10228 & ~i12),
  v3995 = (v3999 & i37) | (v3996 & ~i37),
  v10228 = (v10222 & i13) | (v10229 & ~i13),
  v3996 = (v3998 & i38) | (v3997 & ~i38),
  v10229 = (v10230 & i14) | (v10222 & ~i14),
  v3997 = (v3916 & i39) | (v3998 & ~i39),
  v3998 = (v3961 & i40) | (v3927 & ~i40),
  v3999 = (v3998 & i38) | (v3917 & ~i38),
  v10230 = (v10199 & i23) | (v10178 & ~i23),
  v10231 = (v10237 & i7) | (v10232 & ~i7),
  v10232 = (v10237 & i8) | (v10233 & ~i8),
  v10233 = (v10236 & i9) | (v10234 & ~i9),
  v10234 = (v10153 & i11) | (v10235 & ~i11),
  v10235 = (v10153 & i12) | (v10151 & ~i12),
  v10236 = (v10237 & i10) | (v10234 & ~i10),
  v10237 = (v10169 & i11) | (v10238 & ~i11),
  v10238 = (v10169 & i12) | (v10166 & ~i12),
  v10239 = (v10241 & i4) | (v10240 & ~i4),
  v10240 = (v10242 & i5) | (v10241 & ~i5),
  v10241 = (~v6430 & ~i6) | (v6430 & i6),
  v10242 = (v6430 & i6) | (~v10243 & ~i6),
  v10243 = (v10244 & i30) | (v6430 & ~i30),
  v10244 = v10245 & i31,
  v10245 = (v254 & i32) | (v510 & ~i32),
  v10246 = i6,
  v10247 = (v10315 & i2) | (~v10248 & ~i2),
  v10248 = (v10305 & i3) | (~v10249 & ~i3),
  v10249 = (v10251 & i5) | (~v10250 & ~i5),
  v10250 = (v10146 & i6) | ~i6,
  v10251 = (v10231 & i6) | (v10252 & ~i6),
  v10252 = (v10291 & i7) | (v10253 & ~i7),
  v10253 = (v10263 & i8) | (v10254 & ~i8),
  v10254 = (v10259 & i11) | (v10255 & ~i11),
  v10255 = (v10256 & i12) | ~i12,
  v10256 = (v10257 & ~i13) | i13,
  v10257 = (v10157 & i14) | (v10258 & ~i14),
  v10258 = (v10158 & ~i26) | i26,
  v10259 = (v10260 & ~i12) | i12,
  v10260 = (v10261 & ~i13) | i13,
  v10261 = (v10262 & i14) | ~i14,
  v10262 = (v10158 & i26) | ~i26,
  v10263 = (v10254 & i9) | (v10264 & ~i9),
  v10264 = (v10281 & i10) | (v10265 & ~i10),
  v10265 = (v10275 & i11) | (v10266 & ~i11),
  v10266 = (v10268 & i12) | (v10267 & ~i12),
  v10267 = (v10203 & ~i23) | i23,
  v10268 = (v10267 & i13) | (v10269 & ~i13),
  v10269 = (v10273 & i14) | (v10270 & ~i14),
  v10270 = (v10258 & i23) | (v10271 & ~i23),
  v10271 = (v10258 & i24) | (v10272 & ~i24),
  v10272 = (v10167 & i26) | (v10174 & ~i26),
  v10273 = (v10157 & i23) | (v10274 & ~i23),
  v10274 = (v10157 & i24) | (v10173 & ~i24),
  v10275 = (v10267 & i12) | (v10276 & ~i12),
  v10276 = (v10267 & i13) | (v10277 & ~i13),
  v10277 = (v10278 & i14) | (v10267 & ~i14),
  v10278 = (v10262 & i23) | (v10279 & ~i23),
  v10279 = (v10262 & i24) | (v10280 & ~i24),
  v10280 = (v10174 & i26) | (v10167 & ~i26),
  v10281 = (v10287 & i11) | (v10282 & ~i11),
  v10282 = (v10283 & i12) | (v10185 & ~i12),
  v10283 = (v10185 & i13) | (v10284 & ~i13),
  v10284 = (v10286 & i14) | (v10285 & ~i14),
  v10285 = (v10272 & i24) | (v10258 & ~i24),
  v10286 = (v10173 & i24) | (v10157 & ~i24),
  v10287 = (v10185 & i12) | (v10288 & ~i12),
  v10288 = (v10185 & i13) | (v10289 & ~i13),
  v10289 = (v10290 & i14) | (v10185 & ~i14),
  v10290 = (v10280 & i24) | (v10262 & ~i24),
  v10291 = (v10254 & i8) | (v10292 & ~i8),
  v10292 = (v10254 & i9) | (v10293 & ~i9),
  v10293 = (v10294 & i10) | (v10254 & ~i10),
  v10294 = (v10301 & i11) | (v10295 & ~i11),
  v10295 = (v10297 & i12) | (v10296 & ~i12),
  v10296 = (v10203 & i23) | ~i23,
  v10297 = (v10296 & i13) | (v10298 & ~i13),
  v10298 = (v10300 & i14) | (v10299 & ~i14),
  v10299 = (v10271 & i23) | (v10258 & ~i23),
  v10300 = (v10274 & i23) | (v10157 & ~i23),
  v10301 = (v10296 & i12) | (v10302 & ~i12),
  v10302 = (v10296 & i13) | (v10303 & ~i13),
  v10303 = (v10304 & i14) | (v10296 & ~i14),
  v10304 = (v10279 & i23) | (v10262 & ~i23),
  v10305 = (v10311 & i4) | (v10306 & ~i4),
  v10306 = (v10308 & i5) | (~v10307 & ~i5),
  v10307 = v8608 & i6,
  v10308 = (v6430 & i6) | (~v10309 & ~i6),
  v10309 = (v10310 & i30) | ~i30,
  v10310 = (v10245 & i31) | ~i31,
  v10311 = (v10314 & i5) | (v10312 & ~i5),
  v10312 = (v10313 & i6) | ~i6,
  v10313 = (v10310 & i30) | (~v6430 & ~i30),
  v10314 = v6430 & i6,
  v10315 = i5,
  v10316 = (v10326 & i2) | (~v10317 & ~i2),
  v10317 = (v10321 & i3) | (~v10318 & ~i3),
  v10318 = (v10320 & i4) | (~v10319 & ~i4),
  v10319 = (v10250 & i5) | ~i5,
  v10320 = (v10251 & i5) | (v10252 & ~i5),
  v10321 = (v10323 & i4) | (~v10322 & ~i4),
  v10322 = v10314 & i5,
  v10323 = (v10314 & i5) | (v10324 & ~i5),
  v10324 = v10325 & i6,
  v10325 = v10244 & i30,
  v10326 = i4,
  v10327 = (v10328 & ~i2) | i2,
  v10328 = i3,
  v10329 = (~v10328 & ~i2) | i2,
  v4000 = (v3999 & i37) | (v3998 & ~i37),
  v4001 = (v4000 & i36) | (v4002 & ~i36),
  v4002 = (v3999 & i37) | (v4003 & ~i37),
  v4003 = (v3998 & i38) | (v3916 & ~i38),
  v4004 = (v4005 & i21) | (v27 & ~i21),
  v4005 = (v4006 & i22) | (v3908 & ~i22),
  v4006 = (v4007 & i25) | (v3912 & ~i25),
  v4007 = (v27 & i30) | (v4008 & ~i30),
  v4008 = (v27 & i31) | (v4009 & ~i31),
  v4009 = (~v4010 & ~i32) | i32,
  v4010 = (v4018 & i35) | (v4011 & ~i35),
  v4011 = (v4017 & i36) | (v4012 & ~i36),
  v4012 = (v4016 & i37) | (v4013 & ~i37),
  v4013 = (v4015 & i38) | (v4014 & ~i38),
  v4014 = (v4015 & i39) | (v3916 & ~i39),
  v4015 = (v3961 & i40) | (v3943 & ~i40),
  v4016 = (v4015 & i38) | (v3917 & ~i38),
  v4017 = (v4016 & i37) | (v4015 & ~i37),
  v4018 = (v4017 & i36) | (v4019 & ~i36),
  v4019 = (v4016 & i37) | (v4020 & ~i37),
  v4020 = (v4015 & i38) | (v3916 & ~i38),
  v4021 = (v4022 & i21) | (v27 & ~i21),
  v4022 = (v4023 & i22) | (v3908 & ~i22),
  v4023 = (v4024 & i25) | (v3912 & ~i25),
  v4024 = (v27 & i30) | (v4025 & ~i30),
  v4025 = (v27 & i31) | (v4026 & ~i31),
  v4026 = (~v4027 & ~i32) | i32,
  v4027 = (v4031 & i36) | (v4028 & ~i36),
  v4028 = (v4030 & i37) | (v4029 & ~i37),
  v4029 = (v3961 & i38) | (v3916 & ~i38),
  v4030 = (v3961 & i38) | (v3917 & ~i38),
  v4031 = (v4030 & i37) | (v3961 & ~i37),
  v4032 = (v4096 & i17) | (v4033 & ~i17),
  v4033 = (v4061 & i19) | (v4034 & ~i19),
  v4034 = (v4048 & i20) | (v4035 & ~i20),
  v4035 = (v4036 & i21) | (v27 & ~i21),
  v4036 = (v4037 & i22) | (v3908 & ~i22),
  v4037 = (v4038 & i25) | (v3912 & ~i25),
  v4038 = (v27 & i30) | (v4039 & ~i30),
  v4039 = (v27 & i31) | (v4040 & ~i31),
  v4040 = (~v4041 & ~i32) | i32,
  v4041 = (v4047 & i36) | (v4042 & ~i36),
  v4042 = (v4046 & i37) | (v4043 & ~i37),
  v4043 = (v4045 & i38) | (v4044 & ~i38),
  v4044 = (v3916 & i39) | (v4045 & ~i39),
  v4045 = (v3918 & i41) | (v3928 & ~i41),
  v4046 = (v4045 & i38) | (v3917 & ~i38),
  v4047 = (v4046 & i37) | (v4045 & ~i37),
  v4048 = (v4049 & i21) | (v27 & ~i21),
  v4049 = (v4050 & i22) | (v3908 & ~i22),
  v4050 = (v4051 & i25) | (v3912 & ~i25),
  v4051 = (v27 & i30) | (v4052 & ~i30),
  v4052 = (v27 & i31) | (v4053 & ~i31),
  v4053 = (~v4054 & ~i32) | i32,
  v4054 = (v4060 & i36) | (v4055 & ~i36),
  v4055 = (v4059 & i37) | (v4056 & ~i37),
  v4056 = (v4058 & i38) | (v4057 & ~i38),
  v4057 = (v4058 & i39) | (v3916 & ~i39),
  \*clm_clk_ctl_time0  = ~v10329,
  v4058 = (v3918 & i41) | (v3944 & ~i41),
  \*clm_clk_ctl_time1  = ~v10327,
  v4059 = (v4058 & i38) | (v3917 & ~i38),
  v4060 = (v4059 & i37) | (v4058 & ~i37),
  v4061 = (v4079 & i20) | (v4062 & ~i20),
  v4062 = (v4063 & i21) | (v27 & ~i21),
  v4063 = (v4064 & i22) | (v3908 & ~i22),
  v4064 = (v4065 & i25) | (v3912 & ~i25),
  v4065 = (v27 & i30) | (v4066 & ~i30),
  v4066 = (v27 & i31) | (v4067 & ~i31),
  v4067 = (~v4068 & ~i32) | i32,
  v4068 = (v4075 & i35) | (v4069 & ~i35),
  v4069 = (v4074 & i36) | (v4070 & ~i36),
  v4070 = (v4073 & i37) | (v4071 & ~i37),
  v4071 = (v4072 & i38) | (v3916 & ~i38),
  v4072 = (v4045 & i40) | (v3918 & ~i40),
  v4073 = (v4072 & i38) | (v3917 & ~i38),
  v4074 = (v4073 & i37) | (v4072 & ~i37),
  v4075 = (v4074 & i36) | (v4076 & ~i36),
  v4076 = (v4073 & i37) | (v4077 & ~i37),
  v4077 = (v4072 & i38) | (v4078 & ~i38),
  v4078 = (v3916 & i39) | (v4072 & ~i39),
  v4079 = (v4080 & i21) | (v27 & ~i21),
  v4080 = (v4081 & i22) | (v3908 & ~i22),
  v4081 = (v4082 & i25) | (v3912 & ~i25),
  v4082 = (v27 & i30) | (v4083 & ~i30),
  v4083 = (v27 & i31) | (v4084 & ~i31),
  v4084 = (~v4085 & ~i32) | i32,
  v4085 = (v4092 & i35) | (v4086 & ~i35),
  v4086 = (v4091 & i36) | (v4087 & ~i36),
  v4087 = (v4090 & i37) | (v4088 & ~i37),
  v4088 = (v4089 & i38) | (v3916 & ~i38),
  v4089 = (v4058 & i40) | (v3918 & ~i40),
  v4090 = (v4089 & i38) | (v3917 & ~i38),
  v4091 = (v4090 & i37) | (v4089 & ~i37),
  v4092 = (v4091 & i36) | (v4093 & ~i36),
  v4093 = (v4090 & i37) | (v4094 & ~i37),
  v4094 = (v4089 & i38) | (v4095 & ~i38),
  v4095 = (v4089 & i39) | (v3916 & ~i39),
  v4096 = (v4132 & i19) | (v4097 & ~i19),
  v4097 = (v4115 & i20) | (v4098 & ~i20),
  v4098 = (v4099 & i21) | (v27 & ~i21),
  v4099 = (v4100 & i22) | (v3908 & ~i22),
  v4100 = (v4101 & i25) | (v3912 & ~i25),
  v4101 = (v27 & i30) | (v4102 & ~i30),
  v4102 = (v27 & i31) | (v4103 & ~i31),
  v4103 = (~v4104 & ~i32) | i32,
  v4104 = (v4112 & i35) | (v4105 & ~i35),
  v4105 = (v4111 & i36) | (v4106 & ~i36),
  v4106 = (v4110 & i37) | (v4107 & ~i37),
  v4107 = (v4109 & i38) | (v4108 & ~i38),
  v4108 = (v3916 & i39) | (v4109 & ~i39),
  v4109 = (v3918 & i40) | (v4045 & ~i40),
  v4110 = (v4109 & i38) | (v3917 & ~i38),
  v4111 = (v4110 & i37) | (v4109 & ~i37),
  v4112 = (v4111 & i36) | (v4113 & ~i36),
  v4113 = (v4110 & i37) | (v4114 & ~i37),
  v4114 = (v4109 & i38) | (v3916 & ~i38),
  v4115 = (v4116 & i21) | (v27 & ~i21),
  v4116 = (v4117 & i22) | (v3908 & ~i22),
  v4117 = (v4118 & i25) | (v3912 & ~i25),
  v4118 = (v27 & i30) | (v4119 & ~i30),
  v4119 = (v27 & i31) | (v4120 & ~i31),
  v4120 = (~v4121 & ~i32) | i32,
  v4121 = (v4129 & i35) | (v4122 & ~i35),
  v4122 = (v4128 & i36) | (v4123 & ~i36),
  v4123 = (v4127 & i37) | (v4124 & ~i37),
  v4124 = (v4126 & i38) | (v4125 & ~i38),
  v4125 = (v4126 & i39) | (v3916 & ~i39),
  v4126 = (v3918 & i40) | (v4058 & ~i40),
  v4127 = (v4126 & i38) | (v3917 & ~i38),
  v4128 = (v4127 & i37) | (v4126 & ~i37),
  v4129 = (v4128 & i36) | (v4130 & ~i36),
  v4130 = (v4127 & i37) | (v4131 & ~i37),
  v4131 = (v4126 & i38) | (v3916 & ~i38),
  v4132 = (v4133 & i21) | (v27 & ~i21),
  v4133 = (v4134 & i22) | (v3908 & ~i22),
  v4134 = (v4135 & i25) | (v3912 & ~i25),
  v4135 = (v27 & i30) | (v4136 & ~i30),
  v4136 = (v27 & i31) | (v4137 & ~i31),
  v4137 = (~v4138 & ~i32) | i32,
  v4138 = (v4142 & i36) | (v4139 & ~i36),
  v4139 = (v4141 & i37) | (v4140 & ~i37),
  v4140 = (v3918 & i38) | (v3916 & ~i38),
  v4141 = (v3918 & i38) | (v3917 & ~i38),
  v4142 = (v4141 & i37) | (v3918 & ~i37),
  v4143 = (v4206 & i16) | (v4144 & ~i16),
  v4144 = (v4182 & i17) | (v4145 & ~i17),
  v4145 = (v4165 & i19) | (v4146 & ~i19),
  v4146 = (v4156 & i20) | (v4147 & ~i20),
  v4147 = (v4148 & i21) | (v27 & ~i21),
  v4148 = (v4149 & i22) | (v3908 & ~i22),
  v4149 = (v4150 & i25) | (v3912 & ~i25),
  v4150 = (v27 & i30) | (v4151 & ~i30),
  v4151 = (v27 & i31) | (v4152 & ~i31),
  v4152 = (~v4153 & ~i32) | i32,
  v4153 = (v4154 & i36) | (v3924 & ~i36),
  v4154 = (v3931 & i37) | (v4155 & ~i37),
  v4155 = (v3927 & i38) | (v3916 & ~i38),
  v4156 = (v4157 & i21) | (v27 & ~i21),
  v4157 = (v4158 & i22) | (v3908 & ~i22),
  v4158 = (v4159 & i25) | (v3912 & ~i25),
  v4159 = (v27 & i30) | (v4160 & ~i30),
  v4160 = (v27 & i31) | (v4161 & ~i31),
  v4161 = (~v4162 & ~i32) | i32,
  v4162 = (v4163 & i36) | (v3940 & ~i36),
  v4163 = (v3947 & i37) | (v4164 & ~i37),
  v4164 = (v3943 & i38) | (v3916 & ~i38),
  v4165 = (v4174 & i20) | (v4166 & ~i20),
  v4166 = (v4167 & i21) | (v27 & ~i21),
  v4167 = (v4168 & i22) | (v3908 & ~i22),
  v4168 = (v4169 & i25) | (v3912 & ~i25),
  v4169 = (v27 & i30) | (v4170 & ~i30),
  v4170 = (v27 & i31) | (v4171 & ~i31),
  v4171 = (~v4172 & ~i32) | i32,
  v4172 = (v4173 & i35) | (v3958 & ~i35),
  v4173 = (v3958 & i36) | (v3965 & ~i36),
  v4174 = (v4175 & i21) | (v27 & ~i21),
  v4175 = (v4176 & i22) | (v3908 & ~i22),
  v4176 = (v4177 & i25) | (v3912 & ~i25),
  v4177 = (v27 & i30) | (v4178 & ~i30),
  v4178 = (v27 & i31) | (v4179 & ~i31),
  v4179 = (~v4180 & ~i32) | i32,
  v4180 = (v4181 & i35) | (v3976 & ~i35),
  v4181 = (v3976 & i36) | (v3982 & ~i36),
  v4182 = (v4200 & i19) | (v4183 & ~i19),
  v4183 = (v4192 & i20) | (v4184 & ~i20),
  v4184 = (v4185 & i21) | (v27 & ~i21),
  v4185 = (v4186 & i22) | (v3908 & ~i22),
  v4186 = (v4187 & i25) | (v3912 & ~i25),
  v4187 = (v27 & i30) | (v4188 & ~i30),
  v4188 = (v27 & i31) | (v4189 & ~i31),
  v4189 = (~v4190 & ~i32) | i32,
  v4190 = (v4002 & i35) | (v4191 & ~i35),
  v4191 = (v4002 & i36) | (v3995 & ~i36),
  v4192 = (v4193 & i21) | (v27 & ~i21),
  v4193 = (v4194 & i22) | (v3908 & ~i22),
  v4194 = (v4195 & i25) | (v3912 & ~i25),
  v4195 = (v27 & i30) | (v4196 & ~i30),
  v4196 = (v27 & i31) | (v4197 & ~i31),
  v4197 = (~v4198 & ~i32) | i32,
  v4198 = (v4019 & i35) | (v4199 & ~i35),
  v4199 = (v4019 & i36) | (v4012 & ~i36),
  v4200 = (v4201 & i21) | (v27 & ~i21),
  v4201 = (v4202 & i22) | (v3908 & ~i22),
  v4202 = (v4203 & i25) | (v3912 & ~i25),
  v4203 = (v27 & i30) | (v4204 & ~i30),
  v4204 = (v27 & i31) | (v4205 & ~i31),
  v4205 = (~v4028 & ~i32) | i32,
  v4206 = (v4244 & i17) | (v4207 & ~i17),
  v4207 = (v4227 & i19) | (v4208 & ~i19),
  v4208 = (v4218 & i20) | (v4209 & ~i20),
  v4209 = (v4210 & i21) | (v27 & ~i21),
  v4210 = (v4211 & i22) | (v3908 & ~i22),
  v4211 = (v4212 & i25) | (v3912 & ~i25),
  v4212 = (v27 & i30) | (v4213 & ~i30),
  v4213 = (v27 & i31) | (v4214 & ~i31),
  v4214 = (~v4215 & ~i32) | i32,
  v4215 = (v4216 & i36) | (v4042 & ~i36),
  v4216 = (v4046 & i37) | (v4217 & ~i37),
  v4217 = (v4045 & i38) | (v3916 & ~i38),
  v4218 = (v4219 & i21) | (v27 & ~i21),
  v4219 = (v4220 & i22) | (v3908 & ~i22),
  v4220 = (v4221 & i25) | (v3912 & ~i25),
  v4221 = (v27 & i30) | (v4222 & ~i30),
  v4222 = (v27 & i31) | (v4223 & ~i31),
  v4223 = (~v4224 & ~i32) | i32,
  v4224 = (v4225 & i36) | (v4055 & ~i36),
  v4225 = (v4059 & i37) | (v4226 & ~i37),
  v4226 = (v4058 & i38) | (v3916 & ~i38),
  v4227 = (v4236 & i20) | (v4228 & ~i20),
  v4228 = (v4229 & i21) | (v27 & ~i21),
  v4229 = (v4230 & i22) | (v3908 & ~i22),
  v4230 = (v4231 & i25) | (v3912 & ~i25),
  v4231 = (v27 & i30) | (v4232 & ~i30),
  v4232 = (v27 & i31) | (v4233 & ~i31),
  v4233 = (~v4234 & ~i32) | i32,
  v4234 = (v4235 & i35) | (v4070 & ~i35),
  v4235 = (v4070 & i36) | (v4076 & ~i36),
  v4236 = (v4237 & i21) | (v27 & ~i21),
  v4237 = (v4238 & i22) | (v3908 & ~i22),
  v4238 = (v4239 & i25) | (v3912 & ~i25),
  v4239 = (v27 & i30) | (v4240 & ~i30),
  v4240 = (v27 & i31) | (v4241 & ~i31),
  v4241 = (~v4242 & ~i32) | i32,
  v4242 = (v4243 & i35) | (v4087 & ~i35),
  v4243 = (v4087 & i36) | (v4093 & ~i36),
  v4244 = (v4262 & i19) | (v4245 & ~i19),
  v4245 = (v4254 & i20) | (v4246 & ~i20),
  v4246 = (v4247 & i21) | (v27 & ~i21),
  v4247 = (v4248 & i22) | (v3908 & ~i22),
  v4248 = (v4249 & i25) | (v3912 & ~i25),
  v4249 = (v27 & i30) | (v4250 & ~i30),
  v4250 = (v27 & i31) | (v4251 & ~i31),
  v4251 = (~v4252 & ~i32) | i32,
  v4252 = (v4113 & i35) | (v4253 & ~i35),
  v4253 = (v4113 & i36) | (v4106 & ~i36),
  v4254 = (v4255 & i21) | (v27 & ~i21),
  v4255 = (v4256 & i22) | (v3908 & ~i22),
  v4256 = (v4257 & i25) | (v3912 & ~i25),
  v4257 = (v27 & i30) | (v4258 & ~i30),
  v4258 = (v27 & i31) | (v4259 & ~i31),
  v4259 = (~v4260 & ~i32) | i32,
  v4260 = (v4130 & i35) | (v4261 & ~i35),
  v4261 = (v4130 & i36) | (v4123 & ~i36),
  v4262 = (v4263 & i21) | (v27 & ~i21),
  v4263 = (v4264 & i22) | (v3908 & ~i22),
  v4264 = (v4265 & i25) | (v3912 & ~i25),
  v4265 = (v27 & i30) | (v4266 & ~i30),
  v4266 = (v27 & i31) | (v4267 & ~i31),
  v4267 = (~v4139 & ~i32) | i32,
  v4268 = (v4394 & i15) | (v4269 & ~i15),
  v4269 = (v4332 & i16) | (v4270 & ~i16),
  v4270 = (v4306 & i17) | (v4271 & ~i17),
  v4271 = (v4289 & i19) | (v4272 & ~i19),
  v4272 = (v4281 & i20) | (v4273 & ~i20),
  v4273 = (v4274 & i21) | (v27 & ~i21),
  v4274 = (v4275 & i22) | (v3908 & ~i22),
  v4275 = (v3920 & i25) | (v4276 & ~i25),
  v4276 = (v4277 & i29) | (v3920 & ~i29),
  v4277 = (v27 & i30) | (v4278 & ~i30),
  v4278 = (v27 & i31) | (v4279 & ~i31),
  v4279 = (~v4280 & ~i32) | i32,
  v4280 = (v3915 & i33) | (v3923 & ~i33),
  v4281 = (v4282 & i21) | (v27 & ~i21),
  v4282 = (v4283 & i22) | (v3908 & ~i22),
  v4283 = (v3936 & i25) | (v4284 & ~i25),
  v4284 = (v4285 & i29) | (v3936 & ~i29),
  v4285 = (v27 & i30) | (v4286 & ~i30),
  v4286 = (v27 & i31) | (v4287 & ~i31),
  v4287 = (~v4288 & ~i32) | i32,
  v4288 = (v3915 & i33) | (v3939 & ~i33),
  v4289 = (v4298 & i20) | (v4290 & ~i20),
  v4290 = (v4291 & i21) | (v27 & ~i21),
  v4291 = (v4292 & i22) | (v3908 & ~i22),
  v4292 = (v3953 & i25) | (v4293 & ~i25),
  v4293 = (v4294 & i29) | (v3953 & ~i29),
  v4294 = (v27 & i30) | (v4295 & ~i30),
  v4295 = (v27 & i31) | (v4296 & ~i31),
  v4296 = (~v4297 & ~i32) | i32,
  v4297 = (v3915 & i33) | (v3956 & ~i33),
  v4298 = (v4299 & i21) | (v27 & ~i21),
  v4299 = (v4300 & i22) | (v3908 & ~i22),
  v4300 = (v3971 & i25) | (v4301 & ~i25),
  v4301 = (v4302 & i29) | (v3971 & ~i29),
  v4302 = (v27 & i30) | (v4303 & ~i30),
  v4303 = (v27 & i31) | (v4304 & ~i31),
  v4304 = (~v4305 & ~i32) | i32,
  v4305 = (v3915 & i33) | (v3974 & ~i33),
  v4306 = (v4324 & i19) | (v4307 & ~i19),
  v4307 = (v4316 & i20) | (v4308 & ~i20),
  v4308 = (v4309 & i21) | (v27 & ~i21),
  v4309 = (v4310 & i22) | (v3908 & ~i22),
  v4310 = (v3990 & i25) | (v4311 & ~i25),
  v4311 = (v4312 & i29) | (v3990 & ~i29),
  v4312 = (v27 & i30) | (v4313 & ~i30),
  v4313 = (v27 & i31) | (v4314 & ~i31),
  v4314 = (~v4315 & ~i32) | i32,
  v4315 = (v3915 & i33) | (v3993 & ~i33),
  v4316 = (v4317 & i21) | (v27 & ~i21),
  v4317 = (v4318 & i22) | (v3908 & ~i22),
  v4318 = (v4007 & i25) | (v4319 & ~i25),
  v4319 = (v4320 & i29) | (v4007 & ~i29),
  v4320 = (v27 & i30) | (v4321 & ~i30),
  v4321 = (v27 & i31) | (v4322 & ~i31),
  v4322 = (~v4323 & ~i32) | i32,
  v4323 = (v3915 & i33) | (v4010 & ~i33),
  v4324 = (v4325 & i21) | (v27 & ~i21),
  v4325 = (v4326 & i22) | (v3908 & ~i22),
  v4326 = (v4024 & i25) | (v4327 & ~i25),
  v4327 = (v4328 & i29) | (v4024 & ~i29),
  v4328 = (v27 & i30) | (v4329 & ~i30),
  v4329 = (v27 & i31) | (v4330 & ~i31),
  v4330 = (~v4331 & ~i32) | i32,
  v4331 = (v3915 & i33) | (v4027 & ~i33),
  v4332 = (v4368 & i17) | (v4333 & ~i17),
  v4333 = (v4351 & i19) | (v4334 & ~i19),
  v4334 = (v4343 & i20) | (v4335 & ~i20),
  v4335 = (v4336 & i21) | (v27 & ~i21),
  v4336 = (v4337 & i22) | (v3908 & ~i22),
  v4337 = (v4038 & i25) | (v4338 & ~i25),
  v4338 = (v4339 & i29) | (v4038 & ~i29),
  v4339 = (v27 & i30) | (v4340 & ~i30),
  v4340 = (v27 & i31) | (v4341 & ~i31),
  v4341 = (~v4342 & ~i32) | i32,
  v4342 = (v3915 & i33) | (v4041 & ~i33),
  v4343 = (v4344 & i21) | (v27 & ~i21),
  v4344 = (v4345 & i22) | (v3908 & ~i22),
  v4345 = (v4051 & i25) | (v4346 & ~i25),
  v4346 = (v4347 & i29) | (v4051 & ~i29),
  v4347 = (v27 & i30) | (v4348 & ~i30),
  v4348 = (v27 & i31) | (v4349 & ~i31),
  v4349 = (~v4350 & ~i32) | i32,
  v4350 = (v3915 & i33) | (v4054 & ~i33),
  v4351 = (v4360 & i20) | (v4352 & ~i20),
  v4352 = (v4353 & i21) | (v27 & ~i21),
  v4353 = (v4354 & i22) | (v3908 & ~i22),
  v4354 = (v4065 & i25) | (v4355 & ~i25),
  v4355 = (v4356 & i29) | (v4065 & ~i29),
  v4356 = (v27 & i30) | (v4357 & ~i30),
  v4357 = (v27 & i31) | (v4358 & ~i31),
  v4358 = (~v4359 & ~i32) | i32,
  v4359 = (v3915 & i33) | (v4068 & ~i33),
  v4360 = (v4361 & i21) | (v27 & ~i21),
  v4361 = (v4362 & i22) | (v3908 & ~i22),
  v4362 = (v4082 & i25) | (v4363 & ~i25),
  v4363 = (v4364 & i29) | (v4082 & ~i29),
  v4364 = (v27 & i30) | (v4365 & ~i30),
  v4365 = (v27 & i31) | (v4366 & ~i31),
  v4366 = (~v4367 & ~i32) | i32,
  v4367 = (v3915 & i33) | (v4085 & ~i33),
  v4368 = (v4386 & i19) | (v4369 & ~i19),
  v4369 = (v4378 & i20) | (v4370 & ~i20),
  v4370 = (v4371 & i21) | (v27 & ~i21),
  v4371 = (v4372 & i22) | (v3908 & ~i22),
  v4372 = (v4101 & i25) | (v4373 & ~i25),
  v4373 = (v4374 & i29) | (v4101 & ~i29),
  v4374 = (v27 & i30) | (v4375 & ~i30),
  v4375 = (v27 & i31) | (v4376 & ~i31),
  v4376 = (~v4377 & ~i32) | i32,
  v4377 = (v3915 & i33) | (v4104 & ~i33),
  v4378 = (v4379 & i21) | (v27 & ~i21),
  v4379 = (v4380 & i22) | (v3908 & ~i22),
  v4380 = (v4118 & i25) | (v4381 & ~i25),
  v4381 = (v4382 & i29) | (v4118 & ~i29),
  v4382 = (v27 & i30) | (v4383 & ~i30),
  v4383 = (v27 & i31) | (v4384 & ~i31),
  v4384 = (~v4385 & ~i32) | i32,
  v4385 = (v3915 & i33) | (v4121 & ~i33),
  v4386 = (v4387 & i21) | (v27 & ~i21),
  v4387 = (v4388 & i22) | (v3908 & ~i22),
  v4388 = (v4135 & i25) | (v4389 & ~i25),
  v4389 = (v4390 & i29) | (v4135 & ~i29),
  v4390 = (v27 & i30) | (v4391 & ~i30),
  v4391 = (v27 & i31) | (v4392 & ~i31),
  v4392 = (~v4393 & ~i32) | i32,
  v4393 = (v3915 & i33) | (v4138 & ~i33),
  v4394 = (v4457 & i16) | (v4395 & ~i16),
  v4395 = (v4431 & i17) | (v4396 & ~i17),
  v4396 = (v4414 & i19) | (v4397 & ~i19),
  v4397 = (v4406 & i20) | (v4398 & ~i20),
  v4398 = (v4399 & i21) | (v27 & ~i21),
  v4399 = (v4400 & i22) | (v3908 & ~i22),
  v4400 = (v4150 & i25) | (v4401 & ~i25),
  v4401 = (v4402 & i29) | (v4150 & ~i29),
  v4402 = (v27 & i30) | (v4403 & ~i30),
  v4403 = (v27 & i31) | (v4404 & ~i31),
  v4404 = (~v4405 & ~i32) | i32,
  v4405 = (v3915 & i33) | (v4153 & ~i33),
  v4406 = (v4407 & i21) | (v27 & ~i21),
  v4407 = (v4408 & i22) | (v3908 & ~i22),
  v4408 = (v4159 & i25) | (v4409 & ~i25),
  v4409 = (v4410 & i29) | (v4159 & ~i29),
  v4410 = (v27 & i30) | (v4411 & ~i30),
  v4411 = (v27 & i31) | (v4412 & ~i31),
  v4412 = (~v4413 & ~i32) | i32,
  v4413 = (v3915 & i33) | (v4162 & ~i33),
  v4414 = (v4423 & i20) | (v4415 & ~i20),
  v4415 = (v4416 & i21) | (v27 & ~i21),
  v4416 = (v4417 & i22) | (v3908 & ~i22),
  v4417 = (v4169 & i25) | (v4418 & ~i25),
  v4418 = (v4419 & i29) | (v4169 & ~i29),
  v4419 = (v27 & i30) | (v4420 & ~i30),
  v4420 = (v27 & i31) | (v4421 & ~i31),
  v4421 = (~v4422 & ~i32) | i32,
  v4422 = (v3915 & i33) | (v4172 & ~i33),
  v4423 = (v4424 & i21) | (v27 & ~i21),
  v4424 = (v4425 & i22) | (v3908 & ~i22),
  v4425 = (v4177 & i25) | (v4426 & ~i25),
  v4426 = (v4427 & i29) | (v4177 & ~i29),
  v4427 = (v27 & i30) | (v4428 & ~i30),
  v4428 = (v27 & i31) | (v4429 & ~i31),
  v4429 = (~v4430 & ~i32) | i32,
  v4430 = (v3915 & i33) | (v4180 & ~i33),
  v4431 = (v4449 & i19) | (v4432 & ~i19),
  v4432 = (v4441 & i20) | (v4433 & ~i20),
  v4433 = (v4434 & i21) | (v27 & ~i21),
  v4434 = (v4435 & i22) | (v3908 & ~i22),
  v4435 = (v4187 & i25) | (v4436 & ~i25),
  v4436 = (v4437 & i29) | (v4187 & ~i29),
  v4437 = (v27 & i30) | (v4438 & ~i30),
  v4438 = (v27 & i31) | (v4439 & ~i31),
  v4439 = (~v4440 & ~i32) | i32,
  v4440 = (v3915 & i33) | (v4190 & ~i33),
  v4441 = (v4442 & i21) | (v27 & ~i21),
  v4442 = (v4443 & i22) | (v3908 & ~i22),
  v4443 = (v4195 & i25) | (v4444 & ~i25),
  v4444 = (v4445 & i29) | (v4195 & ~i29),
  v4445 = (v27 & i30) | (v4446 & ~i30),
  v4446 = (v27 & i31) | (v4447 & ~i31),
  v4447 = (~v4448 & ~i32) | i32,
  v4448 = (v3915 & i33) | (v4198 & ~i33),
  v4449 = (v4450 & i21) | (v27 & ~i21),
  v4450 = (v4451 & i22) | (v3908 & ~i22),
  v4451 = (v4203 & i25) | (v4452 & ~i25),
  v4452 = (v4453 & i29) | (v4203 & ~i29),
  v4453 = (v27 & i30) | (v4454 & ~i30),
  v4454 = (v27 & i31) | (v4455 & ~i31),
  v4455 = (~v4456 & ~i32) | i32,
  v4456 = (v3915 & i33) | (v4028 & ~i33),
  v4457 = (v4493 & i17) | (v4458 & ~i17),
  v4458 = (v4476 & i19) | (v4459 & ~i19),
  v4459 = (v4468 & i20) | (v4460 & ~i20),
  v4460 = (v4461 & i21) | (v27 & ~i21),
  v4461 = (v4462 & i22) | (v3908 & ~i22),
  v4462 = (v4212 & i25) | (v4463 & ~i25),
  v4463 = (v4464 & i29) | (v4212 & ~i29),
  v4464 = (v27 & i30) | (v4465 & ~i30),
  v4465 = (v27 & i31) | (v4466 & ~i31),
  v4466 = (~v4467 & ~i32) | i32,
  v4467 = (v3915 & i33) | (v4215 & ~i33),
  v4468 = (v4469 & i21) | (v27 & ~i21),
  v4469 = (v4470 & i22) | (v3908 & ~i22),
  v4470 = (v4221 & i25) | (v4471 & ~i25),
  v4471 = (v4472 & i29) | (v4221 & ~i29),
  v4472 = (v27 & i30) | (v4473 & ~i30),
  v4473 = (v27 & i31) | (v4474 & ~i31),
  v4474 = (~v4475 & ~i32) | i32,
  v4475 = (v3915 & i33) | (v4224 & ~i33),
  v4476 = (v4485 & i20) | (v4477 & ~i20),
  v4477 = (v4478 & i21) | (v27 & ~i21),
  v4478 = (v4479 & i22) | (v3908 & ~i22),
  v4479 = (v4231 & i25) | (v4480 & ~i25),
  v4480 = (v4481 & i29) | (v4231 & ~i29),
  v4481 = (v27 & i30) | (v4482 & ~i30),
  v4482 = (v27 & i31) | (v4483 & ~i31),
  v4483 = (~v4484 & ~i32) | i32,
  v4484 = (v3915 & i33) | (v4234 & ~i33),
  v4485 = (v4486 & i21) | (v27 & ~i21),
  v4486 = (v4487 & i22) | (v3908 & ~i22),
  v4487 = (v4239 & i25) | (v4488 & ~i25),
  v4488 = (v4489 & i29) | (v4239 & ~i29),
  v4489 = (v27 & i30) | (v4490 & ~i30),
  v4490 = (v27 & i31) | (v4491 & ~i31),
  v4491 = (~v4492 & ~i32) | i32,
  v4492 = (v3915 & i33) | (v4242 & ~i33),
  v4493 = (v4511 & i19) | (v4494 & ~i19),
  v4494 = (v4503 & i20) | (v4495 & ~i20),
  v4495 = (v4496 & i21) | (v27 & ~i21),
  v4496 = (v4497 & i22) | (v3908 & ~i22),
  v4497 = (v4249 & i25) | (v4498 & ~i25),
  v4498 = (v4499 & i29) | (v4249 & ~i29),
  v4499 = (v27 & i30) | (v4500 & ~i30),
  v4500 = (v27 & i31) | (v4501 & ~i31),
  v4501 = (~v4502 & ~i32) | i32,
  v4502 = (v3915 & i33) | (v4252 & ~i33),
  v4503 = (v4504 & i21) | (v27 & ~i21),
  v4504 = (v4505 & i22) | (v3908 & ~i22),
  v4505 = (v4257 & i25) | (v4506 & ~i25),
  v4506 = (v4507 & i29) | (v4257 & ~i29),
  v4507 = (v27 & i30) | (v4508 & ~i30),
  v4508 = (v27 & i31) | (v4509 & ~i31),
  v4509 = (~v4510 & ~i32) | i32,
  v4510 = (v3915 & i33) | (v4260 & ~i33),
  v4511 = (v4512 & i21) | (v27 & ~i21),
  v4512 = (v4513 & i22) | (v3908 & ~i22),
  v4513 = (v4265 & i25) | (v4514 & ~i25),
  v4514 = (v4515 & i29) | (v4265 & ~i29),
  v4515 = (v27 & i30) | (v4516 & ~i30),
  v4516 = (v27 & i31) | (v4517 & ~i31),
  v4517 = (~v4518 & ~i32) | i32,
  v4518 = (v3915 & i33) | (v4139 & ~i33),
  v4519 = (v4523 & i11) | (v4520 & ~i11),
  v4520 = (v4523 & i12) | (v4521 & ~i12),
  v4521 = (v4523 & i13) | (v4522 & ~i13),
  v4522 = (v4746 & i14) | (v4523 & ~i14),
  v4523 = (v4635 & i15) | (v4524 & ~i15),
  v4524 = (v4580 & i16) | (v4525 & ~i16),
  v4525 = (v4557 & i17) | (v4526 & ~i17),
  v4526 = (v4542 & i19) | (v4527 & ~i19),
  v4527 = (v4535 & i20) | (v4528 & ~i20),
  v4528 = (v4529 & i21) | (v27 & ~i21),
  v4529 = (v4530 & i22) | (v3908 & ~i22),
  v4530 = (v4531 & i29) | (v3920 & ~i29),
  v4531 = (v27 & i30) | (v4532 & ~i30),
  v4532 = (v27 & i31) | (v4533 & ~i31),
  v4533 = (~v4534 & ~i32) | i32,
  v4534 = (v3923 & i33) | (v3915 & ~i33),
  v4535 = (v4536 & i21) | (v27 & ~i21),
  v4536 = (v4537 & i22) | (v3908 & ~i22),
  v4537 = (v4538 & i29) | (v3936 & ~i29),
  v4538 = (v27 & i30) | (v4539 & ~i30),
  v4539 = (v27 & i31) | (v4540 & ~i31),
  v4540 = (~v4541 & ~i32) | i32,
  v4541 = (v3939 & i33) | (v3915 & ~i33),
  v4542 = (v4550 & i20) | (v4543 & ~i20),
  v4543 = (v4544 & i21) | (v27 & ~i21),
  v4544 = (v4545 & i22) | (v3908 & ~i22),
  v4545 = (v4546 & i29) | (v3953 & ~i29),
  v4546 = (v27 & i30) | (v4547 & ~i30),
  v4547 = (v27 & i31) | (v4548 & ~i31),
  v4548 = (~v4549 & ~i32) | i32,
  v4549 = (v3956 & i33) | (v3915 & ~i33),
  v4550 = (v4551 & i21) | (v27 & ~i21),
  v4551 = (v4552 & i22) | (v3908 & ~i22),
  v4552 = (v4553 & i29) | (v3971 & ~i29),
  v4553 = (v27 & i30) | (v4554 & ~i30),
  v4554 = (v27 & i31) | (v4555 & ~i31),
  v4555 = (~v4556 & ~i32) | i32,
  v4556 = (v3974 & i33) | (v3915 & ~i33),
  v4557 = (v4573 & i19) | (v4558 & ~i19),
  v4558 = (v4566 & i20) | (v4559 & ~i20),
  v4559 = (v4560 & i21) | (v27 & ~i21),
  v4560 = (v4561 & i22) | (v3908 & ~i22),
  v4561 = (v4562 & i29) | (v3990 & ~i29),
  v4562 = (v27 & i30) | (v4563 & ~i30),
  v4563 = (v27 & i31) | (v4564 & ~i31),
  v4564 = (~v4565 & ~i32) | i32,
  v4565 = (v3993 & i33) | (v3915 & ~i33),
  v4566 = (v4567 & i21) | (v27 & ~i21),
  v4567 = (v4568 & i22) | (v3908 & ~i22),
  v4568 = (v4569 & i29) | (v4007 & ~i29),
  v4569 = (v27 & i30) | (v4570 & ~i30),
  v4570 = (v27 & i31) | (v4571 & ~i31),
  v4571 = (~v4572 & ~i32) | i32,
  v4572 = (v4010 & i33) | (v3915 & ~i33),
  v4573 = (v4574 & i21) | (v27 & ~i21),
  v4574 = (v4575 & i22) | (v3908 & ~i22),
  v4575 = (v4576 & i29) | (v4024 & ~i29),
  v4576 = (v27 & i30) | (v4577 & ~i30),
  v4577 = (v27 & i31) | (v4578 & ~i31),
  v4578 = (~v4579 & ~i32) | i32,
  v4579 = (v4027 & i33) | (v3915 & ~i33),
  v4580 = (v4612 & i17) | (v4581 & ~i17),
  v4581 = (v4597 & i19) | (v4582 & ~i19),
  v4582 = (v4590 & i20) | (v4583 & ~i20),
  v4583 = (v4584 & i21) | (v27 & ~i21),
  v4584 = (v4585 & i22) | (v3908 & ~i22),
  v4585 = (v4586 & i29) | (v4038 & ~i29),
  v4586 = (v27 & i30) | (v4587 & ~i30),
  v4587 = (v27 & i31) | (v4588 & ~i31),
  v4588 = (~v4589 & ~i32) | i32,
  v4589 = (v4041 & i33) | (v3915 & ~i33),
  v4590 = (v4591 & i21) | (v27 & ~i21),
  v4591 = (v4592 & i22) | (v3908 & ~i22),
  v4592 = (v4593 & i29) | (v4051 & ~i29),
  v4593 = (v27 & i30) | (v4594 & ~i30),
  v4594 = (v27 & i31) | (v4595 & ~i31),
  v4595 = (~v4596 & ~i32) | i32,
  v4596 = (v4054 & i33) | (v3915 & ~i33),
  v4597 = (v4605 & i20) | (v4598 & ~i20),
  v4598 = (v4599 & i21) | (v27 & ~i21),
  v4599 = (v4600 & i22) | (v3908 & ~i22),
  v4600 = (v4601 & i29) | (v4065 & ~i29),
  v4601 = (v27 & i30) | (v4602 & ~i30),
  v4602 = (v27 & i31) | (v4603 & ~i31),
  v4603 = (~v4604 & ~i32) | i32,
  v4604 = (v4068 & i33) | (v3915 & ~i33),
  v4605 = (v4606 & i21) | (v27 & ~i21),
  v4606 = (v4607 & i22) | (v3908 & ~i22),
  v4607 = (v4608 & i29) | (v4082 & ~i29),
  v4608 = (v27 & i30) | (v4609 & ~i30),
  v4609 = (v27 & i31) | (v4610 & ~i31),
  v4610 = (~v4611 & ~i32) | i32,
  v4611 = (v4085 & i33) | (v3915 & ~i33),
  v4612 = (v4628 & i19) | (v4613 & ~i19),
  v4613 = (v4621 & i20) | (v4614 & ~i20),
  v4614 = (v4615 & i21) | (v27 & ~i21),
  v4615 = (v4616 & i22) | (v3908 & ~i22),
  v4616 = (v4617 & i29) | (v4101 & ~i29),
  v4617 = (v27 & i30) | (v4618 & ~i30),
  v4618 = (v27 & i31) | (v4619 & ~i31),
  v4619 = (~v4620 & ~i32) | i32,
  v4620 = (v4104 & i33) | (v3915 & ~i33),
  v4621 = (v4622 & i21) | (v27 & ~i21),
  v4622 = (v4623 & i22) | (v3908 & ~i22),
  v4623 = (v4624 & i29) | (v4118 & ~i29),
  v4624 = (v27 & i30) | (v4625 & ~i30),
  v4625 = (v27 & i31) | (v4626 & ~i31),
  v4626 = (~v4627 & ~i32) | i32,
  v4627 = (v4121 & i33) | (v3915 & ~i33),
  v4628 = (v4629 & i21) | (v27 & ~i21),
  v4629 = (v4630 & i22) | (v3908 & ~i22),
  v4630 = (v4631 & i29) | (v4135 & ~i29),
  v4631 = (v27 & i30) | (v4632 & ~i30),
  v4632 = (v27 & i31) | (v4633 & ~i31),
  v4633 = (~v4634 & ~i32) | i32,
  v4634 = (v4138 & i33) | (v3915 & ~i33),
  v4635 = (v4691 & i16) | (v4636 & ~i16),
  v4636 = (v4668 & i17) | (v4637 & ~i17),
  v4637 = (v4653 & i19) | (v4638 & ~i19),
  v4638 = (v4646 & i20) | (v4639 & ~i20),
  v4639 = (v4640 & i21) | (v27 & ~i21),
  v4640 = (v4641 & i22) | (v3908 & ~i22),
  v4641 = (v4642 & i29) | (v4150 & ~i29),
  v4642 = (v27 & i30) | (v4643 & ~i30),
  v4643 = (v27 & i31) | (v4644 & ~i31),
  v4644 = (~v4645 & ~i32) | i32,
  v4645 = (v4153 & i33) | (v3915 & ~i33),
  v4646 = (v4647 & i21) | (v27 & ~i21),
  v4647 = (v4648 & i22) | (v3908 & ~i22),
  v4648 = (v4649 & i29) | (v4159 & ~i29),
  v4649 = (v27 & i30) | (v4650 & ~i30),
  v4650 = (v27 & i31) | (v4651 & ~i31),
  v4651 = (~v4652 & ~i32) | i32,
  v4652 = (v4162 & i33) | (v3915 & ~i33),
  v4653 = (v4661 & i20) | (v4654 & ~i20),
  v4654 = (v4655 & i21) | (v27 & ~i21),
  v4655 = (v4656 & i22) | (v3908 & ~i22),
  v4656 = (v4657 & i29) | (v4169 & ~i29),
  v4657 = (v27 & i30) | (v4658 & ~i30),
  v4658 = (v27 & i31) | (v4659 & ~i31),
  v4659 = (~v4660 & ~i32) | i32,
  v4660 = (v4172 & i33) | (v3915 & ~i33),
  v4661 = (v4662 & i21) | (v27 & ~i21),
  v4662 = (v4663 & i22) | (v3908 & ~i22),
  v4663 = (v4664 & i29) | (v4177 & ~i29),
  v4664 = (v27 & i30) | (v4665 & ~i30),
  v4665 = (v27 & i31) | (v4666 & ~i31),
  v4666 = (~v4667 & ~i32) | i32,
  v4667 = (v4180 & i33) | (v3915 & ~i33),
  v4668 = (v4684 & i19) | (v4669 & ~i19),
  v4669 = (v4677 & i20) | (v4670 & ~i20),
  v4670 = (v4671 & i21) | (v27 & ~i21),
  v4671 = (v4672 & i22) | (v3908 & ~i22),
  v4672 = (v4673 & i29) | (v4187 & ~i29),
  v4673 = (v27 & i30) | (v4674 & ~i30),
  v4674 = (v27 & i31) | (v4675 & ~i31),
  v4675 = (~v4676 & ~i32) | i32,
  v4676 = (v4190 & i33) | (v3915 & ~i33),
  v4677 = (v4678 & i21) | (v27 & ~i21),
  v4678 = (v4679 & i22) | (v3908 & ~i22),
  v4679 = (v4680 & i29) | (v4195 & ~i29),
  v4680 = (v27 & i30) | (v4681 & ~i30),
  v4681 = (v27 & i31) | (v4682 & ~i31),
  v4682 = (~v4683 & ~i32) | i32,
  v4683 = (v4198 & i33) | (v3915 & ~i33),
  v4684 = (v4685 & i21) | (v27 & ~i21),
  v4685 = (v4686 & i22) | (v3908 & ~i22),
  v4686 = (v4687 & i29) | (v4203 & ~i29),
  v4687 = (v27 & i30) | (v4688 & ~i30),
  v4688 = (v27 & i31) | (v4689 & ~i31),
  v4689 = (~v4690 & ~i32) | i32,
  v4690 = (v4028 & i33) | (v3915 & ~i33),
  v4691 = (v4723 & i17) | (v4692 & ~i17),
  v4692 = (v4708 & i19) | (v4693 & ~i19),
  v4693 = (v4701 & i20) | (v4694 & ~i20),
  v4694 = (v4695 & i21) | (v27 & ~i21),
  v4695 = (v4696 & i22) | (v3908 & ~i22),
  v4696 = (v4697 & i29) | (v4212 & ~i29),
  v4697 = (v27 & i30) | (v4698 & ~i30),
  v4698 = (v27 & i31) | (v4699 & ~i31),
  v4699 = (~v4700 & ~i32) | i32,
  v4700 = (v4215 & i33) | (v3915 & ~i33),
  v4701 = (v4702 & i21) | (v27 & ~i21),
  v4702 = (v4703 & i22) | (v3908 & ~i22),
  v4703 = (v4704 & i29) | (v4221 & ~i29),
  v4704 = (v27 & i30) | (v4705 & ~i30),
  v4705 = (v27 & i31) | (v4706 & ~i31),
  v4706 = (~v4707 & ~i32) | i32,
  v4707 = (v4224 & i33) | (v3915 & ~i33),
  v4708 = (v4716 & i20) | (v4709 & ~i20),
  v4709 = (v4710 & i21) | (v27 & ~i21),
  v4710 = (v4711 & i22) | (v3908 & ~i22),
  v4711 = (v4712 & i29) | (v4231 & ~i29),
  v4712 = (v27 & i30) | (v4713 & ~i30),
  v4713 = (v27 & i31) | (v4714 & ~i31),
  v4714 = (~v4715 & ~i32) | i32,
  v4715 = (v4234 & i33) | (v3915 & ~i33),
  v4716 = (v4717 & i21) | (v27 & ~i21),
  v4717 = (v4718 & i22) | (v3908 & ~i22),
  v4718 = (v4719 & i29) | (v4239 & ~i29),
  v4719 = (v27 & i30) | (v4720 & ~i30),
  v4720 = (v27 & i31) | (v4721 & ~i31),
  v4721 = (~v4722 & ~i32) | i32,
  v4722 = (v4242 & i33) | (v3915 & ~i33),
  v4723 = (v4739 & i19) | (v4724 & ~i19),
  v4724 = (v4732 & i20) | (v4725 & ~i20),
  v4725 = (v4726 & i21) | (v27 & ~i21),
  v4726 = (v4727 & i22) | (v3908 & ~i22),
  v4727 = (v4728 & i29) | (v4249 & ~i29),
  v4728 = (v27 & i30) | (v4729 & ~i30),
  v4729 = (v27 & i31) | (v4730 & ~i31),
  v4730 = (~v4731 & ~i32) | i32,
  v4731 = (v4252 & i33) | (v3915 & ~i33),
  v4732 = (v4733 & i21) | (v27 & ~i21),
  v4733 = (v4734 & i22) | (v3908 & ~i22),
  v4734 = (v4735 & i29) | (v4257 & ~i29),
  v4735 = (v27 & i30) | (v4736 & ~i30),
  v4736 = (v27 & i31) | (v4737 & ~i31),
  v4737 = (~v4738 & ~i32) | i32,
  v4738 = (v4260 & i33) | (v3915 & ~i33),
  v4739 = (v4740 & i21) | (v27 & ~i21),
  v4740 = (v4741 & i22) | (v3908 & ~i22),
  v4741 = (v4742 & i29) | (v4265 & ~i29),
  v4742 = (v27 & i30) | (v4743 & ~i30),
  v4743 = (v27 & i31) | (v4744 & ~i31),
  v4744 = (~v4745 & ~i32) | i32,
  v4745 = (v4139 & i33) | (v3915 & ~i33),
  v4746 = (v4788 & i15) | (v4747 & ~i15),
  v4747 = (v4768 & i16) | (v4748 & ~i16),
  v4748 = (v4760 & i17) | (v4749 & ~i17),
  v4749 = (v4755 & i19) | (v4750 & ~i19),
  v4750 = (v4753 & i20) | (v4751 & ~i20),
  v4751 = (v4752 & i21) | (v27 & ~i21),
  v4752 = (v3920 & i22) | (v3908 & ~i22),
  v4753 = (v4754 & i21) | (v27 & ~i21),
  v4754 = (v3936 & i22) | (v3908 & ~i22),
  v4755 = (v4758 & i20) | (v4756 & ~i20),
  v4756 = (v4757 & i21) | (v27 & ~i21),
  v4757 = (v3953 & i22) | (v3908 & ~i22),
  v4758 = (v4759 & i21) | (v27 & ~i21),
  v4759 = (v3971 & i22) | (v3908 & ~i22),
  v4760 = (v4766 & i19) | (v4761 & ~i19),
  v4761 = (v4764 & i20) | (v4762 & ~i20),
  v4762 = (v4763 & i21) | (v27 & ~i21),
  v4763 = (v3990 & i22) | (v3908 & ~i22),
  v4764 = (v4765 & i21) | (v27 & ~i21),
  v4765 = (v4007 & i22) | (v3908 & ~i22),
  v4766 = (v4767 & i21) | (v27 & ~i21),
  v4767 = (v4024 & i22) | (v3908 & ~i22),
  v4768 = (v4780 & i17) | (v4769 & ~i17),
  v4769 = (v4775 & i19) | (v4770 & ~i19),
  v4770 = (v4773 & i20) | (v4771 & ~i20),
  v4771 = (v4772 & i21) | (v27 & ~i21),
  v4772 = (v4038 & i22) | (v3908 & ~i22),
  v4773 = (v4774 & i21) | (v27 & ~i21),
  v4774 = (v4051 & i22) | (v3908 & ~i22),
  v4775 = (v4778 & i20) | (v4776 & ~i20),
  v4776 = (v4777 & i21) | (v27 & ~i21),
  v4777 = (v4065 & i22) | (v3908 & ~i22),
  v4778 = (v4779 & i21) | (v27 & ~i21),
  v4779 = (v4082 & i22) | (v3908 & ~i22),
  v4780 = (v4786 & i19) | (v4781 & ~i19),
  v4781 = (v4784 & i20) | (v4782 & ~i20),
  v4782 = (v4783 & i21) | (v27 & ~i21),
  v4783 = (v4101 & i22) | (v3908 & ~i22),
  v4784 = (v4785 & i21) | (v27 & ~i21),
  v4785 = (v4118 & i22) | (v3908 & ~i22),
  v4786 = (v4787 & i21) | (v27 & ~i21),
  v4787 = (v4135 & i22) | (v3908 & ~i22),
  v4788 = (v4809 & i16) | (v4789 & ~i16),
  v4789 = (v4801 & i17) | (v4790 & ~i17),
  v4790 = (v4796 & i19) | (v4791 & ~i19),
  v4791 = (v4794 & i20) | (v4792 & ~i20),
  v4792 = (v4793 & i21) | (v27 & ~i21),
  v4793 = (v4150 & i22) | (v3908 & ~i22),
  v4794 = (v4795 & i21) | (v27 & ~i21),
  v4795 = (v4159 & i22) | (v3908 & ~i22),
  v4796 = (v4799 & i20) | (v4797 & ~i20),
  v4797 = (v4798 & i21) | (v27 & ~i21),
  v4798 = (v4169 & i22) | (v3908 & ~i22),
  v4799 = (v4800 & i21) | (v27 & ~i21),
  v4800 = (v4177 & i22) | (v3908 & ~i22),
  v4801 = (v4807 & i19) | (v4802 & ~i19),
  v4802 = (v4805 & i20) | (v4803 & ~i20),
  v4803 = (v4804 & i21) | (v27 & ~i21),
  v4804 = (v4187 & i22) | (v3908 & ~i22),
  v4805 = (v4806 & i21) | (v27 & ~i21),
  v4806 = (v4195 & i22) | (v3908 & ~i22),
  v4807 = (v4808 & i21) | (v27 & ~i21),
  v4808 = (v4203 & i22) | (v3908 & ~i22),
  v4809 = (v4821 & i17) | (v4810 & ~i17),
  v4810 = (v4816 & i19) | (v4811 & ~i19),
  v4811 = (v4814 & i20) | (v4812 & ~i20),
  v4812 = (v4813 & i21) | (v27 & ~i21),
  v4813 = (v4212 & i22) | (v3908 & ~i22),
  v4814 = (v4815 & i21) | (v27 & ~i21),
  v4815 = (v4221 & i22) | (v3908 & ~i22),
  v4816 = (v4819 & i20) | (v4817 & ~i20),
  v4817 = (v4818 & i21) | (v27 & ~i21),
  v4818 = (v4231 & i22) | (v3908 & ~i22),
  v4819 = (v4820 & i21) | (v27 & ~i21),
  v4820 = (v4239 & i22) | (v3908 & ~i22),
  v4821 = (v4827 & i19) | (v4822 & ~i19),
  v4822 = (v4825 & i20) | (v4823 & ~i20),
  v4823 = (v4824 & i21) | (v27 & ~i21),
  v4824 = (v4249 & i22) | (v3908 & ~i22),
  v4825 = (v4826 & i21) | (v27 & ~i21),
  v4826 = (v4257 & i22) | (v3908 & ~i22),
  v4827 = (v4828 & i21) | (v27 & ~i21),
  v4828 = (v4265 & i22) | (v3908 & ~i22),
  v4829 = (v4833 & i11) | (v4830 & ~i11),
  v4830 = (v4833 & i12) | (v4831 & ~i12),
  v4831 = (v4833 & i13) | (v4832 & ~i13),
  v4832 = (v4835 & i14) | (v4833 & ~i14),
  v4833 = (v4834 & i21) | (v27 & ~i21),
  v4834 = (v3912 & i22) | (v3908 & ~i22),
  v4835 = (v4877 & i15) | (v4836 & ~i15),
  v4836 = (v4857 & i16) | (v4837 & ~i16),
  v4837 = (v4849 & i17) | (v4838 & ~i17),
  v4838 = (v4844 & i19) | (v4839 & ~i19),
  v4839 = (v4842 & i20) | (v4840 & ~i20),
  v4840 = (v4841 & i21) | (v27 & ~i21),
  v4841 = (v4276 & i22) | (v3908 & ~i22),
  v4842 = (v4843 & i21) | (v27 & ~i21),
  v4843 = (v4284 & i22) | (v3908 & ~i22),
  v4844 = (v4847 & i20) | (v4845 & ~i20),
  v4845 = (v4846 & i21) | (v27 & ~i21),
  v4846 = (v4293 & i22) | (v3908 & ~i22),
  v4847 = (v4848 & i21) | (v27 & ~i21),
  v4848 = (v4301 & i22) | (v3908 & ~i22),
  v4849 = (v4855 & i19) | (v4850 & ~i19),
  v4850 = (v4853 & i20) | (v4851 & ~i20),
  v4851 = (v4852 & i21) | (v27 & ~i21),
  v4852 = (v4311 & i22) | (v3908 & ~i22),
  v4853 = (v4854 & i21) | (v27 & ~i21),
  v4854 = (v4319 & i22) | (v3908 & ~i22),
  v4855 = (v4856 & i21) | (v27 & ~i21),
  v4856 = (v4327 & i22) | (v3908 & ~i22),
  v4857 = (v4869 & i17) | (v4858 & ~i17),
  v4858 = (v4864 & i19) | (v4859 & ~i19),
  v4859 = (v4862 & i20) | (v4860 & ~i20),
  v4860 = (v4861 & i21) | (v27 & ~i21),
  v4861 = (v4338 & i22) | (v3908 & ~i22),
  v4862 = (v4863 & i21) | (v27 & ~i21),
  v4863 = (v4346 & i22) | (v3908 & ~i22),
  v4864 = (v4867 & i20) | (v4865 & ~i20),
  v4865 = (v4866 & i21) | (v27 & ~i21),
  v4866 = (v4355 & i22) | (v3908 & ~i22),
  v4867 = (v4868 & i21) | (v27 & ~i21),
  v4868 = (v4363 & i22) | (v3908 & ~i22),
  v4869 = (v4875 & i19) | (v4870 & ~i19),
  v4870 = (v4873 & i20) | (v4871 & ~i20),
  v4871 = (v4872 & i21) | (v27 & ~i21),
  v4872 = (v4373 & i22) | (v3908 & ~i22),
  v4873 = (v4874 & i21) | (v27 & ~i21),
  v4874 = (v4381 & i22) | (v3908 & ~i22),
  v4875 = (v4876 & i21) | (v27 & ~i21),
  v4876 = (v4389 & i22) | (v3908 & ~i22),
  v4877 = (v4898 & i16) | (v4878 & ~i16),
  v4878 = (v4890 & i17) | (v4879 & ~i17),
  v4879 = (v4885 & i19) | (v4880 & ~i19),
  v4880 = (v4883 & i20) | (v4881 & ~i20),
  v4881 = (v4882 & i21) | (v27 & ~i21),
  v4882 = (v4401 & i22) | (v3908 & ~i22),
  v4883 = (v4884 & i21) | (v27 & ~i21),
  v4884 = (v4409 & i22) | (v3908 & ~i22),
  v4885 = (v4888 & i20) | (v4886 & ~i20),
  v4886 = (v4887 & i21) | (v27 & ~i21),
  v4887 = (v4418 & i22) | (v3908 & ~i22),
  v4888 = (v4889 & i21) | (v27 & ~i21),
  v4889 = (v4426 & i22) | (v3908 & ~i22),
  v4890 = (v4896 & i19) | (v4891 & ~i19),
  v4891 = (v4894 & i20) | (v4892 & ~i20),
  v4892 = (v4893 & i21) | (v27 & ~i21),
  v4893 = (v4436 & i22) | (v3908 & ~i22),
  v4894 = (v4895 & i21) | (v27 & ~i21),
  v4895 = (v4444 & i22) | (v3908 & ~i22),
  v4896 = (v4897 & i21) | (v27 & ~i21),
  v4897 = (v4452 & i22) | (v3908 & ~i22),
  v4898 = (v4910 & i17) | (v4899 & ~i17),
  v4899 = (v4905 & i19) | (v4900 & ~i19),
  v4900 = (v4903 & i20) | (v4901 & ~i20),
  v4901 = (v4902 & i21) | (v27 & ~i21),
  v4902 = (v4463 & i22) | (v3908 & ~i22),
  v4903 = (v4904 & i21) | (v27 & ~i21),
  v4904 = (v4471 & i22) | (v3908 & ~i22),
  v4905 = (v4908 & i20) | (v4906 & ~i20),
  v4906 = (v4907 & i21) | (v27 & ~i21),
  v4907 = (v4480 & i22) | (v3908 & ~i22),
  v4908 = (v4909 & i21) | (v27 & ~i21),
  v4909 = (v4488 & i22) | (v3908 & ~i22),
  v4910 = (v4916 & i19) | (v4911 & ~i19),
  v4911 = (v4914 & i20) | (v4912 & ~i20),
  v4912 = (v4913 & i21) | (v27 & ~i21),
  v4913 = (v4498 & i22) | (v3908 & ~i22),
  v4914 = (v4915 & i21) | (v27 & ~i21),
  v4915 = (v4506 & i22) | (v3908 & ~i22),
  v4916 = (v4917 & i21) | (v27 & ~i21),
  v4917 = (v4514 & i22) | (v3908 & ~i22),
  v4918 = (v6282 & i7) | (v4919 & ~i7),
  v4919 = (v5856 & i8) | (v4920 & ~i8),
  v4920 = (v5843 & i9) | (v4921 & ~i9),
  v4921 = (v5419 & i10) | (v4922 & ~i10),
  v4922 = (v5274 & i11) | (v4923 & ~i11),
  v4923 = (v4924 & i12) | (v3899 & ~i12),
  v4924 = (v3901 & i13) | (v4925 & ~i13),
  v4925 = (v5132 & i14) | (v4926 & ~i14),
  v4926 = (v5035 & i15) | (v4927 & ~i15),
  v4927 = (v4987 & i16) | (v4928 & ~i16),
  v4928 = (v4967 & i17) | (v4929 & ~i17),
  v4929 = (v4954 & i19) | (v4930 & ~i19),
  v4930 = (v4948 & i20) | (v4931 & ~i20),
  v4931 = (v4937 & i21) | (v4932 & ~i21),
  v4932 = (v27 & i26) | (v4933 & ~i26),
  v4933 = (v27 & i27) | (v4934 & ~i27),
  v4934 = (v4935 & i30) | (v27 & ~i30),
  v4935 = (v27 & i31) | (~v4936 & ~i31),
  v4936 = (v63 & i32) | ~i32,
  v4937 = (v4941 & i22) | (v4938 & ~i22),
  v4938 = (v3908 & i26) | (v4939 & ~i26),
  v4939 = (v3908 & i27) | (v4940 & ~i27),
  v4940 = (v4935 & i30) | (v3909 & ~i30),
  v4941 = (v4945 & i25) | (v4942 & ~i25),
  v4942 = (v3912 & i26) | (v4943 & ~i26),
  v4943 = (v3912 & i27) | (v4944 & ~i27),
  v4944 = (v4935 & i30) | (v3913 & ~i30),
  v4945 = (v3920 & i26) | (v4946 & ~i26),
  v4946 = (v3920 & i27) | (v4947 & ~i27),
  v4947 = (v4935 & i30) | (v3921 & ~i30),
  v4948 = (v4949 & i21) | (v4932 & ~i21),
  v4949 = (v4950 & i22) | (v4938 & ~i22),
  v4950 = (v4951 & i25) | (v4942 & ~i25),
  v4951 = (v3936 & i26) | (v4952 & ~i26),
  v4952 = (v3936 & i27) | (v4953 & ~i27),
  v4953 = (v4935 & i30) | (v3937 & ~i30),
  v4954 = (v4961 & i20) | (v4955 & ~i20),
  v4955 = (v4956 & i21) | (v4932 & ~i21),
  v4956 = (v4957 & i22) | (v4938 & ~i22),
  v4957 = (v4958 & i25) | (v4942 & ~i25),
  v4958 = (v3953 & i26) | (v4959 & ~i26),
  v4959 = (v3953 & i27) | (v4960 & ~i27),
  v4960 = (v4935 & i30) | (v3954 & ~i30),
  v4961 = (v4962 & i21) | (v4932 & ~i21),
  v4962 = (v4963 & i22) | (v4938 & ~i22),
  v4963 = (v4964 & i25) | (v4942 & ~i25),
  v4964 = (v3971 & i26) | (v4965 & ~i26),
  v4965 = (v3971 & i27) | (v4966 & ~i27),
  v4966 = (v4935 & i30) | (v3972 & ~i30),
  v4967 = (v4981 & i19) | (v4968 & ~i19),
  v4968 = (v4975 & i20) | (v4969 & ~i20),
  v4969 = (v4970 & i21) | (v4932 & ~i21),
  v4970 = (v4971 & i22) | (v4938 & ~i22),
  v4971 = (v4972 & i25) | (v4942 & ~i25),
  v4972 = (v3990 & i26) | (v4973 & ~i26),
  v4973 = (v3990 & i27) | (v4974 & ~i27),
  v4974 = (v4935 & i30) | (v3991 & ~i30),
  v4975 = (v4976 & i21) | (v4932 & ~i21),
  v4976 = (v4977 & i22) | (v4938 & ~i22),
  v4977 = (v4978 & i25) | (v4942 & ~i25),
  v4978 = (v4007 & i26) | (v4979 & ~i26),
  v4979 = (v4007 & i27) | (v4980 & ~i27),
  v4980 = (v4935 & i30) | (v4008 & ~i30),
  v4981 = (v4982 & i21) | (v4932 & ~i21),
  v4982 = (v4983 & i22) | (v4938 & ~i22),
  v4983 = (v4984 & i25) | (v4942 & ~i25),
  v4984 = (v4024 & i26) | (v4985 & ~i26),
  v4985 = (v4024 & i27) | (v4986 & ~i27),
  v4986 = (v4935 & i30) | (v4025 & ~i30),
  v4987 = (v5015 & i17) | (v4988 & ~i17),
  v4988 = (v5002 & i19) | (v4989 & ~i19),
  v4989 = (v4996 & i20) | (v4990 & ~i20),
  v4990 = (v4991 & i21) | (v4932 & ~i21),
  v4991 = (v4992 & i22) | (v4938 & ~i22),
  v4992 = (v4993 & i25) | (v4942 & ~i25),
  v4993 = (v4038 & i26) | (v4994 & ~i26),
  v4994 = (v4038 & i27) | (v4995 & ~i27),
  v4995 = (v4935 & i30) | (v4039 & ~i30),
  v4996 = (v4997 & i21) | (v4932 & ~i21),
  v4997 = (v4998 & i22) | (v4938 & ~i22),
  v4998 = (v4999 & i25) | (v4942 & ~i25),
  v4999 = (v4051 & i26) | (v5000 & ~i26),
  v5000 = (v4051 & i27) | (v5001 & ~i27),
  v5001 = (v4935 & i30) | (v4052 & ~i30),
  v5002 = (v5009 & i20) | (v5003 & ~i20),
  v5003 = (v5004 & i21) | (v4932 & ~i21),
  v5004 = (v5005 & i22) | (v4938 & ~i22),
  v5005 = (v5006 & i25) | (v4942 & ~i25),
  v5006 = (v4065 & i26) | (v5007 & ~i26),
  v5007 = (v4065 & i27) | (v5008 & ~i27),
  v5008 = (v4935 & i30) | (v4066 & ~i30),
  v5009 = (v5010 & i21) | (v4932 & ~i21),
  v5010 = (v5011 & i22) | (v4938 & ~i22),
  v5011 = (v5012 & i25) | (v4942 & ~i25),
  v5012 = (v4082 & i26) | (v5013 & ~i26),
  v5013 = (v4082 & i27) | (v5014 & ~i27),
  v5014 = (v4935 & i30) | (v4083 & ~i30),
  v5015 = (v5029 & i19) | (v5016 & ~i19),
  v5016 = (v5023 & i20) | (v5017 & ~i20),
  v5017 = (v5018 & i21) | (v4932 & ~i21),
  v5018 = (v5019 & i22) | (v4938 & ~i22),
  v5019 = (v5020 & i25) | (v4942 & ~i25),
  v5020 = (v4101 & i26) | (v5021 & ~i26),
  v5021 = (v4101 & i27) | (v5022 & ~i27),
  v5022 = (v4935 & i30) | (v4102 & ~i30),
  v5023 = (v5024 & i21) | (v4932 & ~i21),
  v5024 = (v5025 & i22) | (v4938 & ~i22),
  v5025 = (v5026 & i25) | (v4942 & ~i25),
  v5026 = (v4118 & i26) | (v5027 & ~i26),
  v5027 = (v4118 & i27) | (v5028 & ~i27),
  v5028 = (v4935 & i30) | (v4119 & ~i30),
  v5029 = (v5030 & i21) | (v4932 & ~i21),
  v5030 = (v5031 & i22) | (v4938 & ~i22),
  v5031 = (v5032 & i25) | (v4942 & ~i25),
  v5032 = (v4135 & i26) | (v5033 & ~i26),
  v5033 = (v4135 & i27) | (v5034 & ~i27),
  v5034 = (v4935 & i30) | (v4136 & ~i30),
  v5035 = (v5084 & i16) | (v5036 & ~i16),
  v5036 = (v5064 & i17) | (v5037 & ~i17),
  v5037 = (v5051 & i19) | (v5038 & ~i19),
  v5038 = (v5045 & i20) | (v5039 & ~i20),
  v5039 = (v5040 & i21) | (v4932 & ~i21),
  v5040 = (v5041 & i22) | (v4938 & ~i22),
  v5041 = (v5042 & i25) | (v4942 & ~i25),
  v5042 = (v4150 & i26) | (v5043 & ~i26),
  v5043 = (v4150 & i27) | (v5044 & ~i27),
  v5044 = (v4935 & i30) | (v4151 & ~i30),
  v5045 = (v5046 & i21) | (v4932 & ~i21),
  v5046 = (v5047 & i22) | (v4938 & ~i22),
  v5047 = (v5048 & i25) | (v4942 & ~i25),
  v5048 = (v4159 & i26) | (v5049 & ~i26),
  v5049 = (v4159 & i27) | (v5050 & ~i27),
  v5050 = (v4935 & i30) | (v4160 & ~i30),
  v5051 = (v5058 & i20) | (v5052 & ~i20),
  v5052 = (v5053 & i21) | (v4932 & ~i21),
  v5053 = (v5054 & i22) | (v4938 & ~i22),
  v5054 = (v5055 & i25) | (v4942 & ~i25),
  v5055 = (v4169 & i26) | (v5056 & ~i26),
  v5056 = (v4169 & i27) | (v5057 & ~i27),
  v5057 = (v4935 & i30) | (v4170 & ~i30),
  v5058 = (v5059 & i21) | (v4932 & ~i21),
  v5059 = (v5060 & i22) | (v4938 & ~i22),
  v5060 = (v5061 & i25) | (v4942 & ~i25),
  v5061 = (v4177 & i26) | (v5062 & ~i26),
  v5062 = (v4177 & i27) | (v5063 & ~i27),
  v5063 = (v4935 & i30) | (v4178 & ~i30),
  v5064 = (v5078 & i19) | (v5065 & ~i19),
  v5065 = (v5072 & i20) | (v5066 & ~i20),
  v5066 = (v5067 & i21) | (v4932 & ~i21),
  v5067 = (v5068 & i22) | (v4938 & ~i22),
  v5068 = (v5069 & i25) | (v4942 & ~i25),
  v5069 = (v4187 & i26) | (v5070 & ~i26),
  v5070 = (v4187 & i27) | (v5071 & ~i27),
  v5071 = (v4935 & i30) | (v4188 & ~i30),
  v5072 = (v5073 & i21) | (v4932 & ~i21),
  v5073 = (v5074 & i22) | (v4938 & ~i22),
  v5074 = (v5075 & i25) | (v4942 & ~i25),
  v5075 = (v4195 & i26) | (v5076 & ~i26),
  v5076 = (v4195 & i27) | (v5077 & ~i27),
  v5077 = (v4935 & i30) | (v4196 & ~i30),
  v5078 = (v5079 & i21) | (v4932 & ~i21),
  v5079 = (v5080 & i22) | (v4938 & ~i22),
  v5080 = (v5081 & i25) | (v4942 & ~i25),
  v5081 = (v4203 & i26) | (v5082 & ~i26),
  v5082 = (v4203 & i27) | (v5083 & ~i27),
  v5083 = (v4935 & i30) | (v4204 & ~i30),
  v5084 = (v5112 & i17) | (v5085 & ~i17),
  v5085 = (v5099 & i19) | (v5086 & ~i19),
  v5086 = (v5093 & i20) | (v5087 & ~i20),
  v5087 = (v5088 & i21) | (v4932 & ~i21),
  v5088 = (v5089 & i22) | (v4938 & ~i22),
  v5089 = (v5090 & i25) | (v4942 & ~i25),
  v5090 = (v4212 & i26) | (v5091 & ~i26),
  v5091 = (v4212 & i27) | (v5092 & ~i27),
  v5092 = (v4935 & i30) | (v4213 & ~i30),
  v5093 = (v5094 & i21) | (v4932 & ~i21),
  v5094 = (v5095 & i22) | (v4938 & ~i22),
  v5095 = (v5096 & i25) | (v4942 & ~i25),
  v5096 = (v4221 & i26) | (v5097 & ~i26),
  v5097 = (v4221 & i27) | (v5098 & ~i27),
  v5098 = (v4935 & i30) | (v4222 & ~i30),
  v5099 = (v5106 & i20) | (v5100 & ~i20),
  v5100 = (v5101 & i21) | (v4932 & ~i21),
  v5101 = (v5102 & i22) | (v4938 & ~i22),
  v5102 = (v5103 & i25) | (v4942 & ~i25),
  v5103 = (v4231 & i26) | (v5104 & ~i26),
  v5104 = (v4231 & i27) | (v5105 & ~i27),
  v5105 = (v4935 & i30) | (v4232 & ~i30),
  v5106 = (v5107 & i21) | (v4932 & ~i21),
  v5107 = (v5108 & i22) | (v4938 & ~i22),
  v5108 = (v5109 & i25) | (v4942 & ~i25),
  v5109 = (v4239 & i26) | (v5110 & ~i26),
  v5110 = (v4239 & i27) | (v5111 & ~i27),
  v5111 = (v4935 & i30) | (v4240 & ~i30),
  v5112 = (v5126 & i19) | (v5113 & ~i19),
  v5113 = (v5120 & i20) | (v5114 & ~i20),
  v5114 = (v5115 & i21) | (v4932 & ~i21),
  v5115 = (v5116 & i22) | (v4938 & ~i22),
  v5116 = (v5117 & i25) | (v4942 & ~i25),
  v5117 = (v4249 & i26) | (v5118 & ~i26),
  v5118 = (v4249 & i27) | (v5119 & ~i27),
  v5119 = (v4935 & i30) | (v4250 & ~i30),
  v5120 = (v5121 & i21) | (v4932 & ~i21),
  v5121 = (v5122 & i22) | (v4938 & ~i22),
  v5122 = (v5123 & i25) | (v4942 & ~i25),
  v5123 = (v4257 & i26) | (v5124 & ~i26),
  v5124 = (v4257 & i27) | (v5125 & ~i27),
  v5125 = (v4935 & i30) | (v4258 & ~i30),
  v5126 = (v5127 & i21) | (v4932 & ~i21),
  v5127 = (v5128 & i22) | (v4938 & ~i22),
  v5128 = (v5129 & i25) | (v4942 & ~i25),
  v5129 = (v4265 & i26) | (v5130 & ~i26),
  v5130 = (v4265 & i27) | (v5131 & ~i27),
  v5131 = (v4935 & i30) | (v4266 & ~i30),
  v5132 = (v5205 & i15) | (v5133 & ~i15),
  v5133 = (v5171 & i16) | (v5134 & ~i16),
  v5134 = (v5157 & i17) | (v5135 & ~i17),
  v5135 = (v5148 & i19) | (v5136 & ~i19),
  v5136 = (v5144 & i20) | (v5137 & ~i20),
  v5137 = (v5139 & i21) | (v5138 & ~i21),
  v5138 = (v4934 & i27) | (v27 & ~i27),
  v5139 = (v5141 & i22) | (v5140 & ~i22),
  v5140 = (v4940 & i27) | (v3908 & ~i27),
  v5141 = (v5143 & i25) | (v5142 & ~i25),
  v5142 = (v4944 & i27) | (v3912 & ~i27),
  v5143 = (v4947 & i27) | (v3920 & ~i27),
  v5144 = (v5145 & i21) | (v5138 & ~i21),
  v5145 = (v5146 & i22) | (v5140 & ~i22),
  v5146 = (v5147 & i25) | (v5142 & ~i25),
  v5147 = (v4953 & i27) | (v3936 & ~i27),
  v5148 = (v5153 & i20) | (v5149 & ~i20),
  v5149 = (v5150 & i21) | (v5138 & ~i21),
  v5150 = (v5151 & i22) | (v5140 & ~i22),
  v5151 = (v5152 & i25) | (v5142 & ~i25),
  v5152 = (v4960 & i27) | (v3953 & ~i27),
  v5153 = (v5154 & i21) | (v5138 & ~i21),
  v5154 = (v5155 & i22) | (v5140 & ~i22),
  v5155 = (v5156 & i25) | (v5142 & ~i25),
  v5156 = (v4966 & i27) | (v3971 & ~i27),
  v5157 = (v5167 & i19) | (v5158 & ~i19),
  v5158 = (v5163 & i20) | (v5159 & ~i20),
  v5159 = (v5160 & i21) | (v5138 & ~i21),
  v5160 = (v5161 & i22) | (v5140 & ~i22),
  v5161 = (v5162 & i25) | (v5142 & ~i25),
  v5162 = (v4974 & i27) | (v3990 & ~i27),
  v5163 = (v5164 & i21) | (v5138 & ~i21),
  v5164 = (v5165 & i22) | (v5140 & ~i22),
  v5165 = (v5166 & i25) | (v5142 & ~i25),
  v5166 = (v4980 & i27) | (v4007 & ~i27),
  v5167 = (v5168 & i21) | (v5138 & ~i21),
  v5168 = (v5169 & i22) | (v5140 & ~i22),
  v5169 = (v5170 & i25) | (v5142 & ~i25),
  v5170 = (v4986 & i27) | (v4024 & ~i27),
  v5171 = (v5191 & i17) | (v5172 & ~i17),
  v5172 = (v5182 & i19) | (v5173 & ~i19),
  v5173 = (v5178 & i20) | (v5174 & ~i20),
  v5174 = (v5175 & i21) | (v5138 & ~i21),
  v5175 = (v5176 & i22) | (v5140 & ~i22),
  v5176 = (v5177 & i25) | (v5142 & ~i25),
  v5177 = (v4995 & i27) | (v4038 & ~i27),
  v5178 = (v5179 & i21) | (v5138 & ~i21),
  v5179 = (v5180 & i22) | (v5140 & ~i22),
  v5180 = (v5181 & i25) | (v5142 & ~i25),
  v5181 = (v5001 & i27) | (v4051 & ~i27),
  v5182 = (v5187 & i20) | (v5183 & ~i20),
  v5183 = (v5184 & i21) | (v5138 & ~i21),
  v5184 = (v5185 & i22) | (v5140 & ~i22),
  v5185 = (v5186 & i25) | (v5142 & ~i25),
  v5186 = (v5008 & i27) | (v4065 & ~i27),
  v5187 = (v5188 & i21) | (v5138 & ~i21),
  v5188 = (v5189 & i22) | (v5140 & ~i22),
  v5189 = (v5190 & i25) | (v5142 & ~i25),
  v5190 = (v5014 & i27) | (v4082 & ~i27),
  v5191 = (v5201 & i19) | (v5192 & ~i19),
  v5192 = (v5197 & i20) | (v5193 & ~i20),
  v5193 = (v5194 & i21) | (v5138 & ~i21),
  v5194 = (v5195 & i22) | (v5140 & ~i22),
  v5195 = (v5196 & i25) | (v5142 & ~i25),
  v5196 = (v5022 & i27) | (v4101 & ~i27),
  v5197 = (v5198 & i21) | (v5138 & ~i21),
  v5198 = (v5199 & i22) | (v5140 & ~i22),
  v5199 = (v5200 & i25) | (v5142 & ~i25),
  v5200 = (v5028 & i27) | (v4118 & ~i27),
  v5201 = (v5202 & i21) | (v5138 & ~i21),
  v5202 = (v5203 & i22) | (v5140 & ~i22),
  v5203 = (v5204 & i25) | (v5142 & ~i25),
  v5204 = (v5034 & i27) | (v4135 & ~i27),
  v5205 = (v5240 & i16) | (v5206 & ~i16),
  v5206 = (v5226 & i17) | (v5207 & ~i17),
  v5207 = (v5217 & i19) | (v5208 & ~i19),
  v5208 = (v5213 & i20) | (v5209 & ~i20),
  v5209 = (v5210 & i21) | (v5138 & ~i21),
  v5210 = (v5211 & i22) | (v5140 & ~i22),
  v5211 = (v5212 & i25) | (v5142 & ~i25),
  v5212 = (v5044 & i27) | (v4150 & ~i27),
  v5213 = (v5214 & i21) | (v5138 & ~i21),
  v5214 = (v5215 & i22) | (v5140 & ~i22),
  v5215 = (v5216 & i25) | (v5142 & ~i25),
  v5216 = (v5050 & i27) | (v4159 & ~i27),
  v5217 = (v5222 & i20) | (v5218 & ~i20),
  v5218 = (v5219 & i21) | (v5138 & ~i21),
  v5219 = (v5220 & i22) | (v5140 & ~i22),
  v5220 = (v5221 & i25) | (v5142 & ~i25),
  v5221 = (v5057 & i27) | (v4169 & ~i27),
  v5222 = (v5223 & i21) | (v5138 & ~i21),
  v5223 = (v5224 & i22) | (v5140 & ~i22),
  v5224 = (v5225 & i25) | (v5142 & ~i25),
  v5225 = (v5063 & i27) | (v4177 & ~i27),
  v5226 = (v5236 & i19) | (v5227 & ~i19),
  v5227 = (v5232 & i20) | (v5228 & ~i20),
  v5228 = (v5229 & i21) | (v5138 & ~i21),
  v5229 = (v5230 & i22) | (v5140 & ~i22),
  v5230 = (v5231 & i25) | (v5142 & ~i25),
  v5231 = (v5071 & i27) | (v4187 & ~i27),
  v5232 = (v5233 & i21) | (v5138 & ~i21),
  v5233 = (v5234 & i22) | (v5140 & ~i22),
  v5234 = (v5235 & i25) | (v5142 & ~i25),
  v5235 = (v5077 & i27) | (v4195 & ~i27),
  v5236 = (v5237 & i21) | (v5138 & ~i21),
  v5237 = (v5238 & i22) | (v5140 & ~i22),
  v5238 = (v5239 & i25) | (v5142 & ~i25),
  v5239 = (v5083 & i27) | (v4203 & ~i27),
  v5240 = (v5260 & i17) | (v5241 & ~i17),
  v5241 = (v5251 & i19) | (v5242 & ~i19),
  v5242 = (v5247 & i20) | (v5243 & ~i20),
  v5243 = (v5244 & i21) | (v5138 & ~i21),
  v5244 = (v5245 & i22) | (v5140 & ~i22),
  v5245 = (v5246 & i25) | (v5142 & ~i25),
  v5246 = (v5092 & i27) | (v4212 & ~i27),
  v5247 = (v5248 & i21) | (v5138 & ~i21),
  v5248 = (v5249 & i22) | (v5140 & ~i22),
  v5249 = (v5250 & i25) | (v5142 & ~i25),
  v5250 = (v5098 & i27) | (v4221 & ~i27),
  v5251 = (v5256 & i20) | (v5252 & ~i20),
  v5252 = (v5253 & i21) | (v5138 & ~i21),
  v5253 = (v5254 & i22) | (v5140 & ~i22),
  v5254 = (v5255 & i25) | (v5142 & ~i25),
  v5255 = (v5105 & i27) | (v4231 & ~i27),
  v5256 = (v5257 & i21) | (v5138 & ~i21),
  v5257 = (v5258 & i22) | (v5140 & ~i22),
  v5258 = (v5259 & i25) | (v5142 & ~i25),
  v5259 = (v5111 & i27) | (v4239 & ~i27),
  v5260 = (v5270 & i19) | (v5261 & ~i19),
  v5261 = (v5266 & i20) | (v5262 & ~i20),
  v5262 = (v5263 & i21) | (v5138 & ~i21),
  v5263 = (v5264 & i22) | (v5140 & ~i22),
  v5264 = (v5265 & i25) | (v5142 & ~i25),
  v5265 = (v5119 & i27) | (v4249 & ~i27),
  v5266 = (v5267 & i21) | (v5138 & ~i21),
  v5267 = (v5268 & i22) | (v5140 & ~i22),
  v5268 = (v5269 & i25) | (v5142 & ~i25),
  v5269 = (v5125 & i27) | (v4257 & ~i27),
  v5270 = (v5271 & i21) | (v5138 & ~i21),
  v5271 = (v5272 & i22) | (v5140 & ~i22),
  v5272 = (v5273 & i25) | (v5142 & ~i25),
  v5273 = (v5131 & i27) | (v4265 & ~i27),
  v5274 = (v3901 & i12) | (v5275 & ~i12),
  v5275 = (v3901 & i13) | (v5276 & ~i13),
  v5276 = (v5277 & i14) | (v3901 & ~i14),
  v5277 = (v5350 & i15) | (v5278 & ~i15),
  v5278 = (v5316 & i16) | (v5279 & ~i16),
  v5279 = (v5302 & i17) | (v5280 & ~i17),
  v5280 = (v5293 & i19) | (v5281 & ~i19),
  v5281 = (v5289 & i20) | (v5282 & ~i20),
  v5282 = (v5284 & i21) | (v5283 & ~i21),
  v5283 = (v4933 & i26) | (v27 & ~i26),
  v5284 = (v5286 & i22) | (v5285 & ~i22),
  v5285 = (v4939 & i26) | (v3908 & ~i26),
  v5286 = (v5288 & i25) | (v5287 & ~i25),
  v5287 = (v4943 & i26) | (v3912 & ~i26),
  v5288 = (v4946 & i26) | (v3920 & ~i26),
  v5289 = (v5290 & i21) | (v5283 & ~i21),
  v5290 = (v5291 & i22) | (v5285 & ~i22),
  v5291 = (v5292 & i25) | (v5287 & ~i25),
  v5292 = (v4952 & i26) | (v3936 & ~i26),
  v5293 = (v5298 & i20) | (v5294 & ~i20),
  v5294 = (v5295 & i21) | (v5283 & ~i21),
  v5295 = (v5296 & i22) | (v5285 & ~i22),
  v5296 = (v5297 & i25) | (v5287 & ~i25),
  v5297 = (v4959 & i26) | (v3953 & ~i26),
  v5298 = (v5299 & i21) | (v5283 & ~i21),
  v5299 = (v5300 & i22) | (v5285 & ~i22),
  v5300 = (v5301 & i25) | (v5287 & ~i25),
  v5301 = (v4965 & i26) | (v3971 & ~i26),
  v5302 = (v5312 & i19) | (v5303 & ~i19),
  v5303 = (v5308 & i20) | (v5304 & ~i20),
  v5304 = (v5305 & i21) | (v5283 & ~i21),
  v5305 = (v5306 & i22) | (v5285 & ~i22),
  v5306 = (v5307 & i25) | (v5287 & ~i25),
  v5307 = (v4973 & i26) | (v3990 & ~i26),
  v5308 = (v5309 & i21) | (v5283 & ~i21),
  v5309 = (v5310 & i22) | (v5285 & ~i22),
  v5310 = (v5311 & i25) | (v5287 & ~i25),
  v5311 = (v4979 & i26) | (v4007 & ~i26),
  v5312 = (v5313 & i21) | (v5283 & ~i21),
  v5313 = (v5314 & i22) | (v5285 & ~i22),
  v5314 = (v5315 & i25) | (v5287 & ~i25),
  v5315 = (v4985 & i26) | (v4024 & ~i26),
  v5316 = (v5336 & i17) | (v5317 & ~i17),
  v5317 = (v5327 & i19) | (v5318 & ~i19),
  v5318 = (v5323 & i20) | (v5319 & ~i20),
  v5319 = (v5320 & i21) | (v5283 & ~i21),
  v5320 = (v5321 & i22) | (v5285 & ~i22),
  v5321 = (v5322 & i25) | (v5287 & ~i25),
  v5322 = (v4994 & i26) | (v4038 & ~i26),
  v5323 = (v5324 & i21) | (v5283 & ~i21),
  v5324 = (v5325 & i22) | (v5285 & ~i22),
  v5325 = (v5326 & i25) | (v5287 & ~i25),
  v5326 = (v5000 & i26) | (v4051 & ~i26),
  v5327 = (v5332 & i20) | (v5328 & ~i20),
  v5328 = (v5329 & i21) | (v5283 & ~i21),
  v5329 = (v5330 & i22) | (v5285 & ~i22),
  v5330 = (v5331 & i25) | (v5287 & ~i25),
  v5331 = (v5007 & i26) | (v4065 & ~i26),
  v5332 = (v5333 & i21) | (v5283 & ~i21),
  v5333 = (v5334 & i22) | (v5285 & ~i22),
  v5334 = (v5335 & i25) | (v5287 & ~i25),
  v5335 = (v5013 & i26) | (v4082 & ~i26),
  v5336 = (v5346 & i19) | (v5337 & ~i19),
  v5337 = (v5342 & i20) | (v5338 & ~i20),
  v5338 = (v5339 & i21) | (v5283 & ~i21),
  v5339 = (v5340 & i22) | (v5285 & ~i22),
  v5340 = (v5341 & i25) | (v5287 & ~i25),
  v5341 = (v5021 & i26) | (v4101 & ~i26),
  v5342 = (v5343 & i21) | (v5283 & ~i21),
  v5343 = (v5344 & i22) | (v5285 & ~i22),
  v5344 = (v5345 & i25) | (v5287 & ~i25),
  v5345 = (v5027 & i26) | (v4118 & ~i26),
  v5346 = (v5347 & i21) | (v5283 & ~i21),
  v5347 = (v5348 & i22) | (v5285 & ~i22),
  v5348 = (v5349 & i25) | (v5287 & ~i25),
  v5349 = (v5033 & i26) | (v4135 & ~i26),
  v5350 = (v5385 & i16) | (v5351 & ~i16),
  v5351 = (v5371 & i17) | (v5352 & ~i17),
  v5352 = (v5362 & i19) | (v5353 & ~i19),
  v5353 = (v5358 & i20) | (v5354 & ~i20),
  v5354 = (v5355 & i21) | (v5283 & ~i21),
  v5355 = (v5356 & i22) | (v5285 & ~i22),
  v5356 = (v5357 & i25) | (v5287 & ~i25),
  v5357 = (v5043 & i26) | (v4150 & ~i26),
  v5358 = (v5359 & i21) | (v5283 & ~i21),
  v5359 = (v5360 & i22) | (v5285 & ~i22),
  v5360 = (v5361 & i25) | (v5287 & ~i25),
  v5361 = (v5049 & i26) | (v4159 & ~i26),
  v5362 = (v5367 & i20) | (v5363 & ~i20),
  v5363 = (v5364 & i21) | (v5283 & ~i21),
  v5364 = (v5365 & i22) | (v5285 & ~i22),
  v5365 = (v5366 & i25) | (v5287 & ~i25),
  v5366 = (v5056 & i26) | (v4169 & ~i26),
  v5367 = (v5368 & i21) | (v5283 & ~i21),
  v5368 = (v5369 & i22) | (v5285 & ~i22),
  v5369 = (v5370 & i25) | (v5287 & ~i25),
  v5370 = (v5062 & i26) | (v4177 & ~i26),
  v5371 = (v5381 & i19) | (v5372 & ~i19),
  v5372 = (v5377 & i20) | (v5373 & ~i20),
  v5373 = (v5374 & i21) | (v5283 & ~i21);
always begin
  i2 = \[434] ;
  i3 = \[433] ;
  i4 = \[432] ;
  i5 = \[431] ;
  i6 = \[430] ;
  i7 = \[429] ;
  i8 = \[428] ;
  i9 = \[427] ;
  i10 = \[426] ;
  i11 = \[425] ;
  i12 = \[424] ;
  i13 = \[423] ;
  i14 = \[422] ;
  i29 = \[421] ;
  i30 = \[420] ;
  i31 = \[419] ;
  i32 = \[418] ;
  i33 = \[417] ;
  i34 = \[416] ;
  i35 = \[415] ;
  i36 = \[414] ;
  i37 = \[413] ;
  i38 = \[412] ;
  i39 = \[411] ;
  i40 = \[410] ;
  i41 = \[409] ;
  i42 = \[408] ;
  i43 = \[407] ;
  i44 = \[406] ;
  i45 = \[405] ;
  i46 = \[404] ;
  i47 = \[403] ;
  i48 = \[402] ;
end
initial begin
  i2 = 0;
  i3 = 0;
  i4 = 0;
  i5 = 0;
  i6 = 0;
  i7 = 0;
  i8 = 0;
  i9 = 0;
  i10 = 0;
  i11 = 0;
  i12 = 0;
  i13 = 0;
  i14 = 0;
  i29 = 0;
  i30 = 0;
  i31 = 0;
  i32 = 0;
  i33 = 0;
  i34 = 0;
  i35 = 0;
  i36 = 0;
  i37 = 0;
  i38 = 0;
  i39 = 0;
  i40 = 0;
  i41 = 0;
  i42 = 0;
  i43 = 0;
  i44 = 0;
  i45 = 0;
  i46 = 0;
  i47 = 0;
  i48 = 0;
end
endmodule

