// IWLS benchmark module "unreg" printed on Wed May 29 17:30:25 2002
module unreg(a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, s, t, u, v, w, \xx , y, z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0, o0, p0, q0, r0, s0, t0, u0, v0, w0, x0, y0, z0, a1);
input
  g0,
  h0,
  i0,
  j0,
  k0,
  a,
  b,
  c,
  d,
  e,
  f,
  g,
  h,
  i,
  j,
  k,
  l,
  m,
  n,
  o,
  p,
  q,
  s,
  t,
  u,
  v,
  w,
  \xx ,
  y,
  z,
  a0,
  b0,
  c0,
  d0,
  e0,
  f0;
output
  l0,
  m0,
  n0,
  o0,
  p0,
  q0,
  r0,
  s0,
  t0,
  u0,
  v0,
  w0,
  x0,
  y0,
  z0,
  a1;
wire
  g2,
  i2,
  j2,
  \[10] ,
  \[11] ,
  m2,
  \[12] ,
  \[13] ,
  o2,
  \[14] ,
  \[0] ,
  \[15] ,
  q2,
  \[1] ,
  r2,
  \[2] ,
  \[3] ,
  \[4] ,
  u2,
  \[5] ,
  \[6] ,
  w1,
  w2,
  \[7] ,
  \[8] ,
  y1,
  y2,
  \[9] ,
  z2,
  a2,
  b2,
  e2;
assign
  g2 = (b0 & t) | ((~t & ~g) | s),
  i2 = (c0 & t) | ((~t & ~f) | s),
  j2 = (v & t) | ((~t & ~e) | s),
  \[10]  = (~u & ~f0) | (u & ~q2),
  l0 = \[0] ,
  \[11]  = (~u & ~g0) | (u & ~r2),
  m0 = \[1] ,
  m2 = (e0 & t) | ((~t & ~l) | s),
  \[12]  = (~u & ~h0) | (u & ~u2),
  n0 = \[2] ,
  \[13]  = (~u & ~i0) | (u & ~w2),
  o0 = \[3] ,
  o2 = (f0 & t) | ((~t & ~k) | s),
  \[14]  = (~u & ~j0) | (u & ~y2),
  p0 = \[4] ,
  \[0]  = (~u & ~v) | (u & ~w1),
  \[15]  = (~u & ~k0) | (u & ~z2),
  q0 = \[5] ,
  q2 = (g0 & t) | ((~t & ~j) | s),
  \[1]  = (~u & ~w) | (u & ~y1),
  r0 = \[6] ,
  r2 = (z & t) | ((~t & ~i) | s),
  \[2]  = (~u & ~\xx ) | (u & ~a2),
  s0 = \[7] ,
  \[3]  = (~u & ~y) | (u & ~b2),
  t0 = \[8] ,
  \[4]  = (~u & ~z) | (u & ~e2),
  u0 = \[9] ,
  u2 = (i0 & t) | ((~t & ~p) | s),
  \[5]  = (~u & ~a0) | (u & ~g2),
  v0 = \[10] ,
  \[6]  = (~u & ~b0) | (u & ~i2),
  w0 = \[11] ,
  w1 = (w & t) | ((~t & ~d) | s),
  w2 = (j0 & t) | ((~t & ~o) | s),
  \[7]  = (~u & ~c0) | (u & ~j2),
  x0 = \[12] ,
  \[8]  = (~u & ~d0) | (u & ~m2),
  y0 = \[13] ,
  y1 = (\xx  & t) | ((~t & ~c) | s),
  y2 = (k0 & t) | ((~t & ~n) | s),
  \[9]  = (~u & ~e0) | (u & ~o2),
  z0 = \[14] ,
  z2 = (d0 & t) | ((~t & ~m) | s),
  a1 = \[15] ,
  a2 = (y & t) | ((~t & ~b) | s),
  b2 = (~t & ~a) | ((t & ~q) | s),
  e2 = (a0 & t) | ((~t & ~h) | s);
endmodule

