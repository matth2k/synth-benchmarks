module s1238 (
  CK,
  G0,
  G1,
  G10,
  G11,
  G12,
  G13,
  G2,
  G3,
  G4,
  G5,
  G6,
  G7,
  G8,
  G9,
  G532,
  G546,
  G550,
  G547,
  G548,
  G535,
  G45,
  G551,
  G539,
  G530,
  G552,
  G549,
  G542,
  G537
);
  input CK;
  wire CK;
  input G0;
  wire G0;
  input G1;
  wire G1;
  input G10;
  wire G10;
  input G11;
  wire G11;
  input G12;
  wire G12;
  input G13;
  wire G13;
  input G2;
  wire G2;
  input G3;
  wire G3;
  input G4;
  wire G4;
  input G5;
  wire G5;
  input G6;
  wire G6;
  input G7;
  wire G7;
  input G8;
  wire G8;
  input G9;
  wire G9;
  output G532;
  wire G532;
  output G546;
  wire G546;
  output G550;
  wire G550;
  output G547;
  wire G547;
  output G548;
  wire G548;
  output G535;
  wire G535;
  output G45;
  wire G45;
  output G551;
  wire G551;
  output G539;
  wire G539;
  output G530;
  wire G530;
  output G552;
  wire G552;
  output G549;
  wire G549;
  output G542;
  wire G542;
  output G537;
  wire G537;
  wire __0__;
  wire __1__;
  wire __2__;
  wire __3__;
  wire __4__;
  wire __5__;
  wire __6__;
  wire __7__;
  wire __8__;
  wire __9__;
  wire __10__;
  wire __11__;
  wire __12__;
  wire __13__;
  wire __14__;
  wire __15__;
  wire __16__;
  wire __17__;
  wire __18__;
  wire __19__;
  wire __20__;
  wire __21__;
  wire __22__;
  wire __23__;
  wire __24__;
  wire __25__;
  wire __26__;
  wire __27__;
  wire __28__;
  wire __29__;
  wire __30__;
  wire __31__;
  wire __32__;
  wire __33__;
  wire __34__;
  wire __35__;
  wire __36__;
  wire __37__;
  wire __38__;
  wire __39__;
  wire __40__;
  wire __41__;
  wire __42__;
  wire __43__;
  wire __44__;
  wire __45__;
  wire __47__;
  wire __48__;
  wire __49__;
  wire __50__;
  wire __51__;
  wire __52__;
  wire __53__;
  wire __54__;
  wire __55__;
  wire __56__;
  wire __57__;
  wire __58__;
  wire __59__;
  wire __60__;
  wire __61__;
  wire __62__;
  wire __63__;
  wire __64__;
  wire __65__;
  wire __66__;
  wire __67__;
  wire __68__;
  wire __69__;
  wire __70__;
  wire __71__;
  wire __72__;
  wire __73__;
  wire __75__;
  wire __76__;
  wire __77__;
  wire __78__;
  wire __79__;
  wire __80__;
  wire __81__;
  wire __82__;
  wire __83__;
  wire __84__;
  wire __85__;
  wire __86__;
  wire __87__;
  wire __88__;
  wire __89__;
  wire __90__;
  wire __91__;
  wire __92__;
  wire __93__;
  wire __94__;
  wire __95__;
  wire __96__;
  wire __97__;
  wire __98__;
  wire __99__;
  wire __100__;
  wire __101__;
  wire __102__;
  wire __103__;
  wire __104__;
  wire __105__;
  wire __106__;
  wire __107__;
  wire __108__;
  wire __109__;
  wire __110__;
  wire __111__;
  wire __112__;
  wire __113__;
  wire __114__;
  wire __115__;
  wire __116__;
  wire __117__;
  wire __118__;
  wire __119__;
  wire __120__;
  wire __121__;
  wire __122__;
  wire __123__;
  wire __124__;
  wire __125__;
  wire __126__;
  wire __127__;
  wire __128__;
  wire __129__;
  wire __130__;
  wire __131__;
  wire __132__;
  wire __133__;
  wire __134__;
  wire __135__;
  wire __136__;
  wire __137__;
  wire __138__;
  wire __139__;
  wire __140__;
  wire __141__;
  wire __142__;
  wire __143__;
  wire __144__;
  wire __145__;
  wire __146__;
  wire __147__;
  wire __148__;
  wire __149__;
  wire __150__;
  INV __151__ (
    .I(__13__),
    .O(__0__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __152__ (
    .D(__93__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __153__ (
    .D(__129__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__2__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __154__ (
    .D(__125__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__3__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __155__ (
    .D(__141__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__4__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __156__ (
    .D(__77__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__5__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __157__ (
    .D(__82__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__6__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __158__ (
    .D(__81__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__7__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __159__ (
    .D(__149__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__8__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __160__ (
    .D(__150__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__9__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __161__ (
    .D(__124__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__10__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __162__ (
    .D(__73__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__11__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __163__ (
    .D(__144__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__12__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __164__ (
    .D(__90__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__13__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __165__ (
    .D(__145__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__14__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __166__ (
    .D(__98__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__15__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __167__ (
    .D(__128__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__16__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __168__ (
    .D(__66__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__17__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __169__ (
    .D(__148__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__18__)
  );
  LUT4 #(
    .INIT(16'heff7)
  ) __170__ (
    .I3(G10),
    .I2(G9),
    .I1(G8),
    .I0(G7),
    .O(__19__)
  );
  LUT4 #(
    .INIT(16'h8000)
  ) __171__ (
    .I3(G6),
    .I2(G4),
    .I1(G5),
    .I0(G11),
    .O(__20__)
  );
  LUT5 #(
    .INIT(32'h00004f44)
  ) __172__ (
    .I4(G3),
    .I3(__20__),
    .I2(__19__),
    .I1(__5__),
    .I0(G6),
    .O(__21__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __173__ (
    .I1(G11),
    .I0(G5),
    .O(__22__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __174__ (
    .I2(G6),
    .I1(G3),
    .I0(G4),
    .O(__23__)
  );
  LUT6 #(
    .INIT(64'h1408000000000000)
  ) __175__ (
    .I5(__23__),
    .I4(__22__),
    .I3(G9),
    .I2(G10),
    .I1(G8),
    .I0(G7),
    .O(__24__)
  );
  LUT6 #(
    .INIT(64'h0000000000001000)
  ) __176__ (
    .I5(G10),
    .I4(G8),
    .I3(G9),
    .I2(G5),
    .I1(G7),
    .I0(G11),
    .O(__25__)
  );
  LUT4 #(
    .INIT(16'h8000)
  ) __177__ (
    .I3(G6),
    .I2(G3),
    .I1(G4),
    .I0(__25__),
    .O(__26__)
  );
  LUT5 #(
    .INIT(32'h10000000)
  ) __178__ (
    .I4(G3),
    .I3(G11),
    .I2(__9__),
    .I1(G4),
    .I0(G5),
    .O(__27__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __179__ (
    .I1(G3),
    .I0(G5),
    .O(__28__)
  );
  LUT5 #(
    .INIT(32'h80000000)
  ) __180__ (
    .I4(G10),
    .I3(G9),
    .I2(G8),
    .I1(G7),
    .I0(G11),
    .O(__29__)
  );
  LUT6 #(
    .INIT(64'h1555555500000000)
  ) __181__ (
    .I5(G2),
    .I4(G6),
    .I3(G4),
    .I2(__29__),
    .I1(__28__),
    .I0(__27__),
    .O(__30__)
  );
  LUT6 #(
    .INIT(64'ha00000ff3f3f3f3f)
  ) __182__ (
    .I5(G7),
    .I4(G10),
    .I3(G9),
    .I2(G8),
    .I1(__11__),
    .I0(G11),
    .O(__31__)
  );
  LUT3 #(
    .INIT(8'h0d)
  ) __183__ (
    .I2(G13),
    .I1(__31__),
    .I0(__3__),
    .O(__32__)
  );
  LUT6 #(
    .INIT(64'hfe00fefe00000000)
  ) __184__ (
    .I5(__32__),
    .I4(__30__),
    .I3(__26__),
    .I2(G2),
    .I1(__24__),
    .I0(__21__),
    .O(__33__)
  );
  LUT5 #(
    .INIT(32'h7ff0c2a0)
  ) __185__ (
    .I4(G4),
    .I3(G1),
    .I2(G0),
    .I1(G3),
    .I0(G5),
    .O(__34__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __186__ (
    .I1(G10),
    .I0(G8),
    .O(__35__)
  );
  LUT4 #(
    .INIT(16'hdfc0)
  ) __187__ (
    .I3(G7),
    .I2(G8),
    .I1(__10__),
    .I0(G6),
    .O(__36__)
  );
  LUT6 #(
    .INIT(64'h1111ff1f00000000)
  ) __188__ (
    .I5(G11),
    .I4(__36__),
    .I3(__35__),
    .I2(G9),
    .I1(G6),
    .I0(__11__),
    .O(__37__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __189__ (
    .I1(G8),
    .I0(__10__),
    .O(__38__)
  );
  LUT3 #(
    .INIT(8'h01)
  ) __190__ (
    .I2(G10),
    .I1(G9),
    .I0(G11),
    .O(__39__)
  );
  LUT3 #(
    .INIT(8'h40)
  ) __191__ (
    .I2(G7),
    .I1(__11__),
    .I0(G6),
    .O(__40__)
  );
  LUT4 #(
    .INIT(16'h0305)
  ) __192__ (
    .I3(G3),
    .I2(G4),
    .I1(G0),
    .I0(G5),
    .O(__41__)
  );
  LUT6 #(
    .INIT(64'h0003000a00000000)
  ) __193__ (
    .I5(G9),
    .I4(G8),
    .I3(G7),
    .I2(G11),
    .I1(__10__),
    .I0(G10),
    .O(__42__)
  );
  LUT6 #(
    .INIT(64'h000000fb00000000)
  ) __194__ (
    .I5(__18__),
    .I4(__42__),
    .I3(__41__),
    .I2(__40__),
    .I1(__39__),
    .I0(__38__),
    .O(__43__)
  );
  LUT4 #(
    .INIT(16'h1000)
  ) __195__ (
    .I3(__43__),
    .I2(G12),
    .I1(G13),
    .I0(__37__),
    .O(__44__)
  );
  LUT6 #(
    .INIT(64'hff00000040404040)
  ) __196__ (
    .I5(G2),
    .I4(__44__),
    .I3(__34__),
    .I2(__21__),
    .I1(__33__),
    .I0(G12),
    .O(__45__)
  );
  LUT5 #(
    .INIT(32'h7ffeffff)
  ) __198__ (
    .I4(G9),
    .I3(G10),
    .I2(G8),
    .I1(G7),
    .I0(G11),
    .O(__47__)
  );
  LUT6 #(
    .INIT(64'h4000000000000000)
  ) __199__ (
    .I5(G6),
    .I4(G2),
    .I3(G4),
    .I2(G1),
    .I1(__28__),
    .I0(__47__),
    .O(__48__)
  );
  LUT4 #(
    .INIT(16'h1000)
  ) __200__ (
    .I3(G7),
    .I2(G11),
    .I1(G10),
    .I0(G9),
    .O(__49__)
  );
  LUT6 #(
    .INIT(64'h6001000000000000)
  ) __201__ (
    .I5(G3),
    .I4(__49__),
    .I3(G6),
    .I2(G8),
    .I1(G4),
    .I0(G1),
    .O(__50__)
  );
  LUT4 #(
    .INIT(16'h0080)
  ) __202__ (
    .I3(G10),
    .I2(G9),
    .I1(G8),
    .I0(G11),
    .O(__51__)
  );
  LUT4 #(
    .INIT(16'h0080)
  ) __203__ (
    .I3(G8),
    .I2(G10),
    .I1(G9),
    .I0(G11),
    .O(__52__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __204__ (
    .I1(G6),
    .I0(G3),
    .O(__53__)
  );
  LUT6 #(
    .INIT(64'h00005a4000005040)
  ) __205__ (
    .I5(__53__),
    .I4(G7),
    .I3(__52__),
    .I2(__23__),
    .I1(__51__),
    .I0(G1),
    .O(__54__)
  );
  LUT5 #(
    .INIT(32'h55015555)
  ) __206__ (
    .I4(G2),
    .I3(G5),
    .I2(__54__),
    .I1(__50__),
    .I0(__48__),
    .O(__55__)
  );
  LUT6 #(
    .INIT(64'h8000000000000000)
  ) __207__ (
    .I5(G6),
    .I4(G3),
    .I3(G4),
    .I2(G5),
    .I1(G0),
    .I0(__29__),
    .O(__56__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __208__ (
    .I1(G3),
    .I0(G5),
    .O(__57__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __209__ (
    .I1(G6),
    .I0(G9),
    .O(__58__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __210__ (
    .I1(G10),
    .I0(G8),
    .O(__59__)
  );
  LUT6 #(
    .INIT(64'h4000000000000000)
  ) __211__ (
    .I5(G8),
    .I4(G7),
    .I3(G3),
    .I2(G5),
    .I1(__8__),
    .I0(G10),
    .O(__60__)
  );
  LUT3 #(
    .INIT(8'h04)
  ) __212__ (
    .I2(G4),
    .I1(G11),
    .I0(G0),
    .O(__61__)
  );
  LUT6 #(
    .INIT(64'hffff400000000000)
  ) __213__ (
    .I5(__61__),
    .I4(__60__),
    .I3(__59__),
    .I2(__58__),
    .I1(__57__),
    .I0(G7),
    .O(__62__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __214__ (
    .I1(G2),
    .I0(G1),
    .O(__63__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __215__ (
    .I1(G12),
    .I0(G13),
    .O(__64__)
  );
  LUT6 #(
    .INIT(64'hcf8a000000000000)
  ) __216__ (
    .I5(__64__),
    .I4(__63__),
    .I3(__62__),
    .I2(__43__),
    .I1(__37__),
    .I0(__56__),
    .O(__65__)
  );
  LUT5 #(
    .INIT(32'hff00fff4)
  ) __217__ (
    .I4(G12),
    .I3(__65__),
    .I2(__33__),
    .I1(G13),
    .I0(__55__),
    .O(__66__)
  );
  LUT6 #(
    .INIT(64'h80575575005db37f)
  ) __218__ (
    .I5(G4),
    .I4(G5),
    .I3(G2),
    .I2(G3),
    .I1(G6),
    .I0(G1),
    .O(__67__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __219__ (
    .I1(__31__),
    .I0(__67__),
    .O(__68__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __220__ (
    .I1(G13),
    .I0(G12),
    .O(__69__)
  );
  LUT4 #(
    .INIT(16'h00d0)
  ) __221__ (
    .I3(G13),
    .I2(G12),
    .I1(__37__),
    .I0(__43__),
    .O(__70__)
  );
  LUT5 #(
    .INIT(32'h0000000d)
  ) __222__ (
    .I4(G12),
    .I3(G13),
    .I2(__33__),
    .I1(__31__),
    .I0(__3__),
    .O(__71__)
  );
  LUT6 #(
    .INIT(64'hffffffff40ff4040)
  ) __223__ (
    .I5(__71__),
    .I4(__70__),
    .I3(__65__),
    .I2(__55__),
    .I1(__69__),
    .I0(__68__),
    .O(__72__)
  );
  LUT3 #(
    .INIT(8'hf4)
  ) __224__ (
    .I2(G10),
    .I1(G11),
    .I0(G9),
    .O(__73__)
  );
  LUT6 #(
    .INIT(64'hc5ff10df33ffffff)
  ) __226__ (
    .I5(G6),
    .I4(G10),
    .I3(G9),
    .I2(G8),
    .I1(G7),
    .I0(G11),
    .O(__75__)
  );
  LUT6 #(
    .INIT(64'h4ff4444444444444)
  ) __227__ (
    .I5(G9),
    .I4(__6__),
    .I3(G7),
    .I2(__35__),
    .I1(__44__),
    .I0(__75__),
    .O(__76__)
  );
  LUT6 #(
    .INIT(64'h2000000000000003)
  ) __228__ (
    .I5(G10),
    .I4(G8),
    .I3(G7),
    .I2(G11),
    .I1(G5),
    .I0(G9),
    .O(__77__)
  );
  LUT3 #(
    .INIT(8'h40)
  ) __229__ (
    .I2(G1),
    .I1(G0),
    .I0(G4),
    .O(__78__)
  );
  LUT3 #(
    .INIT(8'h40)
  ) __230__ (
    .I2(G2),
    .I1(G4),
    .I0(G5),
    .O(__79__)
  );
  LUT3 #(
    .INIT(8'h04)
  ) __231__ (
    .I2(G12),
    .I1(__3__),
    .I0(__31__),
    .O(__80__)
  );
  LUT6 #(
    .INIT(64'h0000bfffbfffbfff)
  ) __232__ (
    .I5(__80__),
    .I4(__79__),
    .I3(__43__),
    .I2(G12),
    .I1(__78__),
    .I0(__37__),
    .O(__81__)
  );
  LUT5 #(
    .INIT(32'h0003000a)
  ) __233__ (
    .I4(G13),
    .I3(G12),
    .I2(__31__),
    .I1(__67__),
    .I0(__3__),
    .O(__82__)
  );
  LUT5 #(
    .INIT(32'ha3ff04f7)
  ) __234__ (
    .I4(G9),
    .I3(G10),
    .I2(G8),
    .I1(G11),
    .I0(G7),
    .O(__83__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __235__ (
    .I1(G8),
    .I0(__6__),
    .O(__84__)
  );
  LUT5 #(
    .INIT(32'h70000000)
  ) __236__ (
    .I4(G10),
    .I3(G7),
    .I2(__6__),
    .I1(G9),
    .I0(G8),
    .O(__85__)
  );
  LUT3 #(
    .INIT(8'h40)
  ) __237__ (
    .I2(G9),
    .I1(G7),
    .I0(G10),
    .O(__86__)
  );
  LUT6 #(
    .INIT(64'hfff5fcf0fcf0fcf0)
  ) __238__ (
    .I5(G6),
    .I4(__44__),
    .I3(__86__),
    .I2(__85__),
    .I1(__84__),
    .I0(__83__),
    .O(__87__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __239__ (
    .I1(G10),
    .I0(G7),
    .O(__88__)
  );
  LUT6 #(
    .INIT(64'h00af030f33ff33ff)
  ) __240__ (
    .I5(__44__),
    .I4(G6),
    .I3(__86__),
    .I2(__88__),
    .I1(__84__),
    .I0(G9),
    .O(__89__)
  );
  LUT6 #(
    .INIT(64'ha2aa22aaaaaaaaaa)
  ) __241__ (
    .I5(G10),
    .I4(G9),
    .I3(G8),
    .I2(G7),
    .I1(__6__),
    .I0(__89__),
    .O(__90__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __242__ (
    .I1(G7),
    .I0(G11),
    .O(__91__)
  );
  LUT5 #(
    .INIT(32'h5f5f1f5f)
  ) __243__ (
    .I4(G10),
    .I3(G9),
    .I2(G8),
    .I1(G11),
    .I0(__10__),
    .O(__92__)
  );
  LUT6 #(
    .INIT(64'h07000f0fff00ffff)
  ) __244__ (
    .I5(G8),
    .I4(G6),
    .I3(__92__),
    .I2(__40__),
    .I1(G9),
    .I0(__91__),
    .O(__93__)
  );
  LUT6 #(
    .INIT(64'hf55557df5fff5f5f)
  ) __245__ (
    .I5(G1),
    .I4(G4),
    .I3(G5),
    .I2(G2),
    .I1(G3),
    .I0(G6),
    .O(__94__)
  );
  LUT4 #(
    .INIT(16'h0004)
  ) __246__ (
    .I3(G12),
    .I2(G13),
    .I1(__3__),
    .I0(__31__),
    .O(__95__)
  );
  LUT6 #(
    .INIT(64'h79c8000000000000)
  ) __247__ (
    .I5(G6),
    .I4(__95__),
    .I3(G3),
    .I2(G5),
    .I1(G2),
    .I0(G4),
    .O(__96__)
  );
  LUT6 #(
    .INIT(64'hffffffff40ff4040)
  ) __248__ (
    .I5(__96__),
    .I4(__44__),
    .I3(__1__),
    .I2(__69__),
    .I1(__68__),
    .I0(__94__),
    .O(__97__)
  );
  LUT6 #(
    .INIT(64'hd55555ff5ff777ff)
  ) __249__ (
    .I5(G5),
    .I4(G2),
    .I3(G1),
    .I2(G4),
    .I1(G6),
    .I0(G3),
    .O(__98__)
  );
  LUT5 #(
    .INIT(32'h10000000)
  ) __250__ (
    .I4(G6),
    .I3(G3),
    .I2(G4),
    .I1(__19__),
    .I0(G5),
    .O(__99__)
  );
  LUT5 #(
    .INIT(32'h0000e000)
  ) __251__ (
    .I4(G5),
    .I3(G2),
    .I2(G13),
    .I1(__54__),
    .I0(__50__),
    .O(__100__)
  );
  LUT5 #(
    .INIT(32'h5559ffff)
  ) __252__ (
    .I4(G6),
    .I3(G10),
    .I2(G9),
    .I1(G7),
    .I0(G5),
    .O(__101__)
  );
  LUT5 #(
    .INIT(32'h00f40000)
  ) __253__ (
    .I4(G8),
    .I3(__101__),
    .I2(__33__),
    .I1(G13),
    .I0(__55__),
    .O(__102__)
  );
  LUT6 #(
    .INIT(64'ha000a800a000a000)
  ) __254__ (
    .I5(G6),
    .I4(G9),
    .I3(G8),
    .I2(G0),
    .I1(__4__),
    .I0(__65__),
    .O(__103__)
  );
  LUT6 #(
    .INIT(64'h7ffffffffffffffc)
  ) __255__ (
    .I5(G6),
    .I4(G10),
    .I3(G4),
    .I2(G5),
    .I1(G11),
    .I0(G9),
    .O(__104__)
  );
  LUT6 #(
    .INIT(64'h0300030003005555)
  ) __256__ (
    .I5(G8),
    .I4(G7),
    .I3(G4),
    .I2(G5),
    .I1(__47__),
    .I0(__104__),
    .O(__105__)
  );
  LUT4 #(
    .INIT(16'h0e00)
  ) __257__ (
    .I3(__33__),
    .I2(G12),
    .I1(__105__),
    .I0(__99__),
    .O(__106__)
  );
  LUT6 #(
    .INIT(64'hffffffffffff0f08)
  ) __258__ (
    .I5(__106__),
    .I4(__103__),
    .I3(__102__),
    .I2(G12),
    .I1(__100__),
    .I0(__99__),
    .O(__107__)
  );
  LUT6 #(
    .INIT(64'h3fd8c0f000000000)
  ) __259__ (
    .I5(G5),
    .I4(G0),
    .I3(G3),
    .I2(G1),
    .I1(G4),
    .I0(G2),
    .O(__108__)
  );
  LUT4 #(
    .INIT(16'h7173)
  ) __260__ (
    .I3(G3),
    .I2(G5),
    .I1(G4),
    .I0(G6),
    .O(__109__)
  );
  LUT6 #(
    .INIT(64'h40c04000c0c04000)
  ) __261__ (
    .I5(G2),
    .I4(G4),
    .I3(G1),
    .I2(__69__),
    .I1(__68__),
    .I0(__109__),
    .O(__110__)
  );
  LUT6 #(
    .INIT(64'hffffffffff808080)
  ) __262__ (
    .I5(__110__),
    .I4(__44__),
    .I3(__108__),
    .I2(G4),
    .I1(__95__),
    .I0(__2__),
    .O(__111__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __263__ (
    .I1(G4),
    .I0(G1),
    .O(__112__)
  );
  LUT6 #(
    .INIT(64'h0000000000002080)
  ) __264__ (
    .I5(__31__),
    .I4(__67__),
    .I3(G5),
    .I2(G2),
    .I1(__112__),
    .I0(__69__),
    .O(__113__)
  );
  LUT3 #(
    .INIT(8'h04)
  ) __265__ (
    .I2(G13),
    .I1(G3),
    .I0(__7__),
    .O(__114__)
  );
  LUT6 #(
    .INIT(64'h0000000000008fff)
  ) __266__ (
    .I5(__114__),
    .I4(__113__),
    .I3(__28__),
    .I2(__95__),
    .I1(G2),
    .I0(G4),
    .O(__115__)
  );
  LUT6 #(
    .INIT(64'h0fff88ff00ff00ff)
  ) __267__ (
    .I5(__44__),
    .I4(G0),
    .I3(__115__),
    .I2(__12__),
    .I1(G3),
    .I0(__112__),
    .O(__116__)
  );
  LUT6 #(
    .INIT(64'h5cfbaa0800000000)
  ) __268__ (
    .I5(G0),
    .I4(G4),
    .I3(G3),
    .I2(G2),
    .I1(G5),
    .I0(G1),
    .O(__117__)
  );
  LUT6 #(
    .INIT(64'ha000a30000000000)
  ) __269__ (
    .I5(G6),
    .I4(__19__),
    .I3(G3),
    .I2(G4),
    .I1(G5),
    .I0(__25__),
    .O(__118__)
  );
  LUT4 #(
    .INIT(16'hf400)
  ) __270__ (
    .I3(__118__),
    .I2(__33__),
    .I1(G13),
    .I0(__55__),
    .O(__119__)
  );
  LUT5 #(
    .INIT(32'h80000f0f)
  ) __271__ (
    .I4(G6),
    .I3(G8),
    .I2(G4),
    .I1(G5),
    .I0(G11),
    .O(__120__)
  );
  LUT6 #(
    .INIT(64'hbf00bfbfbfbfbfbf)
  ) __272__ (
    .I5(G13),
    .I4(__68__),
    .I3(__15__),
    .I2(__33__),
    .I1(__120__),
    .I0(G2),
    .O(__121__)
  );
  LUT6 #(
    .INIT(64'hc800880000000000)
  ) __273__ (
    .I5(G6),
    .I4(G3),
    .I3(G4),
    .I2(__33__),
    .I1(__52__),
    .I0(__100__),
    .O(__122__)
  );
  LUT6 #(
    .INIT(64'h88888888fffff8ff)
  ) __274__ (
    .I5(G12),
    .I4(__122__),
    .I3(__121__),
    .I2(__119__),
    .I1(__44__),
    .I0(__117__),
    .O(__123__)
  );
  LUT4 #(
    .INIT(16'h7f30)
  ) __275__ (
    .I3(G10),
    .I2(G11),
    .I1(G7),
    .I0(G9),
    .O(__124__)
  );
  LUT5 #(
    .INIT(32'h7af0fa08)
  ) __276__ (
    .I4(G4),
    .I3(G5),
    .I2(G2),
    .I1(G6),
    .I0(G3),
    .O(__125__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __277__ (
    .I1(G8),
    .I0(G7),
    .O(__126__)
  );
  LUT6 #(
    .INIT(64'h7ffffffffffffffc)
  ) __278__ (
    .I5(G6),
    .I4(G10),
    .I3(G9),
    .I2(G5),
    .I1(G11),
    .I0(G4),
    .O(__127__)
  );
  LUT6 #(
    .INIT(64'hdddddddddddddd0d)
  ) __279__ (
    .I5(G6),
    .I4(G4),
    .I3(G5),
    .I2(__29__),
    .I1(__127__),
    .I0(__126__),
    .O(__128__)
  );
  LUT3 #(
    .INIT(8'h78)
  ) __280__ (
    .I2(G2),
    .I1(G3),
    .I0(G5),
    .O(__129__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __281__ (
    .I1(G3),
    .I0(G0),
    .O(__130__)
  );
  LUT6 #(
    .INIT(64'h0000000070000000)
  ) __282__ (
    .I5(G13),
    .I4(G2),
    .I3(G5),
    .I2(__80__),
    .I1(G3),
    .I0(G4),
    .O(__131__)
  );
  LUT6 #(
    .INIT(64'h00000000dfab0000)
  ) __283__ (
    .I5(G12),
    .I4(G13),
    .I3(G2),
    .I2(G4),
    .I1(G6),
    .I0(G5),
    .O(__132__)
  );
  LUT4 #(
    .INIT(16'h1000)
  ) __284__ (
    .I3(G1),
    .I2(__132__),
    .I1(__31__),
    .I0(__67__),
    .O(__133__)
  );
  LUT6 #(
    .INIT(64'hffffffffffffff40)
  ) __285__ (
    .I5(__114__),
    .I4(__133__),
    .I3(__131__),
    .I2(__44__),
    .I1(__112__),
    .I0(__130__),
    .O(__134__)
  );
  LUT6 #(
    .INIT(64'h00000000000000f4)
  ) __286__ (
    .I5(__19__),
    .I4(G4),
    .I3(G5),
    .I2(__33__),
    .I1(G13),
    .I0(__55__),
    .O(__135__)
  );
  LUT4 #(
    .INIT(16'h1400)
  ) __287__ (
    .I3(G8),
    .I2(G9),
    .I1(G7),
    .I0(G10),
    .O(__136__)
  );
  LUT6 #(
    .INIT(64'h00000000e0000000)
  ) __288__ (
    .I5(G5),
    .I4(G2),
    .I3(G13),
    .I2(__136__),
    .I1(__54__),
    .I0(__50__),
    .O(__137__)
  );
  LUT6 #(
    .INIT(64'h0200000002000300)
  ) __289__ (
    .I5(__16__),
    .I4(G3),
    .I3(__33__),
    .I2(G2),
    .I1(G12),
    .I0(__136__),
    .O(__138__)
  );
  LUT4 #(
    .INIT(16'h8000)
  ) __290__ (
    .I3(G8),
    .I2(__4__),
    .I1(__8__),
    .I0(__65__),
    .O(__139__)
  );
  LUT6 #(
    .INIT(64'hffffffffffff0e00)
  ) __291__ (
    .I5(__139__),
    .I4(__138__),
    .I3(__53__),
    .I2(G12),
    .I1(__137__),
    .I0(__135__),
    .O(__140__)
  );
  LUT4 #(
    .INIT(16'h0100)
  ) __292__ (
    .I3(G7),
    .I2(G10),
    .I1(G4),
    .I0(G0),
    .O(__141__)
  );
  LUT6 #(
    .INIT(64'h79c8000000000000)
  ) __293__ (
    .I5(G11),
    .I4(__6__),
    .I3(G8),
    .I2(G10),
    .I1(G7),
    .I0(G9),
    .O(__142__)
  );
  LUT6 #(
    .INIT(64'hffffffff01000000)
  ) __294__ (
    .I5(__142__),
    .I4(__43__),
    .I3(G12),
    .I2(G13),
    .I1(__37__),
    .I0(__14__),
    .O(__143__)
  );
  LUT5 #(
    .INIT(32'hafbb3f0f)
  ) __295__ (
    .I4(G2),
    .I3(G4),
    .I2(G3),
    .I1(G5),
    .I0(G1),
    .O(__144__)
  );
  LUT6 #(
    .INIT(64'hf55557df5fff5f5f)
  ) __296__ (
    .I5(G6),
    .I4(G9),
    .I3(G10),
    .I2(G7),
    .I1(G8),
    .I0(G11),
    .O(__145__)
  );
  LUT6 #(
    .INIT(64'h000000005575775f)
  ) __297__ (
    .I5(G1),
    .I4(G3),
    .I3(G5),
    .I2(G4),
    .I1(G2),
    .I0(G0),
    .O(__146__)
  );
  LUT6 #(
    .INIT(64'h8003008a00000000)
  ) __298__ (
    .I5(G2),
    .I4(G3),
    .I3(G4),
    .I2(G5),
    .I1(G1),
    .I0(G0),
    .O(__147__)
  );
  LUT6 #(
    .INIT(64'h000000000000fef0)
  ) __299__ (
    .I5(__147__),
    .I4(__146__),
    .I3(G7),
    .I2(G6),
    .I1(G10),
    .I0(__11__),
    .O(__148__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __300__ (
    .I1(G6),
    .I0(G9),
    .O(__149__)
  );
  LUT5 #(
    .INIT(32'h10080002)
  ) __301__ (
    .I4(G6),
    .I3(G10),
    .I2(G9),
    .I1(G8),
    .I0(G7),
    .O(__150__)
  );
  assign G532 = __123__;
  assign G546 = __0__;
  assign G550 = __116__;
  assign G547 = __76__;
  assign G548 = __143__;
  assign G535 = __140__;
  assign G45 = __17__;
  assign G551 = __111__;
  assign G539 = __72__;
  assign G530 = __45__;
  assign G552 = __97__;
  assign G549 = __134__;
  assign G542 = __87__;
  assign G537 = __107__;
endmodule
