module alu_1024(
  input wire a0, input wire b0,
  input wire a1, input wire b1,
  input wire a2, input wire b2,
  input wire a3, input wire b3,
  input wire a4, input wire b4,
  input wire a5, input wire b5,
  input wire a6, input wire b6,
  input wire a7, input wire b7,
  input wire a8, input wire b8,
  input wire a9, input wire b9,
  input wire a10, input wire b10,
  input wire a11, input wire b11,
  input wire a12, input wire b12,
  input wire a13, input wire b13,
  input wire a14, input wire b14,
  input wire a15, input wire b15,
  input wire a16, input wire b16,
  input wire a17, input wire b17,
  input wire a18, input wire b18,
  input wire a19, input wire b19,
  input wire a20, input wire b20,
  input wire a21, input wire b21,
  input wire a22, input wire b22,
  input wire a23, input wire b23,
  input wire a24, input wire b24,
  input wire a25, input wire b25,
  input wire a26, input wire b26,
  input wire a27, input wire b27,
  input wire a28, input wire b28,
  input wire a29, input wire b29,
  input wire a30, input wire b30,
  input wire a31, input wire b31,
  input wire a32, input wire b32,
  input wire a33, input wire b33,
  input wire a34, input wire b34,
  input wire a35, input wire b35,
  input wire a36, input wire b36,
  input wire a37, input wire b37,
  input wire a38, input wire b38,
  input wire a39, input wire b39,
  input wire a40, input wire b40,
  input wire a41, input wire b41,
  input wire a42, input wire b42,
  input wire a43, input wire b43,
  input wire a44, input wire b44,
  input wire a45, input wire b45,
  input wire a46, input wire b46,
  input wire a47, input wire b47,
  input wire a48, input wire b48,
  input wire a49, input wire b49,
  input wire a50, input wire b50,
  input wire a51, input wire b51,
  input wire a52, input wire b52,
  input wire a53, input wire b53,
  input wire a54, input wire b54,
  input wire a55, input wire b55,
  input wire a56, input wire b56,
  input wire a57, input wire b57,
  input wire a58, input wire b58,
  input wire a59, input wire b59,
  input wire a60, input wire b60,
  input wire a61, input wire b61,
  input wire a62, input wire b62,
  input wire a63, input wire b63,
  input wire a64, input wire b64,
  input wire a65, input wire b65,
  input wire a66, input wire b66,
  input wire a67, input wire b67,
  input wire a68, input wire b68,
  input wire a69, input wire b69,
  input wire a70, input wire b70,
  input wire a71, input wire b71,
  input wire a72, input wire b72,
  input wire a73, input wire b73,
  input wire a74, input wire b74,
  input wire a75, input wire b75,
  input wire a76, input wire b76,
  input wire a77, input wire b77,
  input wire a78, input wire b78,
  input wire a79, input wire b79,
  input wire a80, input wire b80,
  input wire a81, input wire b81,
  input wire a82, input wire b82,
  input wire a83, input wire b83,
  input wire a84, input wire b84,
  input wire a85, input wire b85,
  input wire a86, input wire b86,
  input wire a87, input wire b87,
  input wire a88, input wire b88,
  input wire a89, input wire b89,
  input wire a90, input wire b90,
  input wire a91, input wire b91,
  input wire a92, input wire b92,
  input wire a93, input wire b93,
  input wire a94, input wire b94,
  input wire a95, input wire b95,
  input wire a96, input wire b96,
  input wire a97, input wire b97,
  input wire a98, input wire b98,
  input wire a99, input wire b99,
  input wire a100, input wire b100,
  input wire a101, input wire b101,
  input wire a102, input wire b102,
  input wire a103, input wire b103,
  input wire a104, input wire b104,
  input wire a105, input wire b105,
  input wire a106, input wire b106,
  input wire a107, input wire b107,
  input wire a108, input wire b108,
  input wire a109, input wire b109,
  input wire a110, input wire b110,
  input wire a111, input wire b111,
  input wire a112, input wire b112,
  input wire a113, input wire b113,
  input wire a114, input wire b114,
  input wire a115, input wire b115,
  input wire a116, input wire b116,
  input wire a117, input wire b117,
  input wire a118, input wire b118,
  input wire a119, input wire b119,
  input wire a120, input wire b120,
  input wire a121, input wire b121,
  input wire a122, input wire b122,
  input wire a123, input wire b123,
  input wire a124, input wire b124,
  input wire a125, input wire b125,
  input wire a126, input wire b126,
  input wire a127, input wire b127,
  input wire a128, input wire b128,
  input wire a129, input wire b129,
  input wire a130, input wire b130,
  input wire a131, input wire b131,
  input wire a132, input wire b132,
  input wire a133, input wire b133,
  input wire a134, input wire b134,
  input wire a135, input wire b135,
  input wire a136, input wire b136,
  input wire a137, input wire b137,
  input wire a138, input wire b138,
  input wire a139, input wire b139,
  input wire a140, input wire b140,
  input wire a141, input wire b141,
  input wire a142, input wire b142,
  input wire a143, input wire b143,
  input wire a144, input wire b144,
  input wire a145, input wire b145,
  input wire a146, input wire b146,
  input wire a147, input wire b147,
  input wire a148, input wire b148,
  input wire a149, input wire b149,
  input wire a150, input wire b150,
  input wire a151, input wire b151,
  input wire a152, input wire b152,
  input wire a153, input wire b153,
  input wire a154, input wire b154,
  input wire a155, input wire b155,
  input wire a156, input wire b156,
  input wire a157, input wire b157,
  input wire a158, input wire b158,
  input wire a159, input wire b159,
  input wire a160, input wire b160,
  input wire a161, input wire b161,
  input wire a162, input wire b162,
  input wire a163, input wire b163,
  input wire a164, input wire b164,
  input wire a165, input wire b165,
  input wire a166, input wire b166,
  input wire a167, input wire b167,
  input wire a168, input wire b168,
  input wire a169, input wire b169,
  input wire a170, input wire b170,
  input wire a171, input wire b171,
  input wire a172, input wire b172,
  input wire a173, input wire b173,
  input wire a174, input wire b174,
  input wire a175, input wire b175,
  input wire a176, input wire b176,
  input wire a177, input wire b177,
  input wire a178, input wire b178,
  input wire a179, input wire b179,
  input wire a180, input wire b180,
  input wire a181, input wire b181,
  input wire a182, input wire b182,
  input wire a183, input wire b183,
  input wire a184, input wire b184,
  input wire a185, input wire b185,
  input wire a186, input wire b186,
  input wire a187, input wire b187,
  input wire a188, input wire b188,
  input wire a189, input wire b189,
  input wire a190, input wire b190,
  input wire a191, input wire b191,
  input wire a192, input wire b192,
  input wire a193, input wire b193,
  input wire a194, input wire b194,
  input wire a195, input wire b195,
  input wire a196, input wire b196,
  input wire a197, input wire b197,
  input wire a198, input wire b198,
  input wire a199, input wire b199,
  input wire a200, input wire b200,
  input wire a201, input wire b201,
  input wire a202, input wire b202,
  input wire a203, input wire b203,
  input wire a204, input wire b204,
  input wire a205, input wire b205,
  input wire a206, input wire b206,
  input wire a207, input wire b207,
  input wire a208, input wire b208,
  input wire a209, input wire b209,
  input wire a210, input wire b210,
  input wire a211, input wire b211,
  input wire a212, input wire b212,
  input wire a213, input wire b213,
  input wire a214, input wire b214,
  input wire a215, input wire b215,
  input wire a216, input wire b216,
  input wire a217, input wire b217,
  input wire a218, input wire b218,
  input wire a219, input wire b219,
  input wire a220, input wire b220,
  input wire a221, input wire b221,
  input wire a222, input wire b222,
  input wire a223, input wire b223,
  input wire a224, input wire b224,
  input wire a225, input wire b225,
  input wire a226, input wire b226,
  input wire a227, input wire b227,
  input wire a228, input wire b228,
  input wire a229, input wire b229,
  input wire a230, input wire b230,
  input wire a231, input wire b231,
  input wire a232, input wire b232,
  input wire a233, input wire b233,
  input wire a234, input wire b234,
  input wire a235, input wire b235,
  input wire a236, input wire b236,
  input wire a237, input wire b237,
  input wire a238, input wire b238,
  input wire a239, input wire b239,
  input wire a240, input wire b240,
  input wire a241, input wire b241,
  input wire a242, input wire b242,
  input wire a243, input wire b243,
  input wire a244, input wire b244,
  input wire a245, input wire b245,
  input wire a246, input wire b246,
  input wire a247, input wire b247,
  input wire a248, input wire b248,
  input wire a249, input wire b249,
  input wire a250, input wire b250,
  input wire a251, input wire b251,
  input wire a252, input wire b252,
  input wire a253, input wire b253,
  input wire a254, input wire b254,
  input wire a255, input wire b255,
  input wire a256, input wire b256,
  input wire a257, input wire b257,
  input wire a258, input wire b258,
  input wire a259, input wire b259,
  input wire a260, input wire b260,
  input wire a261, input wire b261,
  input wire a262, input wire b262,
  input wire a263, input wire b263,
  input wire a264, input wire b264,
  input wire a265, input wire b265,
  input wire a266, input wire b266,
  input wire a267, input wire b267,
  input wire a268, input wire b268,
  input wire a269, input wire b269,
  input wire a270, input wire b270,
  input wire a271, input wire b271,
  input wire a272, input wire b272,
  input wire a273, input wire b273,
  input wire a274, input wire b274,
  input wire a275, input wire b275,
  input wire a276, input wire b276,
  input wire a277, input wire b277,
  input wire a278, input wire b278,
  input wire a279, input wire b279,
  input wire a280, input wire b280,
  input wire a281, input wire b281,
  input wire a282, input wire b282,
  input wire a283, input wire b283,
  input wire a284, input wire b284,
  input wire a285, input wire b285,
  input wire a286, input wire b286,
  input wire a287, input wire b287,
  input wire a288, input wire b288,
  input wire a289, input wire b289,
  input wire a290, input wire b290,
  input wire a291, input wire b291,
  input wire a292, input wire b292,
  input wire a293, input wire b293,
  input wire a294, input wire b294,
  input wire a295, input wire b295,
  input wire a296, input wire b296,
  input wire a297, input wire b297,
  input wire a298, input wire b298,
  input wire a299, input wire b299,
  input wire a300, input wire b300,
  input wire a301, input wire b301,
  input wire a302, input wire b302,
  input wire a303, input wire b303,
  input wire a304, input wire b304,
  input wire a305, input wire b305,
  input wire a306, input wire b306,
  input wire a307, input wire b307,
  input wire a308, input wire b308,
  input wire a309, input wire b309,
  input wire a310, input wire b310,
  input wire a311, input wire b311,
  input wire a312, input wire b312,
  input wire a313, input wire b313,
  input wire a314, input wire b314,
  input wire a315, input wire b315,
  input wire a316, input wire b316,
  input wire a317, input wire b317,
  input wire a318, input wire b318,
  input wire a319, input wire b319,
  input wire a320, input wire b320,
  input wire a321, input wire b321,
  input wire a322, input wire b322,
  input wire a323, input wire b323,
  input wire a324, input wire b324,
  input wire a325, input wire b325,
  input wire a326, input wire b326,
  input wire a327, input wire b327,
  input wire a328, input wire b328,
  input wire a329, input wire b329,
  input wire a330, input wire b330,
  input wire a331, input wire b331,
  input wire a332, input wire b332,
  input wire a333, input wire b333,
  input wire a334, input wire b334,
  input wire a335, input wire b335,
  input wire a336, input wire b336,
  input wire a337, input wire b337,
  input wire a338, input wire b338,
  input wire a339, input wire b339,
  input wire a340, input wire b340,
  input wire a341, input wire b341,
  input wire a342, input wire b342,
  input wire a343, input wire b343,
  input wire a344, input wire b344,
  input wire a345, input wire b345,
  input wire a346, input wire b346,
  input wire a347, input wire b347,
  input wire a348, input wire b348,
  input wire a349, input wire b349,
  input wire a350, input wire b350,
  input wire a351, input wire b351,
  input wire a352, input wire b352,
  input wire a353, input wire b353,
  input wire a354, input wire b354,
  input wire a355, input wire b355,
  input wire a356, input wire b356,
  input wire a357, input wire b357,
  input wire a358, input wire b358,
  input wire a359, input wire b359,
  input wire a360, input wire b360,
  input wire a361, input wire b361,
  input wire a362, input wire b362,
  input wire a363, input wire b363,
  input wire a364, input wire b364,
  input wire a365, input wire b365,
  input wire a366, input wire b366,
  input wire a367, input wire b367,
  input wire a368, input wire b368,
  input wire a369, input wire b369,
  input wire a370, input wire b370,
  input wire a371, input wire b371,
  input wire a372, input wire b372,
  input wire a373, input wire b373,
  input wire a374, input wire b374,
  input wire a375, input wire b375,
  input wire a376, input wire b376,
  input wire a377, input wire b377,
  input wire a378, input wire b378,
  input wire a379, input wire b379,
  input wire a380, input wire b380,
  input wire a381, input wire b381,
  input wire a382, input wire b382,
  input wire a383, input wire b383,
  input wire a384, input wire b384,
  input wire a385, input wire b385,
  input wire a386, input wire b386,
  input wire a387, input wire b387,
  input wire a388, input wire b388,
  input wire a389, input wire b389,
  input wire a390, input wire b390,
  input wire a391, input wire b391,
  input wire a392, input wire b392,
  input wire a393, input wire b393,
  input wire a394, input wire b394,
  input wire a395, input wire b395,
  input wire a396, input wire b396,
  input wire a397, input wire b397,
  input wire a398, input wire b398,
  input wire a399, input wire b399,
  input wire a400, input wire b400,
  input wire a401, input wire b401,
  input wire a402, input wire b402,
  input wire a403, input wire b403,
  input wire a404, input wire b404,
  input wire a405, input wire b405,
  input wire a406, input wire b406,
  input wire a407, input wire b407,
  input wire a408, input wire b408,
  input wire a409, input wire b409,
  input wire a410, input wire b410,
  input wire a411, input wire b411,
  input wire a412, input wire b412,
  input wire a413, input wire b413,
  input wire a414, input wire b414,
  input wire a415, input wire b415,
  input wire a416, input wire b416,
  input wire a417, input wire b417,
  input wire a418, input wire b418,
  input wire a419, input wire b419,
  input wire a420, input wire b420,
  input wire a421, input wire b421,
  input wire a422, input wire b422,
  input wire a423, input wire b423,
  input wire a424, input wire b424,
  input wire a425, input wire b425,
  input wire a426, input wire b426,
  input wire a427, input wire b427,
  input wire a428, input wire b428,
  input wire a429, input wire b429,
  input wire a430, input wire b430,
  input wire a431, input wire b431,
  input wire a432, input wire b432,
  input wire a433, input wire b433,
  input wire a434, input wire b434,
  input wire a435, input wire b435,
  input wire a436, input wire b436,
  input wire a437, input wire b437,
  input wire a438, input wire b438,
  input wire a439, input wire b439,
  input wire a440, input wire b440,
  input wire a441, input wire b441,
  input wire a442, input wire b442,
  input wire a443, input wire b443,
  input wire a444, input wire b444,
  input wire a445, input wire b445,
  input wire a446, input wire b446,
  input wire a447, input wire b447,
  input wire a448, input wire b448,
  input wire a449, input wire b449,
  input wire a450, input wire b450,
  input wire a451, input wire b451,
  input wire a452, input wire b452,
  input wire a453, input wire b453,
  input wire a454, input wire b454,
  input wire a455, input wire b455,
  input wire a456, input wire b456,
  input wire a457, input wire b457,
  input wire a458, input wire b458,
  input wire a459, input wire b459,
  input wire a460, input wire b460,
  input wire a461, input wire b461,
  input wire a462, input wire b462,
  input wire a463, input wire b463,
  input wire a464, input wire b464,
  input wire a465, input wire b465,
  input wire a466, input wire b466,
  input wire a467, input wire b467,
  input wire a468, input wire b468,
  input wire a469, input wire b469,
  input wire a470, input wire b470,
  input wire a471, input wire b471,
  input wire a472, input wire b472,
  input wire a473, input wire b473,
  input wire a474, input wire b474,
  input wire a475, input wire b475,
  input wire a476, input wire b476,
  input wire a477, input wire b477,
  input wire a478, input wire b478,
  input wire a479, input wire b479,
  input wire a480, input wire b480,
  input wire a481, input wire b481,
  input wire a482, input wire b482,
  input wire a483, input wire b483,
  input wire a484, input wire b484,
  input wire a485, input wire b485,
  input wire a486, input wire b486,
  input wire a487, input wire b487,
  input wire a488, input wire b488,
  input wire a489, input wire b489,
  input wire a490, input wire b490,
  input wire a491, input wire b491,
  input wire a492, input wire b492,
  input wire a493, input wire b493,
  input wire a494, input wire b494,
  input wire a495, input wire b495,
  input wire a496, input wire b496,
  input wire a497, input wire b497,
  input wire a498, input wire b498,
  input wire a499, input wire b499,
  input wire a500, input wire b500,
  input wire a501, input wire b501,
  input wire a502, input wire b502,
  input wire a503, input wire b503,
  input wire a504, input wire b504,
  input wire a505, input wire b505,
  input wire a506, input wire b506,
  input wire a507, input wire b507,
  input wire a508, input wire b508,
  input wire a509, input wire b509,
  input wire a510, input wire b510,
  input wire a511, input wire b511,
  input wire a512, input wire b512,
  input wire a513, input wire b513,
  input wire a514, input wire b514,
  input wire a515, input wire b515,
  input wire a516, input wire b516,
  input wire a517, input wire b517,
  input wire a518, input wire b518,
  input wire a519, input wire b519,
  input wire a520, input wire b520,
  input wire a521, input wire b521,
  input wire a522, input wire b522,
  input wire a523, input wire b523,
  input wire a524, input wire b524,
  input wire a525, input wire b525,
  input wire a526, input wire b526,
  input wire a527, input wire b527,
  input wire a528, input wire b528,
  input wire a529, input wire b529,
  input wire a530, input wire b530,
  input wire a531, input wire b531,
  input wire a532, input wire b532,
  input wire a533, input wire b533,
  input wire a534, input wire b534,
  input wire a535, input wire b535,
  input wire a536, input wire b536,
  input wire a537, input wire b537,
  input wire a538, input wire b538,
  input wire a539, input wire b539,
  input wire a540, input wire b540,
  input wire a541, input wire b541,
  input wire a542, input wire b542,
  input wire a543, input wire b543,
  input wire a544, input wire b544,
  input wire a545, input wire b545,
  input wire a546, input wire b546,
  input wire a547, input wire b547,
  input wire a548, input wire b548,
  input wire a549, input wire b549,
  input wire a550, input wire b550,
  input wire a551, input wire b551,
  input wire a552, input wire b552,
  input wire a553, input wire b553,
  input wire a554, input wire b554,
  input wire a555, input wire b555,
  input wire a556, input wire b556,
  input wire a557, input wire b557,
  input wire a558, input wire b558,
  input wire a559, input wire b559,
  input wire a560, input wire b560,
  input wire a561, input wire b561,
  input wire a562, input wire b562,
  input wire a563, input wire b563,
  input wire a564, input wire b564,
  input wire a565, input wire b565,
  input wire a566, input wire b566,
  input wire a567, input wire b567,
  input wire a568, input wire b568,
  input wire a569, input wire b569,
  input wire a570, input wire b570,
  input wire a571, input wire b571,
  input wire a572, input wire b572,
  input wire a573, input wire b573,
  input wire a574, input wire b574,
  input wire a575, input wire b575,
  input wire a576, input wire b576,
  input wire a577, input wire b577,
  input wire a578, input wire b578,
  input wire a579, input wire b579,
  input wire a580, input wire b580,
  input wire a581, input wire b581,
  input wire a582, input wire b582,
  input wire a583, input wire b583,
  input wire a584, input wire b584,
  input wire a585, input wire b585,
  input wire a586, input wire b586,
  input wire a587, input wire b587,
  input wire a588, input wire b588,
  input wire a589, input wire b589,
  input wire a590, input wire b590,
  input wire a591, input wire b591,
  input wire a592, input wire b592,
  input wire a593, input wire b593,
  input wire a594, input wire b594,
  input wire a595, input wire b595,
  input wire a596, input wire b596,
  input wire a597, input wire b597,
  input wire a598, input wire b598,
  input wire a599, input wire b599,
  input wire a600, input wire b600,
  input wire a601, input wire b601,
  input wire a602, input wire b602,
  input wire a603, input wire b603,
  input wire a604, input wire b604,
  input wire a605, input wire b605,
  input wire a606, input wire b606,
  input wire a607, input wire b607,
  input wire a608, input wire b608,
  input wire a609, input wire b609,
  input wire a610, input wire b610,
  input wire a611, input wire b611,
  input wire a612, input wire b612,
  input wire a613, input wire b613,
  input wire a614, input wire b614,
  input wire a615, input wire b615,
  input wire a616, input wire b616,
  input wire a617, input wire b617,
  input wire a618, input wire b618,
  input wire a619, input wire b619,
  input wire a620, input wire b620,
  input wire a621, input wire b621,
  input wire a622, input wire b622,
  input wire a623, input wire b623,
  input wire a624, input wire b624,
  input wire a625, input wire b625,
  input wire a626, input wire b626,
  input wire a627, input wire b627,
  input wire a628, input wire b628,
  input wire a629, input wire b629,
  input wire a630, input wire b630,
  input wire a631, input wire b631,
  input wire a632, input wire b632,
  input wire a633, input wire b633,
  input wire a634, input wire b634,
  input wire a635, input wire b635,
  input wire a636, input wire b636,
  input wire a637, input wire b637,
  input wire a638, input wire b638,
  input wire a639, input wire b639,
  input wire a640, input wire b640,
  input wire a641, input wire b641,
  input wire a642, input wire b642,
  input wire a643, input wire b643,
  input wire a644, input wire b644,
  input wire a645, input wire b645,
  input wire a646, input wire b646,
  input wire a647, input wire b647,
  input wire a648, input wire b648,
  input wire a649, input wire b649,
  input wire a650, input wire b650,
  input wire a651, input wire b651,
  input wire a652, input wire b652,
  input wire a653, input wire b653,
  input wire a654, input wire b654,
  input wire a655, input wire b655,
  input wire a656, input wire b656,
  input wire a657, input wire b657,
  input wire a658, input wire b658,
  input wire a659, input wire b659,
  input wire a660, input wire b660,
  input wire a661, input wire b661,
  input wire a662, input wire b662,
  input wire a663, input wire b663,
  input wire a664, input wire b664,
  input wire a665, input wire b665,
  input wire a666, input wire b666,
  input wire a667, input wire b667,
  input wire a668, input wire b668,
  input wire a669, input wire b669,
  input wire a670, input wire b670,
  input wire a671, input wire b671,
  input wire a672, input wire b672,
  input wire a673, input wire b673,
  input wire a674, input wire b674,
  input wire a675, input wire b675,
  input wire a676, input wire b676,
  input wire a677, input wire b677,
  input wire a678, input wire b678,
  input wire a679, input wire b679,
  input wire a680, input wire b680,
  input wire a681, input wire b681,
  input wire a682, input wire b682,
  input wire a683, input wire b683,
  input wire a684, input wire b684,
  input wire a685, input wire b685,
  input wire a686, input wire b686,
  input wire a687, input wire b687,
  input wire a688, input wire b688,
  input wire a689, input wire b689,
  input wire a690, input wire b690,
  input wire a691, input wire b691,
  input wire a692, input wire b692,
  input wire a693, input wire b693,
  input wire a694, input wire b694,
  input wire a695, input wire b695,
  input wire a696, input wire b696,
  input wire a697, input wire b697,
  input wire a698, input wire b698,
  input wire a699, input wire b699,
  input wire a700, input wire b700,
  input wire a701, input wire b701,
  input wire a702, input wire b702,
  input wire a703, input wire b703,
  input wire a704, input wire b704,
  input wire a705, input wire b705,
  input wire a706, input wire b706,
  input wire a707, input wire b707,
  input wire a708, input wire b708,
  input wire a709, input wire b709,
  input wire a710, input wire b710,
  input wire a711, input wire b711,
  input wire a712, input wire b712,
  input wire a713, input wire b713,
  input wire a714, input wire b714,
  input wire a715, input wire b715,
  input wire a716, input wire b716,
  input wire a717, input wire b717,
  input wire a718, input wire b718,
  input wire a719, input wire b719,
  input wire a720, input wire b720,
  input wire a721, input wire b721,
  input wire a722, input wire b722,
  input wire a723, input wire b723,
  input wire a724, input wire b724,
  input wire a725, input wire b725,
  input wire a726, input wire b726,
  input wire a727, input wire b727,
  input wire a728, input wire b728,
  input wire a729, input wire b729,
  input wire a730, input wire b730,
  input wire a731, input wire b731,
  input wire a732, input wire b732,
  input wire a733, input wire b733,
  input wire a734, input wire b734,
  input wire a735, input wire b735,
  input wire a736, input wire b736,
  input wire a737, input wire b737,
  input wire a738, input wire b738,
  input wire a739, input wire b739,
  input wire a740, input wire b740,
  input wire a741, input wire b741,
  input wire a742, input wire b742,
  input wire a743, input wire b743,
  input wire a744, input wire b744,
  input wire a745, input wire b745,
  input wire a746, input wire b746,
  input wire a747, input wire b747,
  input wire a748, input wire b748,
  input wire a749, input wire b749,
  input wire a750, input wire b750,
  input wire a751, input wire b751,
  input wire a752, input wire b752,
  input wire a753, input wire b753,
  input wire a754, input wire b754,
  input wire a755, input wire b755,
  input wire a756, input wire b756,
  input wire a757, input wire b757,
  input wire a758, input wire b758,
  input wire a759, input wire b759,
  input wire a760, input wire b760,
  input wire a761, input wire b761,
  input wire a762, input wire b762,
  input wire a763, input wire b763,
  input wire a764, input wire b764,
  input wire a765, input wire b765,
  input wire a766, input wire b766,
  input wire a767, input wire b767,
  input wire a768, input wire b768,
  input wire a769, input wire b769,
  input wire a770, input wire b770,
  input wire a771, input wire b771,
  input wire a772, input wire b772,
  input wire a773, input wire b773,
  input wire a774, input wire b774,
  input wire a775, input wire b775,
  input wire a776, input wire b776,
  input wire a777, input wire b777,
  input wire a778, input wire b778,
  input wire a779, input wire b779,
  input wire a780, input wire b780,
  input wire a781, input wire b781,
  input wire a782, input wire b782,
  input wire a783, input wire b783,
  input wire a784, input wire b784,
  input wire a785, input wire b785,
  input wire a786, input wire b786,
  input wire a787, input wire b787,
  input wire a788, input wire b788,
  input wire a789, input wire b789,
  input wire a790, input wire b790,
  input wire a791, input wire b791,
  input wire a792, input wire b792,
  input wire a793, input wire b793,
  input wire a794, input wire b794,
  input wire a795, input wire b795,
  input wire a796, input wire b796,
  input wire a797, input wire b797,
  input wire a798, input wire b798,
  input wire a799, input wire b799,
  input wire a800, input wire b800,
  input wire a801, input wire b801,
  input wire a802, input wire b802,
  input wire a803, input wire b803,
  input wire a804, input wire b804,
  input wire a805, input wire b805,
  input wire a806, input wire b806,
  input wire a807, input wire b807,
  input wire a808, input wire b808,
  input wire a809, input wire b809,
  input wire a810, input wire b810,
  input wire a811, input wire b811,
  input wire a812, input wire b812,
  input wire a813, input wire b813,
  input wire a814, input wire b814,
  input wire a815, input wire b815,
  input wire a816, input wire b816,
  input wire a817, input wire b817,
  input wire a818, input wire b818,
  input wire a819, input wire b819,
  input wire a820, input wire b820,
  input wire a821, input wire b821,
  input wire a822, input wire b822,
  input wire a823, input wire b823,
  input wire a824, input wire b824,
  input wire a825, input wire b825,
  input wire a826, input wire b826,
  input wire a827, input wire b827,
  input wire a828, input wire b828,
  input wire a829, input wire b829,
  input wire a830, input wire b830,
  input wire a831, input wire b831,
  input wire a832, input wire b832,
  input wire a833, input wire b833,
  input wire a834, input wire b834,
  input wire a835, input wire b835,
  input wire a836, input wire b836,
  input wire a837, input wire b837,
  input wire a838, input wire b838,
  input wire a839, input wire b839,
  input wire a840, input wire b840,
  input wire a841, input wire b841,
  input wire a842, input wire b842,
  input wire a843, input wire b843,
  input wire a844, input wire b844,
  input wire a845, input wire b845,
  input wire a846, input wire b846,
  input wire a847, input wire b847,
  input wire a848, input wire b848,
  input wire a849, input wire b849,
  input wire a850, input wire b850,
  input wire a851, input wire b851,
  input wire a852, input wire b852,
  input wire a853, input wire b853,
  input wire a854, input wire b854,
  input wire a855, input wire b855,
  input wire a856, input wire b856,
  input wire a857, input wire b857,
  input wire a858, input wire b858,
  input wire a859, input wire b859,
  input wire a860, input wire b860,
  input wire a861, input wire b861,
  input wire a862, input wire b862,
  input wire a863, input wire b863,
  input wire a864, input wire b864,
  input wire a865, input wire b865,
  input wire a866, input wire b866,
  input wire a867, input wire b867,
  input wire a868, input wire b868,
  input wire a869, input wire b869,
  input wire a870, input wire b870,
  input wire a871, input wire b871,
  input wire a872, input wire b872,
  input wire a873, input wire b873,
  input wire a874, input wire b874,
  input wire a875, input wire b875,
  input wire a876, input wire b876,
  input wire a877, input wire b877,
  input wire a878, input wire b878,
  input wire a879, input wire b879,
  input wire a880, input wire b880,
  input wire a881, input wire b881,
  input wire a882, input wire b882,
  input wire a883, input wire b883,
  input wire a884, input wire b884,
  input wire a885, input wire b885,
  input wire a886, input wire b886,
  input wire a887, input wire b887,
  input wire a888, input wire b888,
  input wire a889, input wire b889,
  input wire a890, input wire b890,
  input wire a891, input wire b891,
  input wire a892, input wire b892,
  input wire a893, input wire b893,
  input wire a894, input wire b894,
  input wire a895, input wire b895,
  input wire a896, input wire b896,
  input wire a897, input wire b897,
  input wire a898, input wire b898,
  input wire a899, input wire b899,
  input wire a900, input wire b900,
  input wire a901, input wire b901,
  input wire a902, input wire b902,
  input wire a903, input wire b903,
  input wire a904, input wire b904,
  input wire a905, input wire b905,
  input wire a906, input wire b906,
  input wire a907, input wire b907,
  input wire a908, input wire b908,
  input wire a909, input wire b909,
  input wire a910, input wire b910,
  input wire a911, input wire b911,
  input wire a912, input wire b912,
  input wire a913, input wire b913,
  input wire a914, input wire b914,
  input wire a915, input wire b915,
  input wire a916, input wire b916,
  input wire a917, input wire b917,
  input wire a918, input wire b918,
  input wire a919, input wire b919,
  input wire a920, input wire b920,
  input wire a921, input wire b921,
  input wire a922, input wire b922,
  input wire a923, input wire b923,
  input wire a924, input wire b924,
  input wire a925, input wire b925,
  input wire a926, input wire b926,
  input wire a927, input wire b927,
  input wire a928, input wire b928,
  input wire a929, input wire b929,
  input wire a930, input wire b930,
  input wire a931, input wire b931,
  input wire a932, input wire b932,
  input wire a933, input wire b933,
  input wire a934, input wire b934,
  input wire a935, input wire b935,
  input wire a936, input wire b936,
  input wire a937, input wire b937,
  input wire a938, input wire b938,
  input wire a939, input wire b939,
  input wire a940, input wire b940,
  input wire a941, input wire b941,
  input wire a942, input wire b942,
  input wire a943, input wire b943,
  input wire a944, input wire b944,
  input wire a945, input wire b945,
  input wire a946, input wire b946,
  input wire a947, input wire b947,
  input wire a948, input wire b948,
  input wire a949, input wire b949,
  input wire a950, input wire b950,
  input wire a951, input wire b951,
  input wire a952, input wire b952,
  input wire a953, input wire b953,
  input wire a954, input wire b954,
  input wire a955, input wire b955,
  input wire a956, input wire b956,
  input wire a957, input wire b957,
  input wire a958, input wire b958,
  input wire a959, input wire b959,
  input wire a960, input wire b960,
  input wire a961, input wire b961,
  input wire a962, input wire b962,
  input wire a963, input wire b963,
  input wire a964, input wire b964,
  input wire a965, input wire b965,
  input wire a966, input wire b966,
  input wire a967, input wire b967,
  input wire a968, input wire b968,
  input wire a969, input wire b969,
  input wire a970, input wire b970,
  input wire a971, input wire b971,
  input wire a972, input wire b972,
  input wire a973, input wire b973,
  input wire a974, input wire b974,
  input wire a975, input wire b975,
  input wire a976, input wire b976,
  input wire a977, input wire b977,
  input wire a978, input wire b978,
  input wire a979, input wire b979,
  input wire a980, input wire b980,
  input wire a981, input wire b981,
  input wire a982, input wire b982,
  input wire a983, input wire b983,
  input wire a984, input wire b984,
  input wire a985, input wire b985,
  input wire a986, input wire b986,
  input wire a987, input wire b987,
  input wire a988, input wire b988,
  input wire a989, input wire b989,
  input wire a990, input wire b990,
  input wire a991, input wire b991,
  input wire a992, input wire b992,
  input wire a993, input wire b993,
  input wire a994, input wire b994,
  input wire a995, input wire b995,
  input wire a996, input wire b996,
  input wire a997, input wire b997,
  input wire a998, input wire b998,
  input wire a999, input wire b999,
  input wire a1000, input wire b1000,
  input wire a1001, input wire b1001,
  input wire a1002, input wire b1002,
  input wire a1003, input wire b1003,
  input wire a1004, input wire b1004,
  input wire a1005, input wire b1005,
  input wire a1006, input wire b1006,
  input wire a1007, input wire b1007,
  input wire a1008, input wire b1008,
  input wire a1009, input wire b1009,
  input wire a1010, input wire b1010,
  input wire a1011, input wire b1011,
  input wire a1012, input wire b1012,
  input wire a1013, input wire b1013,
  input wire a1014, input wire b1014,
  input wire a1015, input wire b1015,
  input wire a1016, input wire b1016,
  input wire a1017, input wire b1017,
  input wire a1018, input wire b1018,
  input wire a1019, input wire b1019,
  input wire a1020, input wire b1020,
  input wire a1021, input wire b1021,
  input wire a1022, input wire b1022,
  input wire a1023, input wire b1023,
  input wire op0,
  input wire op1,
  output wire y0,
  output wire y1,
  output wire y2,
  output wire y3,
  output wire y4,
  output wire y5,
  output wire y6,
  output wire y7,
  output wire y8,
  output wire y9,
  output wire y10,
  output wire y11,
  output wire y12,
  output wire y13,
  output wire y14,
  output wire y15,
  output wire y16,
  output wire y17,
  output wire y18,
  output wire y19,
  output wire y20,
  output wire y21,
  output wire y22,
  output wire y23,
  output wire y24,
  output wire y25,
  output wire y26,
  output wire y27,
  output wire y28,
  output wire y29,
  output wire y30,
  output wire y31,
  output wire y32,
  output wire y33,
  output wire y34,
  output wire y35,
  output wire y36,
  output wire y37,
  output wire y38,
  output wire y39,
  output wire y40,
  output wire y41,
  output wire y42,
  output wire y43,
  output wire y44,
  output wire y45,
  output wire y46,
  output wire y47,
  output wire y48,
  output wire y49,
  output wire y50,
  output wire y51,
  output wire y52,
  output wire y53,
  output wire y54,
  output wire y55,
  output wire y56,
  output wire y57,
  output wire y58,
  output wire y59,
  output wire y60,
  output wire y61,
  output wire y62,
  output wire y63,
  output wire y64,
  output wire y65,
  output wire y66,
  output wire y67,
  output wire y68,
  output wire y69,
  output wire y70,
  output wire y71,
  output wire y72,
  output wire y73,
  output wire y74,
  output wire y75,
  output wire y76,
  output wire y77,
  output wire y78,
  output wire y79,
  output wire y80,
  output wire y81,
  output wire y82,
  output wire y83,
  output wire y84,
  output wire y85,
  output wire y86,
  output wire y87,
  output wire y88,
  output wire y89,
  output wire y90,
  output wire y91,
  output wire y92,
  output wire y93,
  output wire y94,
  output wire y95,
  output wire y96,
  output wire y97,
  output wire y98,
  output wire y99,
  output wire y100,
  output wire y101,
  output wire y102,
  output wire y103,
  output wire y104,
  output wire y105,
  output wire y106,
  output wire y107,
  output wire y108,
  output wire y109,
  output wire y110,
  output wire y111,
  output wire y112,
  output wire y113,
  output wire y114,
  output wire y115,
  output wire y116,
  output wire y117,
  output wire y118,
  output wire y119,
  output wire y120,
  output wire y121,
  output wire y122,
  output wire y123,
  output wire y124,
  output wire y125,
  output wire y126,
  output wire y127,
  output wire y128,
  output wire y129,
  output wire y130,
  output wire y131,
  output wire y132,
  output wire y133,
  output wire y134,
  output wire y135,
  output wire y136,
  output wire y137,
  output wire y138,
  output wire y139,
  output wire y140,
  output wire y141,
  output wire y142,
  output wire y143,
  output wire y144,
  output wire y145,
  output wire y146,
  output wire y147,
  output wire y148,
  output wire y149,
  output wire y150,
  output wire y151,
  output wire y152,
  output wire y153,
  output wire y154,
  output wire y155,
  output wire y156,
  output wire y157,
  output wire y158,
  output wire y159,
  output wire y160,
  output wire y161,
  output wire y162,
  output wire y163,
  output wire y164,
  output wire y165,
  output wire y166,
  output wire y167,
  output wire y168,
  output wire y169,
  output wire y170,
  output wire y171,
  output wire y172,
  output wire y173,
  output wire y174,
  output wire y175,
  output wire y176,
  output wire y177,
  output wire y178,
  output wire y179,
  output wire y180,
  output wire y181,
  output wire y182,
  output wire y183,
  output wire y184,
  output wire y185,
  output wire y186,
  output wire y187,
  output wire y188,
  output wire y189,
  output wire y190,
  output wire y191,
  output wire y192,
  output wire y193,
  output wire y194,
  output wire y195,
  output wire y196,
  output wire y197,
  output wire y198,
  output wire y199,
  output wire y200,
  output wire y201,
  output wire y202,
  output wire y203,
  output wire y204,
  output wire y205,
  output wire y206,
  output wire y207,
  output wire y208,
  output wire y209,
  output wire y210,
  output wire y211,
  output wire y212,
  output wire y213,
  output wire y214,
  output wire y215,
  output wire y216,
  output wire y217,
  output wire y218,
  output wire y219,
  output wire y220,
  output wire y221,
  output wire y222,
  output wire y223,
  output wire y224,
  output wire y225,
  output wire y226,
  output wire y227,
  output wire y228,
  output wire y229,
  output wire y230,
  output wire y231,
  output wire y232,
  output wire y233,
  output wire y234,
  output wire y235,
  output wire y236,
  output wire y237,
  output wire y238,
  output wire y239,
  output wire y240,
  output wire y241,
  output wire y242,
  output wire y243,
  output wire y244,
  output wire y245,
  output wire y246,
  output wire y247,
  output wire y248,
  output wire y249,
  output wire y250,
  output wire y251,
  output wire y252,
  output wire y253,
  output wire y254,
  output wire y255,
  output wire y256,
  output wire y257,
  output wire y258,
  output wire y259,
  output wire y260,
  output wire y261,
  output wire y262,
  output wire y263,
  output wire y264,
  output wire y265,
  output wire y266,
  output wire y267,
  output wire y268,
  output wire y269,
  output wire y270,
  output wire y271,
  output wire y272,
  output wire y273,
  output wire y274,
  output wire y275,
  output wire y276,
  output wire y277,
  output wire y278,
  output wire y279,
  output wire y280,
  output wire y281,
  output wire y282,
  output wire y283,
  output wire y284,
  output wire y285,
  output wire y286,
  output wire y287,
  output wire y288,
  output wire y289,
  output wire y290,
  output wire y291,
  output wire y292,
  output wire y293,
  output wire y294,
  output wire y295,
  output wire y296,
  output wire y297,
  output wire y298,
  output wire y299,
  output wire y300,
  output wire y301,
  output wire y302,
  output wire y303,
  output wire y304,
  output wire y305,
  output wire y306,
  output wire y307,
  output wire y308,
  output wire y309,
  output wire y310,
  output wire y311,
  output wire y312,
  output wire y313,
  output wire y314,
  output wire y315,
  output wire y316,
  output wire y317,
  output wire y318,
  output wire y319,
  output wire y320,
  output wire y321,
  output wire y322,
  output wire y323,
  output wire y324,
  output wire y325,
  output wire y326,
  output wire y327,
  output wire y328,
  output wire y329,
  output wire y330,
  output wire y331,
  output wire y332,
  output wire y333,
  output wire y334,
  output wire y335,
  output wire y336,
  output wire y337,
  output wire y338,
  output wire y339,
  output wire y340,
  output wire y341,
  output wire y342,
  output wire y343,
  output wire y344,
  output wire y345,
  output wire y346,
  output wire y347,
  output wire y348,
  output wire y349,
  output wire y350,
  output wire y351,
  output wire y352,
  output wire y353,
  output wire y354,
  output wire y355,
  output wire y356,
  output wire y357,
  output wire y358,
  output wire y359,
  output wire y360,
  output wire y361,
  output wire y362,
  output wire y363,
  output wire y364,
  output wire y365,
  output wire y366,
  output wire y367,
  output wire y368,
  output wire y369,
  output wire y370,
  output wire y371,
  output wire y372,
  output wire y373,
  output wire y374,
  output wire y375,
  output wire y376,
  output wire y377,
  output wire y378,
  output wire y379,
  output wire y380,
  output wire y381,
  output wire y382,
  output wire y383,
  output wire y384,
  output wire y385,
  output wire y386,
  output wire y387,
  output wire y388,
  output wire y389,
  output wire y390,
  output wire y391,
  output wire y392,
  output wire y393,
  output wire y394,
  output wire y395,
  output wire y396,
  output wire y397,
  output wire y398,
  output wire y399,
  output wire y400,
  output wire y401,
  output wire y402,
  output wire y403,
  output wire y404,
  output wire y405,
  output wire y406,
  output wire y407,
  output wire y408,
  output wire y409,
  output wire y410,
  output wire y411,
  output wire y412,
  output wire y413,
  output wire y414,
  output wire y415,
  output wire y416,
  output wire y417,
  output wire y418,
  output wire y419,
  output wire y420,
  output wire y421,
  output wire y422,
  output wire y423,
  output wire y424,
  output wire y425,
  output wire y426,
  output wire y427,
  output wire y428,
  output wire y429,
  output wire y430,
  output wire y431,
  output wire y432,
  output wire y433,
  output wire y434,
  output wire y435,
  output wire y436,
  output wire y437,
  output wire y438,
  output wire y439,
  output wire y440,
  output wire y441,
  output wire y442,
  output wire y443,
  output wire y444,
  output wire y445,
  output wire y446,
  output wire y447,
  output wire y448,
  output wire y449,
  output wire y450,
  output wire y451,
  output wire y452,
  output wire y453,
  output wire y454,
  output wire y455,
  output wire y456,
  output wire y457,
  output wire y458,
  output wire y459,
  output wire y460,
  output wire y461,
  output wire y462,
  output wire y463,
  output wire y464,
  output wire y465,
  output wire y466,
  output wire y467,
  output wire y468,
  output wire y469,
  output wire y470,
  output wire y471,
  output wire y472,
  output wire y473,
  output wire y474,
  output wire y475,
  output wire y476,
  output wire y477,
  output wire y478,
  output wire y479,
  output wire y480,
  output wire y481,
  output wire y482,
  output wire y483,
  output wire y484,
  output wire y485,
  output wire y486,
  output wire y487,
  output wire y488,
  output wire y489,
  output wire y490,
  output wire y491,
  output wire y492,
  output wire y493,
  output wire y494,
  output wire y495,
  output wire y496,
  output wire y497,
  output wire y498,
  output wire y499,
  output wire y500,
  output wire y501,
  output wire y502,
  output wire y503,
  output wire y504,
  output wire y505,
  output wire y506,
  output wire y507,
  output wire y508,
  output wire y509,
  output wire y510,
  output wire y511,
  output wire y512,
  output wire y513,
  output wire y514,
  output wire y515,
  output wire y516,
  output wire y517,
  output wire y518,
  output wire y519,
  output wire y520,
  output wire y521,
  output wire y522,
  output wire y523,
  output wire y524,
  output wire y525,
  output wire y526,
  output wire y527,
  output wire y528,
  output wire y529,
  output wire y530,
  output wire y531,
  output wire y532,
  output wire y533,
  output wire y534,
  output wire y535,
  output wire y536,
  output wire y537,
  output wire y538,
  output wire y539,
  output wire y540,
  output wire y541,
  output wire y542,
  output wire y543,
  output wire y544,
  output wire y545,
  output wire y546,
  output wire y547,
  output wire y548,
  output wire y549,
  output wire y550,
  output wire y551,
  output wire y552,
  output wire y553,
  output wire y554,
  output wire y555,
  output wire y556,
  output wire y557,
  output wire y558,
  output wire y559,
  output wire y560,
  output wire y561,
  output wire y562,
  output wire y563,
  output wire y564,
  output wire y565,
  output wire y566,
  output wire y567,
  output wire y568,
  output wire y569,
  output wire y570,
  output wire y571,
  output wire y572,
  output wire y573,
  output wire y574,
  output wire y575,
  output wire y576,
  output wire y577,
  output wire y578,
  output wire y579,
  output wire y580,
  output wire y581,
  output wire y582,
  output wire y583,
  output wire y584,
  output wire y585,
  output wire y586,
  output wire y587,
  output wire y588,
  output wire y589,
  output wire y590,
  output wire y591,
  output wire y592,
  output wire y593,
  output wire y594,
  output wire y595,
  output wire y596,
  output wire y597,
  output wire y598,
  output wire y599,
  output wire y600,
  output wire y601,
  output wire y602,
  output wire y603,
  output wire y604,
  output wire y605,
  output wire y606,
  output wire y607,
  output wire y608,
  output wire y609,
  output wire y610,
  output wire y611,
  output wire y612,
  output wire y613,
  output wire y614,
  output wire y615,
  output wire y616,
  output wire y617,
  output wire y618,
  output wire y619,
  output wire y620,
  output wire y621,
  output wire y622,
  output wire y623,
  output wire y624,
  output wire y625,
  output wire y626,
  output wire y627,
  output wire y628,
  output wire y629,
  output wire y630,
  output wire y631,
  output wire y632,
  output wire y633,
  output wire y634,
  output wire y635,
  output wire y636,
  output wire y637,
  output wire y638,
  output wire y639,
  output wire y640,
  output wire y641,
  output wire y642,
  output wire y643,
  output wire y644,
  output wire y645,
  output wire y646,
  output wire y647,
  output wire y648,
  output wire y649,
  output wire y650,
  output wire y651,
  output wire y652,
  output wire y653,
  output wire y654,
  output wire y655,
  output wire y656,
  output wire y657,
  output wire y658,
  output wire y659,
  output wire y660,
  output wire y661,
  output wire y662,
  output wire y663,
  output wire y664,
  output wire y665,
  output wire y666,
  output wire y667,
  output wire y668,
  output wire y669,
  output wire y670,
  output wire y671,
  output wire y672,
  output wire y673,
  output wire y674,
  output wire y675,
  output wire y676,
  output wire y677,
  output wire y678,
  output wire y679,
  output wire y680,
  output wire y681,
  output wire y682,
  output wire y683,
  output wire y684,
  output wire y685,
  output wire y686,
  output wire y687,
  output wire y688,
  output wire y689,
  output wire y690,
  output wire y691,
  output wire y692,
  output wire y693,
  output wire y694,
  output wire y695,
  output wire y696,
  output wire y697,
  output wire y698,
  output wire y699,
  output wire y700,
  output wire y701,
  output wire y702,
  output wire y703,
  output wire y704,
  output wire y705,
  output wire y706,
  output wire y707,
  output wire y708,
  output wire y709,
  output wire y710,
  output wire y711,
  output wire y712,
  output wire y713,
  output wire y714,
  output wire y715,
  output wire y716,
  output wire y717,
  output wire y718,
  output wire y719,
  output wire y720,
  output wire y721,
  output wire y722,
  output wire y723,
  output wire y724,
  output wire y725,
  output wire y726,
  output wire y727,
  output wire y728,
  output wire y729,
  output wire y730,
  output wire y731,
  output wire y732,
  output wire y733,
  output wire y734,
  output wire y735,
  output wire y736,
  output wire y737,
  output wire y738,
  output wire y739,
  output wire y740,
  output wire y741,
  output wire y742,
  output wire y743,
  output wire y744,
  output wire y745,
  output wire y746,
  output wire y747,
  output wire y748,
  output wire y749,
  output wire y750,
  output wire y751,
  output wire y752,
  output wire y753,
  output wire y754,
  output wire y755,
  output wire y756,
  output wire y757,
  output wire y758,
  output wire y759,
  output wire y760,
  output wire y761,
  output wire y762,
  output wire y763,
  output wire y764,
  output wire y765,
  output wire y766,
  output wire y767,
  output wire y768,
  output wire y769,
  output wire y770,
  output wire y771,
  output wire y772,
  output wire y773,
  output wire y774,
  output wire y775,
  output wire y776,
  output wire y777,
  output wire y778,
  output wire y779,
  output wire y780,
  output wire y781,
  output wire y782,
  output wire y783,
  output wire y784,
  output wire y785,
  output wire y786,
  output wire y787,
  output wire y788,
  output wire y789,
  output wire y790,
  output wire y791,
  output wire y792,
  output wire y793,
  output wire y794,
  output wire y795,
  output wire y796,
  output wire y797,
  output wire y798,
  output wire y799,
  output wire y800,
  output wire y801,
  output wire y802,
  output wire y803,
  output wire y804,
  output wire y805,
  output wire y806,
  output wire y807,
  output wire y808,
  output wire y809,
  output wire y810,
  output wire y811,
  output wire y812,
  output wire y813,
  output wire y814,
  output wire y815,
  output wire y816,
  output wire y817,
  output wire y818,
  output wire y819,
  output wire y820,
  output wire y821,
  output wire y822,
  output wire y823,
  output wire y824,
  output wire y825,
  output wire y826,
  output wire y827,
  output wire y828,
  output wire y829,
  output wire y830,
  output wire y831,
  output wire y832,
  output wire y833,
  output wire y834,
  output wire y835,
  output wire y836,
  output wire y837,
  output wire y838,
  output wire y839,
  output wire y840,
  output wire y841,
  output wire y842,
  output wire y843,
  output wire y844,
  output wire y845,
  output wire y846,
  output wire y847,
  output wire y848,
  output wire y849,
  output wire y850,
  output wire y851,
  output wire y852,
  output wire y853,
  output wire y854,
  output wire y855,
  output wire y856,
  output wire y857,
  output wire y858,
  output wire y859,
  output wire y860,
  output wire y861,
  output wire y862,
  output wire y863,
  output wire y864,
  output wire y865,
  output wire y866,
  output wire y867,
  output wire y868,
  output wire y869,
  output wire y870,
  output wire y871,
  output wire y872,
  output wire y873,
  output wire y874,
  output wire y875,
  output wire y876,
  output wire y877,
  output wire y878,
  output wire y879,
  output wire y880,
  output wire y881,
  output wire y882,
  output wire y883,
  output wire y884,
  output wire y885,
  output wire y886,
  output wire y887,
  output wire y888,
  output wire y889,
  output wire y890,
  output wire y891,
  output wire y892,
  output wire y893,
  output wire y894,
  output wire y895,
  output wire y896,
  output wire y897,
  output wire y898,
  output wire y899,
  output wire y900,
  output wire y901,
  output wire y902,
  output wire y903,
  output wire y904,
  output wire y905,
  output wire y906,
  output wire y907,
  output wire y908,
  output wire y909,
  output wire y910,
  output wire y911,
  output wire y912,
  output wire y913,
  output wire y914,
  output wire y915,
  output wire y916,
  output wire y917,
  output wire y918,
  output wire y919,
  output wire y920,
  output wire y921,
  output wire y922,
  output wire y923,
  output wire y924,
  output wire y925,
  output wire y926,
  output wire y927,
  output wire y928,
  output wire y929,
  output wire y930,
  output wire y931,
  output wire y932,
  output wire y933,
  output wire y934,
  output wire y935,
  output wire y936,
  output wire y937,
  output wire y938,
  output wire y939,
  output wire y940,
  output wire y941,
  output wire y942,
  output wire y943,
  output wire y944,
  output wire y945,
  output wire y946,
  output wire y947,
  output wire y948,
  output wire y949,
  output wire y950,
  output wire y951,
  output wire y952,
  output wire y953,
  output wire y954,
  output wire y955,
  output wire y956,
  output wire y957,
  output wire y958,
  output wire y959,
  output wire y960,
  output wire y961,
  output wire y962,
  output wire y963,
  output wire y964,
  output wire y965,
  output wire y966,
  output wire y967,
  output wire y968,
  output wire y969,
  output wire y970,
  output wire y971,
  output wire y972,
  output wire y973,
  output wire y974,
  output wire y975,
  output wire y976,
  output wire y977,
  output wire y978,
  output wire y979,
  output wire y980,
  output wire y981,
  output wire y982,
  output wire y983,
  output wire y984,
  output wire y985,
  output wire y986,
  output wire y987,
  output wire y988,
  output wire y989,
  output wire y990,
  output wire y991,
  output wire y992,
  output wire y993,
  output wire y994,
  output wire y995,
  output wire y996,
  output wire y997,
  output wire y998,
  output wire y999,
  output wire y1000,
  output wire y1001,
  output wire y1002,
  output wire y1003,
  output wire y1004,
  output wire y1005,
  output wire y1006,
  output wire y1007,
  output wire y1008,
  output wire y1009,
  output wire y1010,
  output wire y1011,
  output wire y1012,
  output wire y1013,
  output wire y1014,
  output wire y1015,
  output wire y1016,
  output wire y1017,
  output wire y1018,
  output wire y1019,
  output wire y1020,
  output wire y1021,
  output wire y1022,
  output wire y1023
);
  wire add_sel, sub_sel, and_sel, or_sel;
  assign add_sel = ~op1 & ~op0;
  assign sub_sel = ~op1 & op0;
  assign and_sel = op1 & ~op0;
  assign or_sel  = op1 & op0;
  wire c0;
  wire c1;
  wire c2;
  wire c3;
  wire c4;
  wire c5;
  wire c6;
  wire c7;
  wire c8;
  wire c9;
  wire c10;
  wire c11;
  wire c12;
  wire c13;
  wire c14;
  wire c15;
  wire c16;
  wire c17;
  wire c18;
  wire c19;
  wire c20;
  wire c21;
  wire c22;
  wire c23;
  wire c24;
  wire c25;
  wire c26;
  wire c27;
  wire c28;
  wire c29;
  wire c30;
  wire c31;
  wire c32;
  wire c33;
  wire c34;
  wire c35;
  wire c36;
  wire c37;
  wire c38;
  wire c39;
  wire c40;
  wire c41;
  wire c42;
  wire c43;
  wire c44;
  wire c45;
  wire c46;
  wire c47;
  wire c48;
  wire c49;
  wire c50;
  wire c51;
  wire c52;
  wire c53;
  wire c54;
  wire c55;
  wire c56;
  wire c57;
  wire c58;
  wire c59;
  wire c60;
  wire c61;
  wire c62;
  wire c63;
  wire c64;
  wire c65;
  wire c66;
  wire c67;
  wire c68;
  wire c69;
  wire c70;
  wire c71;
  wire c72;
  wire c73;
  wire c74;
  wire c75;
  wire c76;
  wire c77;
  wire c78;
  wire c79;
  wire c80;
  wire c81;
  wire c82;
  wire c83;
  wire c84;
  wire c85;
  wire c86;
  wire c87;
  wire c88;
  wire c89;
  wire c90;
  wire c91;
  wire c92;
  wire c93;
  wire c94;
  wire c95;
  wire c96;
  wire c97;
  wire c98;
  wire c99;
  wire c100;
  wire c101;
  wire c102;
  wire c103;
  wire c104;
  wire c105;
  wire c106;
  wire c107;
  wire c108;
  wire c109;
  wire c110;
  wire c111;
  wire c112;
  wire c113;
  wire c114;
  wire c115;
  wire c116;
  wire c117;
  wire c118;
  wire c119;
  wire c120;
  wire c121;
  wire c122;
  wire c123;
  wire c124;
  wire c125;
  wire c126;
  wire c127;
  wire c128;
  wire c129;
  wire c130;
  wire c131;
  wire c132;
  wire c133;
  wire c134;
  wire c135;
  wire c136;
  wire c137;
  wire c138;
  wire c139;
  wire c140;
  wire c141;
  wire c142;
  wire c143;
  wire c144;
  wire c145;
  wire c146;
  wire c147;
  wire c148;
  wire c149;
  wire c150;
  wire c151;
  wire c152;
  wire c153;
  wire c154;
  wire c155;
  wire c156;
  wire c157;
  wire c158;
  wire c159;
  wire c160;
  wire c161;
  wire c162;
  wire c163;
  wire c164;
  wire c165;
  wire c166;
  wire c167;
  wire c168;
  wire c169;
  wire c170;
  wire c171;
  wire c172;
  wire c173;
  wire c174;
  wire c175;
  wire c176;
  wire c177;
  wire c178;
  wire c179;
  wire c180;
  wire c181;
  wire c182;
  wire c183;
  wire c184;
  wire c185;
  wire c186;
  wire c187;
  wire c188;
  wire c189;
  wire c190;
  wire c191;
  wire c192;
  wire c193;
  wire c194;
  wire c195;
  wire c196;
  wire c197;
  wire c198;
  wire c199;
  wire c200;
  wire c201;
  wire c202;
  wire c203;
  wire c204;
  wire c205;
  wire c206;
  wire c207;
  wire c208;
  wire c209;
  wire c210;
  wire c211;
  wire c212;
  wire c213;
  wire c214;
  wire c215;
  wire c216;
  wire c217;
  wire c218;
  wire c219;
  wire c220;
  wire c221;
  wire c222;
  wire c223;
  wire c224;
  wire c225;
  wire c226;
  wire c227;
  wire c228;
  wire c229;
  wire c230;
  wire c231;
  wire c232;
  wire c233;
  wire c234;
  wire c235;
  wire c236;
  wire c237;
  wire c238;
  wire c239;
  wire c240;
  wire c241;
  wire c242;
  wire c243;
  wire c244;
  wire c245;
  wire c246;
  wire c247;
  wire c248;
  wire c249;
  wire c250;
  wire c251;
  wire c252;
  wire c253;
  wire c254;
  wire c255;
  wire c256;
  wire c257;
  wire c258;
  wire c259;
  wire c260;
  wire c261;
  wire c262;
  wire c263;
  wire c264;
  wire c265;
  wire c266;
  wire c267;
  wire c268;
  wire c269;
  wire c270;
  wire c271;
  wire c272;
  wire c273;
  wire c274;
  wire c275;
  wire c276;
  wire c277;
  wire c278;
  wire c279;
  wire c280;
  wire c281;
  wire c282;
  wire c283;
  wire c284;
  wire c285;
  wire c286;
  wire c287;
  wire c288;
  wire c289;
  wire c290;
  wire c291;
  wire c292;
  wire c293;
  wire c294;
  wire c295;
  wire c296;
  wire c297;
  wire c298;
  wire c299;
  wire c300;
  wire c301;
  wire c302;
  wire c303;
  wire c304;
  wire c305;
  wire c306;
  wire c307;
  wire c308;
  wire c309;
  wire c310;
  wire c311;
  wire c312;
  wire c313;
  wire c314;
  wire c315;
  wire c316;
  wire c317;
  wire c318;
  wire c319;
  wire c320;
  wire c321;
  wire c322;
  wire c323;
  wire c324;
  wire c325;
  wire c326;
  wire c327;
  wire c328;
  wire c329;
  wire c330;
  wire c331;
  wire c332;
  wire c333;
  wire c334;
  wire c335;
  wire c336;
  wire c337;
  wire c338;
  wire c339;
  wire c340;
  wire c341;
  wire c342;
  wire c343;
  wire c344;
  wire c345;
  wire c346;
  wire c347;
  wire c348;
  wire c349;
  wire c350;
  wire c351;
  wire c352;
  wire c353;
  wire c354;
  wire c355;
  wire c356;
  wire c357;
  wire c358;
  wire c359;
  wire c360;
  wire c361;
  wire c362;
  wire c363;
  wire c364;
  wire c365;
  wire c366;
  wire c367;
  wire c368;
  wire c369;
  wire c370;
  wire c371;
  wire c372;
  wire c373;
  wire c374;
  wire c375;
  wire c376;
  wire c377;
  wire c378;
  wire c379;
  wire c380;
  wire c381;
  wire c382;
  wire c383;
  wire c384;
  wire c385;
  wire c386;
  wire c387;
  wire c388;
  wire c389;
  wire c390;
  wire c391;
  wire c392;
  wire c393;
  wire c394;
  wire c395;
  wire c396;
  wire c397;
  wire c398;
  wire c399;
  wire c400;
  wire c401;
  wire c402;
  wire c403;
  wire c404;
  wire c405;
  wire c406;
  wire c407;
  wire c408;
  wire c409;
  wire c410;
  wire c411;
  wire c412;
  wire c413;
  wire c414;
  wire c415;
  wire c416;
  wire c417;
  wire c418;
  wire c419;
  wire c420;
  wire c421;
  wire c422;
  wire c423;
  wire c424;
  wire c425;
  wire c426;
  wire c427;
  wire c428;
  wire c429;
  wire c430;
  wire c431;
  wire c432;
  wire c433;
  wire c434;
  wire c435;
  wire c436;
  wire c437;
  wire c438;
  wire c439;
  wire c440;
  wire c441;
  wire c442;
  wire c443;
  wire c444;
  wire c445;
  wire c446;
  wire c447;
  wire c448;
  wire c449;
  wire c450;
  wire c451;
  wire c452;
  wire c453;
  wire c454;
  wire c455;
  wire c456;
  wire c457;
  wire c458;
  wire c459;
  wire c460;
  wire c461;
  wire c462;
  wire c463;
  wire c464;
  wire c465;
  wire c466;
  wire c467;
  wire c468;
  wire c469;
  wire c470;
  wire c471;
  wire c472;
  wire c473;
  wire c474;
  wire c475;
  wire c476;
  wire c477;
  wire c478;
  wire c479;
  wire c480;
  wire c481;
  wire c482;
  wire c483;
  wire c484;
  wire c485;
  wire c486;
  wire c487;
  wire c488;
  wire c489;
  wire c490;
  wire c491;
  wire c492;
  wire c493;
  wire c494;
  wire c495;
  wire c496;
  wire c497;
  wire c498;
  wire c499;
  wire c500;
  wire c501;
  wire c502;
  wire c503;
  wire c504;
  wire c505;
  wire c506;
  wire c507;
  wire c508;
  wire c509;
  wire c510;
  wire c511;
  wire c512;
  wire c513;
  wire c514;
  wire c515;
  wire c516;
  wire c517;
  wire c518;
  wire c519;
  wire c520;
  wire c521;
  wire c522;
  wire c523;
  wire c524;
  wire c525;
  wire c526;
  wire c527;
  wire c528;
  wire c529;
  wire c530;
  wire c531;
  wire c532;
  wire c533;
  wire c534;
  wire c535;
  wire c536;
  wire c537;
  wire c538;
  wire c539;
  wire c540;
  wire c541;
  wire c542;
  wire c543;
  wire c544;
  wire c545;
  wire c546;
  wire c547;
  wire c548;
  wire c549;
  wire c550;
  wire c551;
  wire c552;
  wire c553;
  wire c554;
  wire c555;
  wire c556;
  wire c557;
  wire c558;
  wire c559;
  wire c560;
  wire c561;
  wire c562;
  wire c563;
  wire c564;
  wire c565;
  wire c566;
  wire c567;
  wire c568;
  wire c569;
  wire c570;
  wire c571;
  wire c572;
  wire c573;
  wire c574;
  wire c575;
  wire c576;
  wire c577;
  wire c578;
  wire c579;
  wire c580;
  wire c581;
  wire c582;
  wire c583;
  wire c584;
  wire c585;
  wire c586;
  wire c587;
  wire c588;
  wire c589;
  wire c590;
  wire c591;
  wire c592;
  wire c593;
  wire c594;
  wire c595;
  wire c596;
  wire c597;
  wire c598;
  wire c599;
  wire c600;
  wire c601;
  wire c602;
  wire c603;
  wire c604;
  wire c605;
  wire c606;
  wire c607;
  wire c608;
  wire c609;
  wire c610;
  wire c611;
  wire c612;
  wire c613;
  wire c614;
  wire c615;
  wire c616;
  wire c617;
  wire c618;
  wire c619;
  wire c620;
  wire c621;
  wire c622;
  wire c623;
  wire c624;
  wire c625;
  wire c626;
  wire c627;
  wire c628;
  wire c629;
  wire c630;
  wire c631;
  wire c632;
  wire c633;
  wire c634;
  wire c635;
  wire c636;
  wire c637;
  wire c638;
  wire c639;
  wire c640;
  wire c641;
  wire c642;
  wire c643;
  wire c644;
  wire c645;
  wire c646;
  wire c647;
  wire c648;
  wire c649;
  wire c650;
  wire c651;
  wire c652;
  wire c653;
  wire c654;
  wire c655;
  wire c656;
  wire c657;
  wire c658;
  wire c659;
  wire c660;
  wire c661;
  wire c662;
  wire c663;
  wire c664;
  wire c665;
  wire c666;
  wire c667;
  wire c668;
  wire c669;
  wire c670;
  wire c671;
  wire c672;
  wire c673;
  wire c674;
  wire c675;
  wire c676;
  wire c677;
  wire c678;
  wire c679;
  wire c680;
  wire c681;
  wire c682;
  wire c683;
  wire c684;
  wire c685;
  wire c686;
  wire c687;
  wire c688;
  wire c689;
  wire c690;
  wire c691;
  wire c692;
  wire c693;
  wire c694;
  wire c695;
  wire c696;
  wire c697;
  wire c698;
  wire c699;
  wire c700;
  wire c701;
  wire c702;
  wire c703;
  wire c704;
  wire c705;
  wire c706;
  wire c707;
  wire c708;
  wire c709;
  wire c710;
  wire c711;
  wire c712;
  wire c713;
  wire c714;
  wire c715;
  wire c716;
  wire c717;
  wire c718;
  wire c719;
  wire c720;
  wire c721;
  wire c722;
  wire c723;
  wire c724;
  wire c725;
  wire c726;
  wire c727;
  wire c728;
  wire c729;
  wire c730;
  wire c731;
  wire c732;
  wire c733;
  wire c734;
  wire c735;
  wire c736;
  wire c737;
  wire c738;
  wire c739;
  wire c740;
  wire c741;
  wire c742;
  wire c743;
  wire c744;
  wire c745;
  wire c746;
  wire c747;
  wire c748;
  wire c749;
  wire c750;
  wire c751;
  wire c752;
  wire c753;
  wire c754;
  wire c755;
  wire c756;
  wire c757;
  wire c758;
  wire c759;
  wire c760;
  wire c761;
  wire c762;
  wire c763;
  wire c764;
  wire c765;
  wire c766;
  wire c767;
  wire c768;
  wire c769;
  wire c770;
  wire c771;
  wire c772;
  wire c773;
  wire c774;
  wire c775;
  wire c776;
  wire c777;
  wire c778;
  wire c779;
  wire c780;
  wire c781;
  wire c782;
  wire c783;
  wire c784;
  wire c785;
  wire c786;
  wire c787;
  wire c788;
  wire c789;
  wire c790;
  wire c791;
  wire c792;
  wire c793;
  wire c794;
  wire c795;
  wire c796;
  wire c797;
  wire c798;
  wire c799;
  wire c800;
  wire c801;
  wire c802;
  wire c803;
  wire c804;
  wire c805;
  wire c806;
  wire c807;
  wire c808;
  wire c809;
  wire c810;
  wire c811;
  wire c812;
  wire c813;
  wire c814;
  wire c815;
  wire c816;
  wire c817;
  wire c818;
  wire c819;
  wire c820;
  wire c821;
  wire c822;
  wire c823;
  wire c824;
  wire c825;
  wire c826;
  wire c827;
  wire c828;
  wire c829;
  wire c830;
  wire c831;
  wire c832;
  wire c833;
  wire c834;
  wire c835;
  wire c836;
  wire c837;
  wire c838;
  wire c839;
  wire c840;
  wire c841;
  wire c842;
  wire c843;
  wire c844;
  wire c845;
  wire c846;
  wire c847;
  wire c848;
  wire c849;
  wire c850;
  wire c851;
  wire c852;
  wire c853;
  wire c854;
  wire c855;
  wire c856;
  wire c857;
  wire c858;
  wire c859;
  wire c860;
  wire c861;
  wire c862;
  wire c863;
  wire c864;
  wire c865;
  wire c866;
  wire c867;
  wire c868;
  wire c869;
  wire c870;
  wire c871;
  wire c872;
  wire c873;
  wire c874;
  wire c875;
  wire c876;
  wire c877;
  wire c878;
  wire c879;
  wire c880;
  wire c881;
  wire c882;
  wire c883;
  wire c884;
  wire c885;
  wire c886;
  wire c887;
  wire c888;
  wire c889;
  wire c890;
  wire c891;
  wire c892;
  wire c893;
  wire c894;
  wire c895;
  wire c896;
  wire c897;
  wire c898;
  wire c899;
  wire c900;
  wire c901;
  wire c902;
  wire c903;
  wire c904;
  wire c905;
  wire c906;
  wire c907;
  wire c908;
  wire c909;
  wire c910;
  wire c911;
  wire c912;
  wire c913;
  wire c914;
  wire c915;
  wire c916;
  wire c917;
  wire c918;
  wire c919;
  wire c920;
  wire c921;
  wire c922;
  wire c923;
  wire c924;
  wire c925;
  wire c926;
  wire c927;
  wire c928;
  wire c929;
  wire c930;
  wire c931;
  wire c932;
  wire c933;
  wire c934;
  wire c935;
  wire c936;
  wire c937;
  wire c938;
  wire c939;
  wire c940;
  wire c941;
  wire c942;
  wire c943;
  wire c944;
  wire c945;
  wire c946;
  wire c947;
  wire c948;
  wire c949;
  wire c950;
  wire c951;
  wire c952;
  wire c953;
  wire c954;
  wire c955;
  wire c956;
  wire c957;
  wire c958;
  wire c959;
  wire c960;
  wire c961;
  wire c962;
  wire c963;
  wire c964;
  wire c965;
  wire c966;
  wire c967;
  wire c968;
  wire c969;
  wire c970;
  wire c971;
  wire c972;
  wire c973;
  wire c974;
  wire c975;
  wire c976;
  wire c977;
  wire c978;
  wire c979;
  wire c980;
  wire c981;
  wire c982;
  wire c983;
  wire c984;
  wire c985;
  wire c986;
  wire c987;
  wire c988;
  wire c989;
  wire c990;
  wire c991;
  wire c992;
  wire c993;
  wire c994;
  wire c995;
  wire c996;
  wire c997;
  wire c998;
  wire c999;
  wire c1000;
  wire c1001;
  wire c1002;
  wire c1003;
  wire c1004;
  wire c1005;
  wire c1006;
  wire c1007;
  wire c1008;
  wire c1009;
  wire c1010;
  wire c1011;
  wire c1012;
  wire c1013;
  wire c1014;
  wire c1015;
  wire c1016;
  wire c1017;
  wire c1018;
  wire c1019;
  wire c1020;
  wire c1021;
  wire c1022;
  wire c1023;
  wire c1024;
  assign c0 = 1'b0;
  wire s0, sub0, and0, or0;
  wire b_inv0;
  assign b_inv0 = ~b0;
  assign s0  = a0 ^ b0 ^ c0;
  assign sub0 = a0 ^ b_inv0 ^ c0;
  assign and0 = a0 & b0;
  assign or0  = a0 | b0;
  assign c1 = (a0 & b0) | (a0 & c0) | (b0 & c0);
  wire c_sub1;
  assign c_sub1 = (a0 & b_inv0) | (a0 & c0) | (b_inv0 & c0);
  wire s1, sub1, and1, or1;
  wire b_inv1;
  assign b_inv1 = ~b1;
  assign s1  = a1 ^ b1 ^ c1;
  assign sub1 = a1 ^ b_inv1 ^ c1;
  assign and1 = a1 & b1;
  assign or1  = a1 | b1;
  assign c2 = (a1 & b1) | (a1 & c1) | (b1 & c1);
  wire c_sub2;
  assign c_sub2 = (a1 & b_inv1) | (a1 & c1) | (b_inv1 & c1);
  wire s2, sub2, and2, or2;
  wire b_inv2;
  assign b_inv2 = ~b2;
  assign s2  = a2 ^ b2 ^ c2;
  assign sub2 = a2 ^ b_inv2 ^ c2;
  assign and2 = a2 & b2;
  assign or2  = a2 | b2;
  assign c3 = (a2 & b2) | (a2 & c2) | (b2 & c2);
  wire c_sub3;
  assign c_sub3 = (a2 & b_inv2) | (a2 & c2) | (b_inv2 & c2);
  wire s3, sub3, and3, or3;
  wire b_inv3;
  assign b_inv3 = ~b3;
  assign s3  = a3 ^ b3 ^ c3;
  assign sub3 = a3 ^ b_inv3 ^ c3;
  assign and3 = a3 & b3;
  assign or3  = a3 | b3;
  assign c4 = (a3 & b3) | (a3 & c3) | (b3 & c3);
  wire c_sub4;
  assign c_sub4 = (a3 & b_inv3) | (a3 & c3) | (b_inv3 & c3);
  wire s4, sub4, and4, or4;
  wire b_inv4;
  assign b_inv4 = ~b4;
  assign s4  = a4 ^ b4 ^ c4;
  assign sub4 = a4 ^ b_inv4 ^ c4;
  assign and4 = a4 & b4;
  assign or4  = a4 | b4;
  assign c5 = (a4 & b4) | (a4 & c4) | (b4 & c4);
  wire c_sub5;
  assign c_sub5 = (a4 & b_inv4) | (a4 & c4) | (b_inv4 & c4);
  wire s5, sub5, and5, or5;
  wire b_inv5;
  assign b_inv5 = ~b5;
  assign s5  = a5 ^ b5 ^ c5;
  assign sub5 = a5 ^ b_inv5 ^ c5;
  assign and5 = a5 & b5;
  assign or5  = a5 | b5;
  assign c6 = (a5 & b5) | (a5 & c5) | (b5 & c5);
  wire c_sub6;
  assign c_sub6 = (a5 & b_inv5) | (a5 & c5) | (b_inv5 & c5);
  wire s6, sub6, and6, or6;
  wire b_inv6;
  assign b_inv6 = ~b6;
  assign s6  = a6 ^ b6 ^ c6;
  assign sub6 = a6 ^ b_inv6 ^ c6;
  assign and6 = a6 & b6;
  assign or6  = a6 | b6;
  assign c7 = (a6 & b6) | (a6 & c6) | (b6 & c6);
  wire c_sub7;
  assign c_sub7 = (a6 & b_inv6) | (a6 & c6) | (b_inv6 & c6);
  wire s7, sub7, and7, or7;
  wire b_inv7;
  assign b_inv7 = ~b7;
  assign s7  = a7 ^ b7 ^ c7;
  assign sub7 = a7 ^ b_inv7 ^ c7;
  assign and7 = a7 & b7;
  assign or7  = a7 | b7;
  assign c8 = (a7 & b7) | (a7 & c7) | (b7 & c7);
  wire c_sub8;
  assign c_sub8 = (a7 & b_inv7) | (a7 & c7) | (b_inv7 & c7);
  wire s8, sub8, and8, or8;
  wire b_inv8;
  assign b_inv8 = ~b8;
  assign s8  = a8 ^ b8 ^ c8;
  assign sub8 = a8 ^ b_inv8 ^ c8;
  assign and8 = a8 & b8;
  assign or8  = a8 | b8;
  assign c9 = (a8 & b8) | (a8 & c8) | (b8 & c8);
  wire c_sub9;
  assign c_sub9 = (a8 & b_inv8) | (a8 & c8) | (b_inv8 & c8);
  wire s9, sub9, and9, or9;
  wire b_inv9;
  assign b_inv9 = ~b9;
  assign s9  = a9 ^ b9 ^ c9;
  assign sub9 = a9 ^ b_inv9 ^ c9;
  assign and9 = a9 & b9;
  assign or9  = a9 | b9;
  assign c10 = (a9 & b9) | (a9 & c9) | (b9 & c9);
  wire c_sub10;
  assign c_sub10 = (a9 & b_inv9) | (a9 & c9) | (b_inv9 & c9);
  wire s10, sub10, and10, or10;
  wire b_inv10;
  assign b_inv10 = ~b10;
  assign s10  = a10 ^ b10 ^ c10;
  assign sub10 = a10 ^ b_inv10 ^ c10;
  assign and10 = a10 & b10;
  assign or10  = a10 | b10;
  assign c11 = (a10 & b10) | (a10 & c10) | (b10 & c10);
  wire c_sub11;
  assign c_sub11 = (a10 & b_inv10) | (a10 & c10) | (b_inv10 & c10);
  wire s11, sub11, and11, or11;
  wire b_inv11;
  assign b_inv11 = ~b11;
  assign s11  = a11 ^ b11 ^ c11;
  assign sub11 = a11 ^ b_inv11 ^ c11;
  assign and11 = a11 & b11;
  assign or11  = a11 | b11;
  assign c12 = (a11 & b11) | (a11 & c11) | (b11 & c11);
  wire c_sub12;
  assign c_sub12 = (a11 & b_inv11) | (a11 & c11) | (b_inv11 & c11);
  wire s12, sub12, and12, or12;
  wire b_inv12;
  assign b_inv12 = ~b12;
  assign s12  = a12 ^ b12 ^ c12;
  assign sub12 = a12 ^ b_inv12 ^ c12;
  assign and12 = a12 & b12;
  assign or12  = a12 | b12;
  assign c13 = (a12 & b12) | (a12 & c12) | (b12 & c12);
  wire c_sub13;
  assign c_sub13 = (a12 & b_inv12) | (a12 & c12) | (b_inv12 & c12);
  wire s13, sub13, and13, or13;
  wire b_inv13;
  assign b_inv13 = ~b13;
  assign s13  = a13 ^ b13 ^ c13;
  assign sub13 = a13 ^ b_inv13 ^ c13;
  assign and13 = a13 & b13;
  assign or13  = a13 | b13;
  assign c14 = (a13 & b13) | (a13 & c13) | (b13 & c13);
  wire c_sub14;
  assign c_sub14 = (a13 & b_inv13) | (a13 & c13) | (b_inv13 & c13);
  wire s14, sub14, and14, or14;
  wire b_inv14;
  assign b_inv14 = ~b14;
  assign s14  = a14 ^ b14 ^ c14;
  assign sub14 = a14 ^ b_inv14 ^ c14;
  assign and14 = a14 & b14;
  assign or14  = a14 | b14;
  assign c15 = (a14 & b14) | (a14 & c14) | (b14 & c14);
  wire c_sub15;
  assign c_sub15 = (a14 & b_inv14) | (a14 & c14) | (b_inv14 & c14);
  wire s15, sub15, and15, or15;
  wire b_inv15;
  assign b_inv15 = ~b15;
  assign s15  = a15 ^ b15 ^ c15;
  assign sub15 = a15 ^ b_inv15 ^ c15;
  assign and15 = a15 & b15;
  assign or15  = a15 | b15;
  assign c16 = (a15 & b15) | (a15 & c15) | (b15 & c15);
  wire c_sub16;
  assign c_sub16 = (a15 & b_inv15) | (a15 & c15) | (b_inv15 & c15);
  wire s16, sub16, and16, or16;
  wire b_inv16;
  assign b_inv16 = ~b16;
  assign s16  = a16 ^ b16 ^ c16;
  assign sub16 = a16 ^ b_inv16 ^ c16;
  assign and16 = a16 & b16;
  assign or16  = a16 | b16;
  assign c17 = (a16 & b16) | (a16 & c16) | (b16 & c16);
  wire c_sub17;
  assign c_sub17 = (a16 & b_inv16) | (a16 & c16) | (b_inv16 & c16);
  wire s17, sub17, and17, or17;
  wire b_inv17;
  assign b_inv17 = ~b17;
  assign s17  = a17 ^ b17 ^ c17;
  assign sub17 = a17 ^ b_inv17 ^ c17;
  assign and17 = a17 & b17;
  assign or17  = a17 | b17;
  assign c18 = (a17 & b17) | (a17 & c17) | (b17 & c17);
  wire c_sub18;
  assign c_sub18 = (a17 & b_inv17) | (a17 & c17) | (b_inv17 & c17);
  wire s18, sub18, and18, or18;
  wire b_inv18;
  assign b_inv18 = ~b18;
  assign s18  = a18 ^ b18 ^ c18;
  assign sub18 = a18 ^ b_inv18 ^ c18;
  assign and18 = a18 & b18;
  assign or18  = a18 | b18;
  assign c19 = (a18 & b18) | (a18 & c18) | (b18 & c18);
  wire c_sub19;
  assign c_sub19 = (a18 & b_inv18) | (a18 & c18) | (b_inv18 & c18);
  wire s19, sub19, and19, or19;
  wire b_inv19;
  assign b_inv19 = ~b19;
  assign s19  = a19 ^ b19 ^ c19;
  assign sub19 = a19 ^ b_inv19 ^ c19;
  assign and19 = a19 & b19;
  assign or19  = a19 | b19;
  assign c20 = (a19 & b19) | (a19 & c19) | (b19 & c19);
  wire c_sub20;
  assign c_sub20 = (a19 & b_inv19) | (a19 & c19) | (b_inv19 & c19);
  wire s20, sub20, and20, or20;
  wire b_inv20;
  assign b_inv20 = ~b20;
  assign s20  = a20 ^ b20 ^ c20;
  assign sub20 = a20 ^ b_inv20 ^ c20;
  assign and20 = a20 & b20;
  assign or20  = a20 | b20;
  assign c21 = (a20 & b20) | (a20 & c20) | (b20 & c20);
  wire c_sub21;
  assign c_sub21 = (a20 & b_inv20) | (a20 & c20) | (b_inv20 & c20);
  wire s21, sub21, and21, or21;
  wire b_inv21;
  assign b_inv21 = ~b21;
  assign s21  = a21 ^ b21 ^ c21;
  assign sub21 = a21 ^ b_inv21 ^ c21;
  assign and21 = a21 & b21;
  assign or21  = a21 | b21;
  assign c22 = (a21 & b21) | (a21 & c21) | (b21 & c21);
  wire c_sub22;
  assign c_sub22 = (a21 & b_inv21) | (a21 & c21) | (b_inv21 & c21);
  wire s22, sub22, and22, or22;
  wire b_inv22;
  assign b_inv22 = ~b22;
  assign s22  = a22 ^ b22 ^ c22;
  assign sub22 = a22 ^ b_inv22 ^ c22;
  assign and22 = a22 & b22;
  assign or22  = a22 | b22;
  assign c23 = (a22 & b22) | (a22 & c22) | (b22 & c22);
  wire c_sub23;
  assign c_sub23 = (a22 & b_inv22) | (a22 & c22) | (b_inv22 & c22);
  wire s23, sub23, and23, or23;
  wire b_inv23;
  assign b_inv23 = ~b23;
  assign s23  = a23 ^ b23 ^ c23;
  assign sub23 = a23 ^ b_inv23 ^ c23;
  assign and23 = a23 & b23;
  assign or23  = a23 | b23;
  assign c24 = (a23 & b23) | (a23 & c23) | (b23 & c23);
  wire c_sub24;
  assign c_sub24 = (a23 & b_inv23) | (a23 & c23) | (b_inv23 & c23);
  wire s24, sub24, and24, or24;
  wire b_inv24;
  assign b_inv24 = ~b24;
  assign s24  = a24 ^ b24 ^ c24;
  assign sub24 = a24 ^ b_inv24 ^ c24;
  assign and24 = a24 & b24;
  assign or24  = a24 | b24;
  assign c25 = (a24 & b24) | (a24 & c24) | (b24 & c24);
  wire c_sub25;
  assign c_sub25 = (a24 & b_inv24) | (a24 & c24) | (b_inv24 & c24);
  wire s25, sub25, and25, or25;
  wire b_inv25;
  assign b_inv25 = ~b25;
  assign s25  = a25 ^ b25 ^ c25;
  assign sub25 = a25 ^ b_inv25 ^ c25;
  assign and25 = a25 & b25;
  assign or25  = a25 | b25;
  assign c26 = (a25 & b25) | (a25 & c25) | (b25 & c25);
  wire c_sub26;
  assign c_sub26 = (a25 & b_inv25) | (a25 & c25) | (b_inv25 & c25);
  wire s26, sub26, and26, or26;
  wire b_inv26;
  assign b_inv26 = ~b26;
  assign s26  = a26 ^ b26 ^ c26;
  assign sub26 = a26 ^ b_inv26 ^ c26;
  assign and26 = a26 & b26;
  assign or26  = a26 | b26;
  assign c27 = (a26 & b26) | (a26 & c26) | (b26 & c26);
  wire c_sub27;
  assign c_sub27 = (a26 & b_inv26) | (a26 & c26) | (b_inv26 & c26);
  wire s27, sub27, and27, or27;
  wire b_inv27;
  assign b_inv27 = ~b27;
  assign s27  = a27 ^ b27 ^ c27;
  assign sub27 = a27 ^ b_inv27 ^ c27;
  assign and27 = a27 & b27;
  assign or27  = a27 | b27;
  assign c28 = (a27 & b27) | (a27 & c27) | (b27 & c27);
  wire c_sub28;
  assign c_sub28 = (a27 & b_inv27) | (a27 & c27) | (b_inv27 & c27);
  wire s28, sub28, and28, or28;
  wire b_inv28;
  assign b_inv28 = ~b28;
  assign s28  = a28 ^ b28 ^ c28;
  assign sub28 = a28 ^ b_inv28 ^ c28;
  assign and28 = a28 & b28;
  assign or28  = a28 | b28;
  assign c29 = (a28 & b28) | (a28 & c28) | (b28 & c28);
  wire c_sub29;
  assign c_sub29 = (a28 & b_inv28) | (a28 & c28) | (b_inv28 & c28);
  wire s29, sub29, and29, or29;
  wire b_inv29;
  assign b_inv29 = ~b29;
  assign s29  = a29 ^ b29 ^ c29;
  assign sub29 = a29 ^ b_inv29 ^ c29;
  assign and29 = a29 & b29;
  assign or29  = a29 | b29;
  assign c30 = (a29 & b29) | (a29 & c29) | (b29 & c29);
  wire c_sub30;
  assign c_sub30 = (a29 & b_inv29) | (a29 & c29) | (b_inv29 & c29);
  wire s30, sub30, and30, or30;
  wire b_inv30;
  assign b_inv30 = ~b30;
  assign s30  = a30 ^ b30 ^ c30;
  assign sub30 = a30 ^ b_inv30 ^ c30;
  assign and30 = a30 & b30;
  assign or30  = a30 | b30;
  assign c31 = (a30 & b30) | (a30 & c30) | (b30 & c30);
  wire c_sub31;
  assign c_sub31 = (a30 & b_inv30) | (a30 & c30) | (b_inv30 & c30);
  wire s31, sub31, and31, or31;
  wire b_inv31;
  assign b_inv31 = ~b31;
  assign s31  = a31 ^ b31 ^ c31;
  assign sub31 = a31 ^ b_inv31 ^ c31;
  assign and31 = a31 & b31;
  assign or31  = a31 | b31;
  assign c32 = (a31 & b31) | (a31 & c31) | (b31 & c31);
  wire c_sub32;
  assign c_sub32 = (a31 & b_inv31) | (a31 & c31) | (b_inv31 & c31);
  wire s32, sub32, and32, or32;
  wire b_inv32;
  assign b_inv32 = ~b32;
  assign s32  = a32 ^ b32 ^ c32;
  assign sub32 = a32 ^ b_inv32 ^ c32;
  assign and32 = a32 & b32;
  assign or32  = a32 | b32;
  assign c33 = (a32 & b32) | (a32 & c32) | (b32 & c32);
  wire c_sub33;
  assign c_sub33 = (a32 & b_inv32) | (a32 & c32) | (b_inv32 & c32);
  wire s33, sub33, and33, or33;
  wire b_inv33;
  assign b_inv33 = ~b33;
  assign s33  = a33 ^ b33 ^ c33;
  assign sub33 = a33 ^ b_inv33 ^ c33;
  assign and33 = a33 & b33;
  assign or33  = a33 | b33;
  assign c34 = (a33 & b33) | (a33 & c33) | (b33 & c33);
  wire c_sub34;
  assign c_sub34 = (a33 & b_inv33) | (a33 & c33) | (b_inv33 & c33);
  wire s34, sub34, and34, or34;
  wire b_inv34;
  assign b_inv34 = ~b34;
  assign s34  = a34 ^ b34 ^ c34;
  assign sub34 = a34 ^ b_inv34 ^ c34;
  assign and34 = a34 & b34;
  assign or34  = a34 | b34;
  assign c35 = (a34 & b34) | (a34 & c34) | (b34 & c34);
  wire c_sub35;
  assign c_sub35 = (a34 & b_inv34) | (a34 & c34) | (b_inv34 & c34);
  wire s35, sub35, and35, or35;
  wire b_inv35;
  assign b_inv35 = ~b35;
  assign s35  = a35 ^ b35 ^ c35;
  assign sub35 = a35 ^ b_inv35 ^ c35;
  assign and35 = a35 & b35;
  assign or35  = a35 | b35;
  assign c36 = (a35 & b35) | (a35 & c35) | (b35 & c35);
  wire c_sub36;
  assign c_sub36 = (a35 & b_inv35) | (a35 & c35) | (b_inv35 & c35);
  wire s36, sub36, and36, or36;
  wire b_inv36;
  assign b_inv36 = ~b36;
  assign s36  = a36 ^ b36 ^ c36;
  assign sub36 = a36 ^ b_inv36 ^ c36;
  assign and36 = a36 & b36;
  assign or36  = a36 | b36;
  assign c37 = (a36 & b36) | (a36 & c36) | (b36 & c36);
  wire c_sub37;
  assign c_sub37 = (a36 & b_inv36) | (a36 & c36) | (b_inv36 & c36);
  wire s37, sub37, and37, or37;
  wire b_inv37;
  assign b_inv37 = ~b37;
  assign s37  = a37 ^ b37 ^ c37;
  assign sub37 = a37 ^ b_inv37 ^ c37;
  assign and37 = a37 & b37;
  assign or37  = a37 | b37;
  assign c38 = (a37 & b37) | (a37 & c37) | (b37 & c37);
  wire c_sub38;
  assign c_sub38 = (a37 & b_inv37) | (a37 & c37) | (b_inv37 & c37);
  wire s38, sub38, and38, or38;
  wire b_inv38;
  assign b_inv38 = ~b38;
  assign s38  = a38 ^ b38 ^ c38;
  assign sub38 = a38 ^ b_inv38 ^ c38;
  assign and38 = a38 & b38;
  assign or38  = a38 | b38;
  assign c39 = (a38 & b38) | (a38 & c38) | (b38 & c38);
  wire c_sub39;
  assign c_sub39 = (a38 & b_inv38) | (a38 & c38) | (b_inv38 & c38);
  wire s39, sub39, and39, or39;
  wire b_inv39;
  assign b_inv39 = ~b39;
  assign s39  = a39 ^ b39 ^ c39;
  assign sub39 = a39 ^ b_inv39 ^ c39;
  assign and39 = a39 & b39;
  assign or39  = a39 | b39;
  assign c40 = (a39 & b39) | (a39 & c39) | (b39 & c39);
  wire c_sub40;
  assign c_sub40 = (a39 & b_inv39) | (a39 & c39) | (b_inv39 & c39);
  wire s40, sub40, and40, or40;
  wire b_inv40;
  assign b_inv40 = ~b40;
  assign s40  = a40 ^ b40 ^ c40;
  assign sub40 = a40 ^ b_inv40 ^ c40;
  assign and40 = a40 & b40;
  assign or40  = a40 | b40;
  assign c41 = (a40 & b40) | (a40 & c40) | (b40 & c40);
  wire c_sub41;
  assign c_sub41 = (a40 & b_inv40) | (a40 & c40) | (b_inv40 & c40);
  wire s41, sub41, and41, or41;
  wire b_inv41;
  assign b_inv41 = ~b41;
  assign s41  = a41 ^ b41 ^ c41;
  assign sub41 = a41 ^ b_inv41 ^ c41;
  assign and41 = a41 & b41;
  assign or41  = a41 | b41;
  assign c42 = (a41 & b41) | (a41 & c41) | (b41 & c41);
  wire c_sub42;
  assign c_sub42 = (a41 & b_inv41) | (a41 & c41) | (b_inv41 & c41);
  wire s42, sub42, and42, or42;
  wire b_inv42;
  assign b_inv42 = ~b42;
  assign s42  = a42 ^ b42 ^ c42;
  assign sub42 = a42 ^ b_inv42 ^ c42;
  assign and42 = a42 & b42;
  assign or42  = a42 | b42;
  assign c43 = (a42 & b42) | (a42 & c42) | (b42 & c42);
  wire c_sub43;
  assign c_sub43 = (a42 & b_inv42) | (a42 & c42) | (b_inv42 & c42);
  wire s43, sub43, and43, or43;
  wire b_inv43;
  assign b_inv43 = ~b43;
  assign s43  = a43 ^ b43 ^ c43;
  assign sub43 = a43 ^ b_inv43 ^ c43;
  assign and43 = a43 & b43;
  assign or43  = a43 | b43;
  assign c44 = (a43 & b43) | (a43 & c43) | (b43 & c43);
  wire c_sub44;
  assign c_sub44 = (a43 & b_inv43) | (a43 & c43) | (b_inv43 & c43);
  wire s44, sub44, and44, or44;
  wire b_inv44;
  assign b_inv44 = ~b44;
  assign s44  = a44 ^ b44 ^ c44;
  assign sub44 = a44 ^ b_inv44 ^ c44;
  assign and44 = a44 & b44;
  assign or44  = a44 | b44;
  assign c45 = (a44 & b44) | (a44 & c44) | (b44 & c44);
  wire c_sub45;
  assign c_sub45 = (a44 & b_inv44) | (a44 & c44) | (b_inv44 & c44);
  wire s45, sub45, and45, or45;
  wire b_inv45;
  assign b_inv45 = ~b45;
  assign s45  = a45 ^ b45 ^ c45;
  assign sub45 = a45 ^ b_inv45 ^ c45;
  assign and45 = a45 & b45;
  assign or45  = a45 | b45;
  assign c46 = (a45 & b45) | (a45 & c45) | (b45 & c45);
  wire c_sub46;
  assign c_sub46 = (a45 & b_inv45) | (a45 & c45) | (b_inv45 & c45);
  wire s46, sub46, and46, or46;
  wire b_inv46;
  assign b_inv46 = ~b46;
  assign s46  = a46 ^ b46 ^ c46;
  assign sub46 = a46 ^ b_inv46 ^ c46;
  assign and46 = a46 & b46;
  assign or46  = a46 | b46;
  assign c47 = (a46 & b46) | (a46 & c46) | (b46 & c46);
  wire c_sub47;
  assign c_sub47 = (a46 & b_inv46) | (a46 & c46) | (b_inv46 & c46);
  wire s47, sub47, and47, or47;
  wire b_inv47;
  assign b_inv47 = ~b47;
  assign s47  = a47 ^ b47 ^ c47;
  assign sub47 = a47 ^ b_inv47 ^ c47;
  assign and47 = a47 & b47;
  assign or47  = a47 | b47;
  assign c48 = (a47 & b47) | (a47 & c47) | (b47 & c47);
  wire c_sub48;
  assign c_sub48 = (a47 & b_inv47) | (a47 & c47) | (b_inv47 & c47);
  wire s48, sub48, and48, or48;
  wire b_inv48;
  assign b_inv48 = ~b48;
  assign s48  = a48 ^ b48 ^ c48;
  assign sub48 = a48 ^ b_inv48 ^ c48;
  assign and48 = a48 & b48;
  assign or48  = a48 | b48;
  assign c49 = (a48 & b48) | (a48 & c48) | (b48 & c48);
  wire c_sub49;
  assign c_sub49 = (a48 & b_inv48) | (a48 & c48) | (b_inv48 & c48);
  wire s49, sub49, and49, or49;
  wire b_inv49;
  assign b_inv49 = ~b49;
  assign s49  = a49 ^ b49 ^ c49;
  assign sub49 = a49 ^ b_inv49 ^ c49;
  assign and49 = a49 & b49;
  assign or49  = a49 | b49;
  assign c50 = (a49 & b49) | (a49 & c49) | (b49 & c49);
  wire c_sub50;
  assign c_sub50 = (a49 & b_inv49) | (a49 & c49) | (b_inv49 & c49);
  wire s50, sub50, and50, or50;
  wire b_inv50;
  assign b_inv50 = ~b50;
  assign s50  = a50 ^ b50 ^ c50;
  assign sub50 = a50 ^ b_inv50 ^ c50;
  assign and50 = a50 & b50;
  assign or50  = a50 | b50;
  assign c51 = (a50 & b50) | (a50 & c50) | (b50 & c50);
  wire c_sub51;
  assign c_sub51 = (a50 & b_inv50) | (a50 & c50) | (b_inv50 & c50);
  wire s51, sub51, and51, or51;
  wire b_inv51;
  assign b_inv51 = ~b51;
  assign s51  = a51 ^ b51 ^ c51;
  assign sub51 = a51 ^ b_inv51 ^ c51;
  assign and51 = a51 & b51;
  assign or51  = a51 | b51;
  assign c52 = (a51 & b51) | (a51 & c51) | (b51 & c51);
  wire c_sub52;
  assign c_sub52 = (a51 & b_inv51) | (a51 & c51) | (b_inv51 & c51);
  wire s52, sub52, and52, or52;
  wire b_inv52;
  assign b_inv52 = ~b52;
  assign s52  = a52 ^ b52 ^ c52;
  assign sub52 = a52 ^ b_inv52 ^ c52;
  assign and52 = a52 & b52;
  assign or52  = a52 | b52;
  assign c53 = (a52 & b52) | (a52 & c52) | (b52 & c52);
  wire c_sub53;
  assign c_sub53 = (a52 & b_inv52) | (a52 & c52) | (b_inv52 & c52);
  wire s53, sub53, and53, or53;
  wire b_inv53;
  assign b_inv53 = ~b53;
  assign s53  = a53 ^ b53 ^ c53;
  assign sub53 = a53 ^ b_inv53 ^ c53;
  assign and53 = a53 & b53;
  assign or53  = a53 | b53;
  assign c54 = (a53 & b53) | (a53 & c53) | (b53 & c53);
  wire c_sub54;
  assign c_sub54 = (a53 & b_inv53) | (a53 & c53) | (b_inv53 & c53);
  wire s54, sub54, and54, or54;
  wire b_inv54;
  assign b_inv54 = ~b54;
  assign s54  = a54 ^ b54 ^ c54;
  assign sub54 = a54 ^ b_inv54 ^ c54;
  assign and54 = a54 & b54;
  assign or54  = a54 | b54;
  assign c55 = (a54 & b54) | (a54 & c54) | (b54 & c54);
  wire c_sub55;
  assign c_sub55 = (a54 & b_inv54) | (a54 & c54) | (b_inv54 & c54);
  wire s55, sub55, and55, or55;
  wire b_inv55;
  assign b_inv55 = ~b55;
  assign s55  = a55 ^ b55 ^ c55;
  assign sub55 = a55 ^ b_inv55 ^ c55;
  assign and55 = a55 & b55;
  assign or55  = a55 | b55;
  assign c56 = (a55 & b55) | (a55 & c55) | (b55 & c55);
  wire c_sub56;
  assign c_sub56 = (a55 & b_inv55) | (a55 & c55) | (b_inv55 & c55);
  wire s56, sub56, and56, or56;
  wire b_inv56;
  assign b_inv56 = ~b56;
  assign s56  = a56 ^ b56 ^ c56;
  assign sub56 = a56 ^ b_inv56 ^ c56;
  assign and56 = a56 & b56;
  assign or56  = a56 | b56;
  assign c57 = (a56 & b56) | (a56 & c56) | (b56 & c56);
  wire c_sub57;
  assign c_sub57 = (a56 & b_inv56) | (a56 & c56) | (b_inv56 & c56);
  wire s57, sub57, and57, or57;
  wire b_inv57;
  assign b_inv57 = ~b57;
  assign s57  = a57 ^ b57 ^ c57;
  assign sub57 = a57 ^ b_inv57 ^ c57;
  assign and57 = a57 & b57;
  assign or57  = a57 | b57;
  assign c58 = (a57 & b57) | (a57 & c57) | (b57 & c57);
  wire c_sub58;
  assign c_sub58 = (a57 & b_inv57) | (a57 & c57) | (b_inv57 & c57);
  wire s58, sub58, and58, or58;
  wire b_inv58;
  assign b_inv58 = ~b58;
  assign s58  = a58 ^ b58 ^ c58;
  assign sub58 = a58 ^ b_inv58 ^ c58;
  assign and58 = a58 & b58;
  assign or58  = a58 | b58;
  assign c59 = (a58 & b58) | (a58 & c58) | (b58 & c58);
  wire c_sub59;
  assign c_sub59 = (a58 & b_inv58) | (a58 & c58) | (b_inv58 & c58);
  wire s59, sub59, and59, or59;
  wire b_inv59;
  assign b_inv59 = ~b59;
  assign s59  = a59 ^ b59 ^ c59;
  assign sub59 = a59 ^ b_inv59 ^ c59;
  assign and59 = a59 & b59;
  assign or59  = a59 | b59;
  assign c60 = (a59 & b59) | (a59 & c59) | (b59 & c59);
  wire c_sub60;
  assign c_sub60 = (a59 & b_inv59) | (a59 & c59) | (b_inv59 & c59);
  wire s60, sub60, and60, or60;
  wire b_inv60;
  assign b_inv60 = ~b60;
  assign s60  = a60 ^ b60 ^ c60;
  assign sub60 = a60 ^ b_inv60 ^ c60;
  assign and60 = a60 & b60;
  assign or60  = a60 | b60;
  assign c61 = (a60 & b60) | (a60 & c60) | (b60 & c60);
  wire c_sub61;
  assign c_sub61 = (a60 & b_inv60) | (a60 & c60) | (b_inv60 & c60);
  wire s61, sub61, and61, or61;
  wire b_inv61;
  assign b_inv61 = ~b61;
  assign s61  = a61 ^ b61 ^ c61;
  assign sub61 = a61 ^ b_inv61 ^ c61;
  assign and61 = a61 & b61;
  assign or61  = a61 | b61;
  assign c62 = (a61 & b61) | (a61 & c61) | (b61 & c61);
  wire c_sub62;
  assign c_sub62 = (a61 & b_inv61) | (a61 & c61) | (b_inv61 & c61);
  wire s62, sub62, and62, or62;
  wire b_inv62;
  assign b_inv62 = ~b62;
  assign s62  = a62 ^ b62 ^ c62;
  assign sub62 = a62 ^ b_inv62 ^ c62;
  assign and62 = a62 & b62;
  assign or62  = a62 | b62;
  assign c63 = (a62 & b62) | (a62 & c62) | (b62 & c62);
  wire c_sub63;
  assign c_sub63 = (a62 & b_inv62) | (a62 & c62) | (b_inv62 & c62);
  wire s63, sub63, and63, or63;
  wire b_inv63;
  assign b_inv63 = ~b63;
  assign s63  = a63 ^ b63 ^ c63;
  assign sub63 = a63 ^ b_inv63 ^ c63;
  assign and63 = a63 & b63;
  assign or63  = a63 | b63;
  assign c64 = (a63 & b63) | (a63 & c63) | (b63 & c63);
  wire c_sub64;
  assign c_sub64 = (a63 & b_inv63) | (a63 & c63) | (b_inv63 & c63);
  wire s64, sub64, and64, or64;
  wire b_inv64;
  assign b_inv64 = ~b64;
  assign s64  = a64 ^ b64 ^ c64;
  assign sub64 = a64 ^ b_inv64 ^ c64;
  assign and64 = a64 & b64;
  assign or64  = a64 | b64;
  assign c65 = (a64 & b64) | (a64 & c64) | (b64 & c64);
  wire c_sub65;
  assign c_sub65 = (a64 & b_inv64) | (a64 & c64) | (b_inv64 & c64);
  wire s65, sub65, and65, or65;
  wire b_inv65;
  assign b_inv65 = ~b65;
  assign s65  = a65 ^ b65 ^ c65;
  assign sub65 = a65 ^ b_inv65 ^ c65;
  assign and65 = a65 & b65;
  assign or65  = a65 | b65;
  assign c66 = (a65 & b65) | (a65 & c65) | (b65 & c65);
  wire c_sub66;
  assign c_sub66 = (a65 & b_inv65) | (a65 & c65) | (b_inv65 & c65);
  wire s66, sub66, and66, or66;
  wire b_inv66;
  assign b_inv66 = ~b66;
  assign s66  = a66 ^ b66 ^ c66;
  assign sub66 = a66 ^ b_inv66 ^ c66;
  assign and66 = a66 & b66;
  assign or66  = a66 | b66;
  assign c67 = (a66 & b66) | (a66 & c66) | (b66 & c66);
  wire c_sub67;
  assign c_sub67 = (a66 & b_inv66) | (a66 & c66) | (b_inv66 & c66);
  wire s67, sub67, and67, or67;
  wire b_inv67;
  assign b_inv67 = ~b67;
  assign s67  = a67 ^ b67 ^ c67;
  assign sub67 = a67 ^ b_inv67 ^ c67;
  assign and67 = a67 & b67;
  assign or67  = a67 | b67;
  assign c68 = (a67 & b67) | (a67 & c67) | (b67 & c67);
  wire c_sub68;
  assign c_sub68 = (a67 & b_inv67) | (a67 & c67) | (b_inv67 & c67);
  wire s68, sub68, and68, or68;
  wire b_inv68;
  assign b_inv68 = ~b68;
  assign s68  = a68 ^ b68 ^ c68;
  assign sub68 = a68 ^ b_inv68 ^ c68;
  assign and68 = a68 & b68;
  assign or68  = a68 | b68;
  assign c69 = (a68 & b68) | (a68 & c68) | (b68 & c68);
  wire c_sub69;
  assign c_sub69 = (a68 & b_inv68) | (a68 & c68) | (b_inv68 & c68);
  wire s69, sub69, and69, or69;
  wire b_inv69;
  assign b_inv69 = ~b69;
  assign s69  = a69 ^ b69 ^ c69;
  assign sub69 = a69 ^ b_inv69 ^ c69;
  assign and69 = a69 & b69;
  assign or69  = a69 | b69;
  assign c70 = (a69 & b69) | (a69 & c69) | (b69 & c69);
  wire c_sub70;
  assign c_sub70 = (a69 & b_inv69) | (a69 & c69) | (b_inv69 & c69);
  wire s70, sub70, and70, or70;
  wire b_inv70;
  assign b_inv70 = ~b70;
  assign s70  = a70 ^ b70 ^ c70;
  assign sub70 = a70 ^ b_inv70 ^ c70;
  assign and70 = a70 & b70;
  assign or70  = a70 | b70;
  assign c71 = (a70 & b70) | (a70 & c70) | (b70 & c70);
  wire c_sub71;
  assign c_sub71 = (a70 & b_inv70) | (a70 & c70) | (b_inv70 & c70);
  wire s71, sub71, and71, or71;
  wire b_inv71;
  assign b_inv71 = ~b71;
  assign s71  = a71 ^ b71 ^ c71;
  assign sub71 = a71 ^ b_inv71 ^ c71;
  assign and71 = a71 & b71;
  assign or71  = a71 | b71;
  assign c72 = (a71 & b71) | (a71 & c71) | (b71 & c71);
  wire c_sub72;
  assign c_sub72 = (a71 & b_inv71) | (a71 & c71) | (b_inv71 & c71);
  wire s72, sub72, and72, or72;
  wire b_inv72;
  assign b_inv72 = ~b72;
  assign s72  = a72 ^ b72 ^ c72;
  assign sub72 = a72 ^ b_inv72 ^ c72;
  assign and72 = a72 & b72;
  assign or72  = a72 | b72;
  assign c73 = (a72 & b72) | (a72 & c72) | (b72 & c72);
  wire c_sub73;
  assign c_sub73 = (a72 & b_inv72) | (a72 & c72) | (b_inv72 & c72);
  wire s73, sub73, and73, or73;
  wire b_inv73;
  assign b_inv73 = ~b73;
  assign s73  = a73 ^ b73 ^ c73;
  assign sub73 = a73 ^ b_inv73 ^ c73;
  assign and73 = a73 & b73;
  assign or73  = a73 | b73;
  assign c74 = (a73 & b73) | (a73 & c73) | (b73 & c73);
  wire c_sub74;
  assign c_sub74 = (a73 & b_inv73) | (a73 & c73) | (b_inv73 & c73);
  wire s74, sub74, and74, or74;
  wire b_inv74;
  assign b_inv74 = ~b74;
  assign s74  = a74 ^ b74 ^ c74;
  assign sub74 = a74 ^ b_inv74 ^ c74;
  assign and74 = a74 & b74;
  assign or74  = a74 | b74;
  assign c75 = (a74 & b74) | (a74 & c74) | (b74 & c74);
  wire c_sub75;
  assign c_sub75 = (a74 & b_inv74) | (a74 & c74) | (b_inv74 & c74);
  wire s75, sub75, and75, or75;
  wire b_inv75;
  assign b_inv75 = ~b75;
  assign s75  = a75 ^ b75 ^ c75;
  assign sub75 = a75 ^ b_inv75 ^ c75;
  assign and75 = a75 & b75;
  assign or75  = a75 | b75;
  assign c76 = (a75 & b75) | (a75 & c75) | (b75 & c75);
  wire c_sub76;
  assign c_sub76 = (a75 & b_inv75) | (a75 & c75) | (b_inv75 & c75);
  wire s76, sub76, and76, or76;
  wire b_inv76;
  assign b_inv76 = ~b76;
  assign s76  = a76 ^ b76 ^ c76;
  assign sub76 = a76 ^ b_inv76 ^ c76;
  assign and76 = a76 & b76;
  assign or76  = a76 | b76;
  assign c77 = (a76 & b76) | (a76 & c76) | (b76 & c76);
  wire c_sub77;
  assign c_sub77 = (a76 & b_inv76) | (a76 & c76) | (b_inv76 & c76);
  wire s77, sub77, and77, or77;
  wire b_inv77;
  assign b_inv77 = ~b77;
  assign s77  = a77 ^ b77 ^ c77;
  assign sub77 = a77 ^ b_inv77 ^ c77;
  assign and77 = a77 & b77;
  assign or77  = a77 | b77;
  assign c78 = (a77 & b77) | (a77 & c77) | (b77 & c77);
  wire c_sub78;
  assign c_sub78 = (a77 & b_inv77) | (a77 & c77) | (b_inv77 & c77);
  wire s78, sub78, and78, or78;
  wire b_inv78;
  assign b_inv78 = ~b78;
  assign s78  = a78 ^ b78 ^ c78;
  assign sub78 = a78 ^ b_inv78 ^ c78;
  assign and78 = a78 & b78;
  assign or78  = a78 | b78;
  assign c79 = (a78 & b78) | (a78 & c78) | (b78 & c78);
  wire c_sub79;
  assign c_sub79 = (a78 & b_inv78) | (a78 & c78) | (b_inv78 & c78);
  wire s79, sub79, and79, or79;
  wire b_inv79;
  assign b_inv79 = ~b79;
  assign s79  = a79 ^ b79 ^ c79;
  assign sub79 = a79 ^ b_inv79 ^ c79;
  assign and79 = a79 & b79;
  assign or79  = a79 | b79;
  assign c80 = (a79 & b79) | (a79 & c79) | (b79 & c79);
  wire c_sub80;
  assign c_sub80 = (a79 & b_inv79) | (a79 & c79) | (b_inv79 & c79);
  wire s80, sub80, and80, or80;
  wire b_inv80;
  assign b_inv80 = ~b80;
  assign s80  = a80 ^ b80 ^ c80;
  assign sub80 = a80 ^ b_inv80 ^ c80;
  assign and80 = a80 & b80;
  assign or80  = a80 | b80;
  assign c81 = (a80 & b80) | (a80 & c80) | (b80 & c80);
  wire c_sub81;
  assign c_sub81 = (a80 & b_inv80) | (a80 & c80) | (b_inv80 & c80);
  wire s81, sub81, and81, or81;
  wire b_inv81;
  assign b_inv81 = ~b81;
  assign s81  = a81 ^ b81 ^ c81;
  assign sub81 = a81 ^ b_inv81 ^ c81;
  assign and81 = a81 & b81;
  assign or81  = a81 | b81;
  assign c82 = (a81 & b81) | (a81 & c81) | (b81 & c81);
  wire c_sub82;
  assign c_sub82 = (a81 & b_inv81) | (a81 & c81) | (b_inv81 & c81);
  wire s82, sub82, and82, or82;
  wire b_inv82;
  assign b_inv82 = ~b82;
  assign s82  = a82 ^ b82 ^ c82;
  assign sub82 = a82 ^ b_inv82 ^ c82;
  assign and82 = a82 & b82;
  assign or82  = a82 | b82;
  assign c83 = (a82 & b82) | (a82 & c82) | (b82 & c82);
  wire c_sub83;
  assign c_sub83 = (a82 & b_inv82) | (a82 & c82) | (b_inv82 & c82);
  wire s83, sub83, and83, or83;
  wire b_inv83;
  assign b_inv83 = ~b83;
  assign s83  = a83 ^ b83 ^ c83;
  assign sub83 = a83 ^ b_inv83 ^ c83;
  assign and83 = a83 & b83;
  assign or83  = a83 | b83;
  assign c84 = (a83 & b83) | (a83 & c83) | (b83 & c83);
  wire c_sub84;
  assign c_sub84 = (a83 & b_inv83) | (a83 & c83) | (b_inv83 & c83);
  wire s84, sub84, and84, or84;
  wire b_inv84;
  assign b_inv84 = ~b84;
  assign s84  = a84 ^ b84 ^ c84;
  assign sub84 = a84 ^ b_inv84 ^ c84;
  assign and84 = a84 & b84;
  assign or84  = a84 | b84;
  assign c85 = (a84 & b84) | (a84 & c84) | (b84 & c84);
  wire c_sub85;
  assign c_sub85 = (a84 & b_inv84) | (a84 & c84) | (b_inv84 & c84);
  wire s85, sub85, and85, or85;
  wire b_inv85;
  assign b_inv85 = ~b85;
  assign s85  = a85 ^ b85 ^ c85;
  assign sub85 = a85 ^ b_inv85 ^ c85;
  assign and85 = a85 & b85;
  assign or85  = a85 | b85;
  assign c86 = (a85 & b85) | (a85 & c85) | (b85 & c85);
  wire c_sub86;
  assign c_sub86 = (a85 & b_inv85) | (a85 & c85) | (b_inv85 & c85);
  wire s86, sub86, and86, or86;
  wire b_inv86;
  assign b_inv86 = ~b86;
  assign s86  = a86 ^ b86 ^ c86;
  assign sub86 = a86 ^ b_inv86 ^ c86;
  assign and86 = a86 & b86;
  assign or86  = a86 | b86;
  assign c87 = (a86 & b86) | (a86 & c86) | (b86 & c86);
  wire c_sub87;
  assign c_sub87 = (a86 & b_inv86) | (a86 & c86) | (b_inv86 & c86);
  wire s87, sub87, and87, or87;
  wire b_inv87;
  assign b_inv87 = ~b87;
  assign s87  = a87 ^ b87 ^ c87;
  assign sub87 = a87 ^ b_inv87 ^ c87;
  assign and87 = a87 & b87;
  assign or87  = a87 | b87;
  assign c88 = (a87 & b87) | (a87 & c87) | (b87 & c87);
  wire c_sub88;
  assign c_sub88 = (a87 & b_inv87) | (a87 & c87) | (b_inv87 & c87);
  wire s88, sub88, and88, or88;
  wire b_inv88;
  assign b_inv88 = ~b88;
  assign s88  = a88 ^ b88 ^ c88;
  assign sub88 = a88 ^ b_inv88 ^ c88;
  assign and88 = a88 & b88;
  assign or88  = a88 | b88;
  assign c89 = (a88 & b88) | (a88 & c88) | (b88 & c88);
  wire c_sub89;
  assign c_sub89 = (a88 & b_inv88) | (a88 & c88) | (b_inv88 & c88);
  wire s89, sub89, and89, or89;
  wire b_inv89;
  assign b_inv89 = ~b89;
  assign s89  = a89 ^ b89 ^ c89;
  assign sub89 = a89 ^ b_inv89 ^ c89;
  assign and89 = a89 & b89;
  assign or89  = a89 | b89;
  assign c90 = (a89 & b89) | (a89 & c89) | (b89 & c89);
  wire c_sub90;
  assign c_sub90 = (a89 & b_inv89) | (a89 & c89) | (b_inv89 & c89);
  wire s90, sub90, and90, or90;
  wire b_inv90;
  assign b_inv90 = ~b90;
  assign s90  = a90 ^ b90 ^ c90;
  assign sub90 = a90 ^ b_inv90 ^ c90;
  assign and90 = a90 & b90;
  assign or90  = a90 | b90;
  assign c91 = (a90 & b90) | (a90 & c90) | (b90 & c90);
  wire c_sub91;
  assign c_sub91 = (a90 & b_inv90) | (a90 & c90) | (b_inv90 & c90);
  wire s91, sub91, and91, or91;
  wire b_inv91;
  assign b_inv91 = ~b91;
  assign s91  = a91 ^ b91 ^ c91;
  assign sub91 = a91 ^ b_inv91 ^ c91;
  assign and91 = a91 & b91;
  assign or91  = a91 | b91;
  assign c92 = (a91 & b91) | (a91 & c91) | (b91 & c91);
  wire c_sub92;
  assign c_sub92 = (a91 & b_inv91) | (a91 & c91) | (b_inv91 & c91);
  wire s92, sub92, and92, or92;
  wire b_inv92;
  assign b_inv92 = ~b92;
  assign s92  = a92 ^ b92 ^ c92;
  assign sub92 = a92 ^ b_inv92 ^ c92;
  assign and92 = a92 & b92;
  assign or92  = a92 | b92;
  assign c93 = (a92 & b92) | (a92 & c92) | (b92 & c92);
  wire c_sub93;
  assign c_sub93 = (a92 & b_inv92) | (a92 & c92) | (b_inv92 & c92);
  wire s93, sub93, and93, or93;
  wire b_inv93;
  assign b_inv93 = ~b93;
  assign s93  = a93 ^ b93 ^ c93;
  assign sub93 = a93 ^ b_inv93 ^ c93;
  assign and93 = a93 & b93;
  assign or93  = a93 | b93;
  assign c94 = (a93 & b93) | (a93 & c93) | (b93 & c93);
  wire c_sub94;
  assign c_sub94 = (a93 & b_inv93) | (a93 & c93) | (b_inv93 & c93);
  wire s94, sub94, and94, or94;
  wire b_inv94;
  assign b_inv94 = ~b94;
  assign s94  = a94 ^ b94 ^ c94;
  assign sub94 = a94 ^ b_inv94 ^ c94;
  assign and94 = a94 & b94;
  assign or94  = a94 | b94;
  assign c95 = (a94 & b94) | (a94 & c94) | (b94 & c94);
  wire c_sub95;
  assign c_sub95 = (a94 & b_inv94) | (a94 & c94) | (b_inv94 & c94);
  wire s95, sub95, and95, or95;
  wire b_inv95;
  assign b_inv95 = ~b95;
  assign s95  = a95 ^ b95 ^ c95;
  assign sub95 = a95 ^ b_inv95 ^ c95;
  assign and95 = a95 & b95;
  assign or95  = a95 | b95;
  assign c96 = (a95 & b95) | (a95 & c95) | (b95 & c95);
  wire c_sub96;
  assign c_sub96 = (a95 & b_inv95) | (a95 & c95) | (b_inv95 & c95);
  wire s96, sub96, and96, or96;
  wire b_inv96;
  assign b_inv96 = ~b96;
  assign s96  = a96 ^ b96 ^ c96;
  assign sub96 = a96 ^ b_inv96 ^ c96;
  assign and96 = a96 & b96;
  assign or96  = a96 | b96;
  assign c97 = (a96 & b96) | (a96 & c96) | (b96 & c96);
  wire c_sub97;
  assign c_sub97 = (a96 & b_inv96) | (a96 & c96) | (b_inv96 & c96);
  wire s97, sub97, and97, or97;
  wire b_inv97;
  assign b_inv97 = ~b97;
  assign s97  = a97 ^ b97 ^ c97;
  assign sub97 = a97 ^ b_inv97 ^ c97;
  assign and97 = a97 & b97;
  assign or97  = a97 | b97;
  assign c98 = (a97 & b97) | (a97 & c97) | (b97 & c97);
  wire c_sub98;
  assign c_sub98 = (a97 & b_inv97) | (a97 & c97) | (b_inv97 & c97);
  wire s98, sub98, and98, or98;
  wire b_inv98;
  assign b_inv98 = ~b98;
  assign s98  = a98 ^ b98 ^ c98;
  assign sub98 = a98 ^ b_inv98 ^ c98;
  assign and98 = a98 & b98;
  assign or98  = a98 | b98;
  assign c99 = (a98 & b98) | (a98 & c98) | (b98 & c98);
  wire c_sub99;
  assign c_sub99 = (a98 & b_inv98) | (a98 & c98) | (b_inv98 & c98);
  wire s99, sub99, and99, or99;
  wire b_inv99;
  assign b_inv99 = ~b99;
  assign s99  = a99 ^ b99 ^ c99;
  assign sub99 = a99 ^ b_inv99 ^ c99;
  assign and99 = a99 & b99;
  assign or99  = a99 | b99;
  assign c100 = (a99 & b99) | (a99 & c99) | (b99 & c99);
  wire c_sub100;
  assign c_sub100 = (a99 & b_inv99) | (a99 & c99) | (b_inv99 & c99);
  wire s100, sub100, and100, or100;
  wire b_inv100;
  assign b_inv100 = ~b100;
  assign s100  = a100 ^ b100 ^ c100;
  assign sub100 = a100 ^ b_inv100 ^ c100;
  assign and100 = a100 & b100;
  assign or100  = a100 | b100;
  assign c101 = (a100 & b100) | (a100 & c100) | (b100 & c100);
  wire c_sub101;
  assign c_sub101 = (a100 & b_inv100) | (a100 & c100) | (b_inv100 & c100);
  wire s101, sub101, and101, or101;
  wire b_inv101;
  assign b_inv101 = ~b101;
  assign s101  = a101 ^ b101 ^ c101;
  assign sub101 = a101 ^ b_inv101 ^ c101;
  assign and101 = a101 & b101;
  assign or101  = a101 | b101;
  assign c102 = (a101 & b101) | (a101 & c101) | (b101 & c101);
  wire c_sub102;
  assign c_sub102 = (a101 & b_inv101) | (a101 & c101) | (b_inv101 & c101);
  wire s102, sub102, and102, or102;
  wire b_inv102;
  assign b_inv102 = ~b102;
  assign s102  = a102 ^ b102 ^ c102;
  assign sub102 = a102 ^ b_inv102 ^ c102;
  assign and102 = a102 & b102;
  assign or102  = a102 | b102;
  assign c103 = (a102 & b102) | (a102 & c102) | (b102 & c102);
  wire c_sub103;
  assign c_sub103 = (a102 & b_inv102) | (a102 & c102) | (b_inv102 & c102);
  wire s103, sub103, and103, or103;
  wire b_inv103;
  assign b_inv103 = ~b103;
  assign s103  = a103 ^ b103 ^ c103;
  assign sub103 = a103 ^ b_inv103 ^ c103;
  assign and103 = a103 & b103;
  assign or103  = a103 | b103;
  assign c104 = (a103 & b103) | (a103 & c103) | (b103 & c103);
  wire c_sub104;
  assign c_sub104 = (a103 & b_inv103) | (a103 & c103) | (b_inv103 & c103);
  wire s104, sub104, and104, or104;
  wire b_inv104;
  assign b_inv104 = ~b104;
  assign s104  = a104 ^ b104 ^ c104;
  assign sub104 = a104 ^ b_inv104 ^ c104;
  assign and104 = a104 & b104;
  assign or104  = a104 | b104;
  assign c105 = (a104 & b104) | (a104 & c104) | (b104 & c104);
  wire c_sub105;
  assign c_sub105 = (a104 & b_inv104) | (a104 & c104) | (b_inv104 & c104);
  wire s105, sub105, and105, or105;
  wire b_inv105;
  assign b_inv105 = ~b105;
  assign s105  = a105 ^ b105 ^ c105;
  assign sub105 = a105 ^ b_inv105 ^ c105;
  assign and105 = a105 & b105;
  assign or105  = a105 | b105;
  assign c106 = (a105 & b105) | (a105 & c105) | (b105 & c105);
  wire c_sub106;
  assign c_sub106 = (a105 & b_inv105) | (a105 & c105) | (b_inv105 & c105);
  wire s106, sub106, and106, or106;
  wire b_inv106;
  assign b_inv106 = ~b106;
  assign s106  = a106 ^ b106 ^ c106;
  assign sub106 = a106 ^ b_inv106 ^ c106;
  assign and106 = a106 & b106;
  assign or106  = a106 | b106;
  assign c107 = (a106 & b106) | (a106 & c106) | (b106 & c106);
  wire c_sub107;
  assign c_sub107 = (a106 & b_inv106) | (a106 & c106) | (b_inv106 & c106);
  wire s107, sub107, and107, or107;
  wire b_inv107;
  assign b_inv107 = ~b107;
  assign s107  = a107 ^ b107 ^ c107;
  assign sub107 = a107 ^ b_inv107 ^ c107;
  assign and107 = a107 & b107;
  assign or107  = a107 | b107;
  assign c108 = (a107 & b107) | (a107 & c107) | (b107 & c107);
  wire c_sub108;
  assign c_sub108 = (a107 & b_inv107) | (a107 & c107) | (b_inv107 & c107);
  wire s108, sub108, and108, or108;
  wire b_inv108;
  assign b_inv108 = ~b108;
  assign s108  = a108 ^ b108 ^ c108;
  assign sub108 = a108 ^ b_inv108 ^ c108;
  assign and108 = a108 & b108;
  assign or108  = a108 | b108;
  assign c109 = (a108 & b108) | (a108 & c108) | (b108 & c108);
  wire c_sub109;
  assign c_sub109 = (a108 & b_inv108) | (a108 & c108) | (b_inv108 & c108);
  wire s109, sub109, and109, or109;
  wire b_inv109;
  assign b_inv109 = ~b109;
  assign s109  = a109 ^ b109 ^ c109;
  assign sub109 = a109 ^ b_inv109 ^ c109;
  assign and109 = a109 & b109;
  assign or109  = a109 | b109;
  assign c110 = (a109 & b109) | (a109 & c109) | (b109 & c109);
  wire c_sub110;
  assign c_sub110 = (a109 & b_inv109) | (a109 & c109) | (b_inv109 & c109);
  wire s110, sub110, and110, or110;
  wire b_inv110;
  assign b_inv110 = ~b110;
  assign s110  = a110 ^ b110 ^ c110;
  assign sub110 = a110 ^ b_inv110 ^ c110;
  assign and110 = a110 & b110;
  assign or110  = a110 | b110;
  assign c111 = (a110 & b110) | (a110 & c110) | (b110 & c110);
  wire c_sub111;
  assign c_sub111 = (a110 & b_inv110) | (a110 & c110) | (b_inv110 & c110);
  wire s111, sub111, and111, or111;
  wire b_inv111;
  assign b_inv111 = ~b111;
  assign s111  = a111 ^ b111 ^ c111;
  assign sub111 = a111 ^ b_inv111 ^ c111;
  assign and111 = a111 & b111;
  assign or111  = a111 | b111;
  assign c112 = (a111 & b111) | (a111 & c111) | (b111 & c111);
  wire c_sub112;
  assign c_sub112 = (a111 & b_inv111) | (a111 & c111) | (b_inv111 & c111);
  wire s112, sub112, and112, or112;
  wire b_inv112;
  assign b_inv112 = ~b112;
  assign s112  = a112 ^ b112 ^ c112;
  assign sub112 = a112 ^ b_inv112 ^ c112;
  assign and112 = a112 & b112;
  assign or112  = a112 | b112;
  assign c113 = (a112 & b112) | (a112 & c112) | (b112 & c112);
  wire c_sub113;
  assign c_sub113 = (a112 & b_inv112) | (a112 & c112) | (b_inv112 & c112);
  wire s113, sub113, and113, or113;
  wire b_inv113;
  assign b_inv113 = ~b113;
  assign s113  = a113 ^ b113 ^ c113;
  assign sub113 = a113 ^ b_inv113 ^ c113;
  assign and113 = a113 & b113;
  assign or113  = a113 | b113;
  assign c114 = (a113 & b113) | (a113 & c113) | (b113 & c113);
  wire c_sub114;
  assign c_sub114 = (a113 & b_inv113) | (a113 & c113) | (b_inv113 & c113);
  wire s114, sub114, and114, or114;
  wire b_inv114;
  assign b_inv114 = ~b114;
  assign s114  = a114 ^ b114 ^ c114;
  assign sub114 = a114 ^ b_inv114 ^ c114;
  assign and114 = a114 & b114;
  assign or114  = a114 | b114;
  assign c115 = (a114 & b114) | (a114 & c114) | (b114 & c114);
  wire c_sub115;
  assign c_sub115 = (a114 & b_inv114) | (a114 & c114) | (b_inv114 & c114);
  wire s115, sub115, and115, or115;
  wire b_inv115;
  assign b_inv115 = ~b115;
  assign s115  = a115 ^ b115 ^ c115;
  assign sub115 = a115 ^ b_inv115 ^ c115;
  assign and115 = a115 & b115;
  assign or115  = a115 | b115;
  assign c116 = (a115 & b115) | (a115 & c115) | (b115 & c115);
  wire c_sub116;
  assign c_sub116 = (a115 & b_inv115) | (a115 & c115) | (b_inv115 & c115);
  wire s116, sub116, and116, or116;
  wire b_inv116;
  assign b_inv116 = ~b116;
  assign s116  = a116 ^ b116 ^ c116;
  assign sub116 = a116 ^ b_inv116 ^ c116;
  assign and116 = a116 & b116;
  assign or116  = a116 | b116;
  assign c117 = (a116 & b116) | (a116 & c116) | (b116 & c116);
  wire c_sub117;
  assign c_sub117 = (a116 & b_inv116) | (a116 & c116) | (b_inv116 & c116);
  wire s117, sub117, and117, or117;
  wire b_inv117;
  assign b_inv117 = ~b117;
  assign s117  = a117 ^ b117 ^ c117;
  assign sub117 = a117 ^ b_inv117 ^ c117;
  assign and117 = a117 & b117;
  assign or117  = a117 | b117;
  assign c118 = (a117 & b117) | (a117 & c117) | (b117 & c117);
  wire c_sub118;
  assign c_sub118 = (a117 & b_inv117) | (a117 & c117) | (b_inv117 & c117);
  wire s118, sub118, and118, or118;
  wire b_inv118;
  assign b_inv118 = ~b118;
  assign s118  = a118 ^ b118 ^ c118;
  assign sub118 = a118 ^ b_inv118 ^ c118;
  assign and118 = a118 & b118;
  assign or118  = a118 | b118;
  assign c119 = (a118 & b118) | (a118 & c118) | (b118 & c118);
  wire c_sub119;
  assign c_sub119 = (a118 & b_inv118) | (a118 & c118) | (b_inv118 & c118);
  wire s119, sub119, and119, or119;
  wire b_inv119;
  assign b_inv119 = ~b119;
  assign s119  = a119 ^ b119 ^ c119;
  assign sub119 = a119 ^ b_inv119 ^ c119;
  assign and119 = a119 & b119;
  assign or119  = a119 | b119;
  assign c120 = (a119 & b119) | (a119 & c119) | (b119 & c119);
  wire c_sub120;
  assign c_sub120 = (a119 & b_inv119) | (a119 & c119) | (b_inv119 & c119);
  wire s120, sub120, and120, or120;
  wire b_inv120;
  assign b_inv120 = ~b120;
  assign s120  = a120 ^ b120 ^ c120;
  assign sub120 = a120 ^ b_inv120 ^ c120;
  assign and120 = a120 & b120;
  assign or120  = a120 | b120;
  assign c121 = (a120 & b120) | (a120 & c120) | (b120 & c120);
  wire c_sub121;
  assign c_sub121 = (a120 & b_inv120) | (a120 & c120) | (b_inv120 & c120);
  wire s121, sub121, and121, or121;
  wire b_inv121;
  assign b_inv121 = ~b121;
  assign s121  = a121 ^ b121 ^ c121;
  assign sub121 = a121 ^ b_inv121 ^ c121;
  assign and121 = a121 & b121;
  assign or121  = a121 | b121;
  assign c122 = (a121 & b121) | (a121 & c121) | (b121 & c121);
  wire c_sub122;
  assign c_sub122 = (a121 & b_inv121) | (a121 & c121) | (b_inv121 & c121);
  wire s122, sub122, and122, or122;
  wire b_inv122;
  assign b_inv122 = ~b122;
  assign s122  = a122 ^ b122 ^ c122;
  assign sub122 = a122 ^ b_inv122 ^ c122;
  assign and122 = a122 & b122;
  assign or122  = a122 | b122;
  assign c123 = (a122 & b122) | (a122 & c122) | (b122 & c122);
  wire c_sub123;
  assign c_sub123 = (a122 & b_inv122) | (a122 & c122) | (b_inv122 & c122);
  wire s123, sub123, and123, or123;
  wire b_inv123;
  assign b_inv123 = ~b123;
  assign s123  = a123 ^ b123 ^ c123;
  assign sub123 = a123 ^ b_inv123 ^ c123;
  assign and123 = a123 & b123;
  assign or123  = a123 | b123;
  assign c124 = (a123 & b123) | (a123 & c123) | (b123 & c123);
  wire c_sub124;
  assign c_sub124 = (a123 & b_inv123) | (a123 & c123) | (b_inv123 & c123);
  wire s124, sub124, and124, or124;
  wire b_inv124;
  assign b_inv124 = ~b124;
  assign s124  = a124 ^ b124 ^ c124;
  assign sub124 = a124 ^ b_inv124 ^ c124;
  assign and124 = a124 & b124;
  assign or124  = a124 | b124;
  assign c125 = (a124 & b124) | (a124 & c124) | (b124 & c124);
  wire c_sub125;
  assign c_sub125 = (a124 & b_inv124) | (a124 & c124) | (b_inv124 & c124);
  wire s125, sub125, and125, or125;
  wire b_inv125;
  assign b_inv125 = ~b125;
  assign s125  = a125 ^ b125 ^ c125;
  assign sub125 = a125 ^ b_inv125 ^ c125;
  assign and125 = a125 & b125;
  assign or125  = a125 | b125;
  assign c126 = (a125 & b125) | (a125 & c125) | (b125 & c125);
  wire c_sub126;
  assign c_sub126 = (a125 & b_inv125) | (a125 & c125) | (b_inv125 & c125);
  wire s126, sub126, and126, or126;
  wire b_inv126;
  assign b_inv126 = ~b126;
  assign s126  = a126 ^ b126 ^ c126;
  assign sub126 = a126 ^ b_inv126 ^ c126;
  assign and126 = a126 & b126;
  assign or126  = a126 | b126;
  assign c127 = (a126 & b126) | (a126 & c126) | (b126 & c126);
  wire c_sub127;
  assign c_sub127 = (a126 & b_inv126) | (a126 & c126) | (b_inv126 & c126);
  wire s127, sub127, and127, or127;
  wire b_inv127;
  assign b_inv127 = ~b127;
  assign s127  = a127 ^ b127 ^ c127;
  assign sub127 = a127 ^ b_inv127 ^ c127;
  assign and127 = a127 & b127;
  assign or127  = a127 | b127;
  assign c128 = (a127 & b127) | (a127 & c127) | (b127 & c127);
  wire c_sub128;
  assign c_sub128 = (a127 & b_inv127) | (a127 & c127) | (b_inv127 & c127);
  wire s128, sub128, and128, or128;
  wire b_inv128;
  assign b_inv128 = ~b128;
  assign s128  = a128 ^ b128 ^ c128;
  assign sub128 = a128 ^ b_inv128 ^ c128;
  assign and128 = a128 & b128;
  assign or128  = a128 | b128;
  assign c129 = (a128 & b128) | (a128 & c128) | (b128 & c128);
  wire c_sub129;
  assign c_sub129 = (a128 & b_inv128) | (a128 & c128) | (b_inv128 & c128);
  wire s129, sub129, and129, or129;
  wire b_inv129;
  assign b_inv129 = ~b129;
  assign s129  = a129 ^ b129 ^ c129;
  assign sub129 = a129 ^ b_inv129 ^ c129;
  assign and129 = a129 & b129;
  assign or129  = a129 | b129;
  assign c130 = (a129 & b129) | (a129 & c129) | (b129 & c129);
  wire c_sub130;
  assign c_sub130 = (a129 & b_inv129) | (a129 & c129) | (b_inv129 & c129);
  wire s130, sub130, and130, or130;
  wire b_inv130;
  assign b_inv130 = ~b130;
  assign s130  = a130 ^ b130 ^ c130;
  assign sub130 = a130 ^ b_inv130 ^ c130;
  assign and130 = a130 & b130;
  assign or130  = a130 | b130;
  assign c131 = (a130 & b130) | (a130 & c130) | (b130 & c130);
  wire c_sub131;
  assign c_sub131 = (a130 & b_inv130) | (a130 & c130) | (b_inv130 & c130);
  wire s131, sub131, and131, or131;
  wire b_inv131;
  assign b_inv131 = ~b131;
  assign s131  = a131 ^ b131 ^ c131;
  assign sub131 = a131 ^ b_inv131 ^ c131;
  assign and131 = a131 & b131;
  assign or131  = a131 | b131;
  assign c132 = (a131 & b131) | (a131 & c131) | (b131 & c131);
  wire c_sub132;
  assign c_sub132 = (a131 & b_inv131) | (a131 & c131) | (b_inv131 & c131);
  wire s132, sub132, and132, or132;
  wire b_inv132;
  assign b_inv132 = ~b132;
  assign s132  = a132 ^ b132 ^ c132;
  assign sub132 = a132 ^ b_inv132 ^ c132;
  assign and132 = a132 & b132;
  assign or132  = a132 | b132;
  assign c133 = (a132 & b132) | (a132 & c132) | (b132 & c132);
  wire c_sub133;
  assign c_sub133 = (a132 & b_inv132) | (a132 & c132) | (b_inv132 & c132);
  wire s133, sub133, and133, or133;
  wire b_inv133;
  assign b_inv133 = ~b133;
  assign s133  = a133 ^ b133 ^ c133;
  assign sub133 = a133 ^ b_inv133 ^ c133;
  assign and133 = a133 & b133;
  assign or133  = a133 | b133;
  assign c134 = (a133 & b133) | (a133 & c133) | (b133 & c133);
  wire c_sub134;
  assign c_sub134 = (a133 & b_inv133) | (a133 & c133) | (b_inv133 & c133);
  wire s134, sub134, and134, or134;
  wire b_inv134;
  assign b_inv134 = ~b134;
  assign s134  = a134 ^ b134 ^ c134;
  assign sub134 = a134 ^ b_inv134 ^ c134;
  assign and134 = a134 & b134;
  assign or134  = a134 | b134;
  assign c135 = (a134 & b134) | (a134 & c134) | (b134 & c134);
  wire c_sub135;
  assign c_sub135 = (a134 & b_inv134) | (a134 & c134) | (b_inv134 & c134);
  wire s135, sub135, and135, or135;
  wire b_inv135;
  assign b_inv135 = ~b135;
  assign s135  = a135 ^ b135 ^ c135;
  assign sub135 = a135 ^ b_inv135 ^ c135;
  assign and135 = a135 & b135;
  assign or135  = a135 | b135;
  assign c136 = (a135 & b135) | (a135 & c135) | (b135 & c135);
  wire c_sub136;
  assign c_sub136 = (a135 & b_inv135) | (a135 & c135) | (b_inv135 & c135);
  wire s136, sub136, and136, or136;
  wire b_inv136;
  assign b_inv136 = ~b136;
  assign s136  = a136 ^ b136 ^ c136;
  assign sub136 = a136 ^ b_inv136 ^ c136;
  assign and136 = a136 & b136;
  assign or136  = a136 | b136;
  assign c137 = (a136 & b136) | (a136 & c136) | (b136 & c136);
  wire c_sub137;
  assign c_sub137 = (a136 & b_inv136) | (a136 & c136) | (b_inv136 & c136);
  wire s137, sub137, and137, or137;
  wire b_inv137;
  assign b_inv137 = ~b137;
  assign s137  = a137 ^ b137 ^ c137;
  assign sub137 = a137 ^ b_inv137 ^ c137;
  assign and137 = a137 & b137;
  assign or137  = a137 | b137;
  assign c138 = (a137 & b137) | (a137 & c137) | (b137 & c137);
  wire c_sub138;
  assign c_sub138 = (a137 & b_inv137) | (a137 & c137) | (b_inv137 & c137);
  wire s138, sub138, and138, or138;
  wire b_inv138;
  assign b_inv138 = ~b138;
  assign s138  = a138 ^ b138 ^ c138;
  assign sub138 = a138 ^ b_inv138 ^ c138;
  assign and138 = a138 & b138;
  assign or138  = a138 | b138;
  assign c139 = (a138 & b138) | (a138 & c138) | (b138 & c138);
  wire c_sub139;
  assign c_sub139 = (a138 & b_inv138) | (a138 & c138) | (b_inv138 & c138);
  wire s139, sub139, and139, or139;
  wire b_inv139;
  assign b_inv139 = ~b139;
  assign s139  = a139 ^ b139 ^ c139;
  assign sub139 = a139 ^ b_inv139 ^ c139;
  assign and139 = a139 & b139;
  assign or139  = a139 | b139;
  assign c140 = (a139 & b139) | (a139 & c139) | (b139 & c139);
  wire c_sub140;
  assign c_sub140 = (a139 & b_inv139) | (a139 & c139) | (b_inv139 & c139);
  wire s140, sub140, and140, or140;
  wire b_inv140;
  assign b_inv140 = ~b140;
  assign s140  = a140 ^ b140 ^ c140;
  assign sub140 = a140 ^ b_inv140 ^ c140;
  assign and140 = a140 & b140;
  assign or140  = a140 | b140;
  assign c141 = (a140 & b140) | (a140 & c140) | (b140 & c140);
  wire c_sub141;
  assign c_sub141 = (a140 & b_inv140) | (a140 & c140) | (b_inv140 & c140);
  wire s141, sub141, and141, or141;
  wire b_inv141;
  assign b_inv141 = ~b141;
  assign s141  = a141 ^ b141 ^ c141;
  assign sub141 = a141 ^ b_inv141 ^ c141;
  assign and141 = a141 & b141;
  assign or141  = a141 | b141;
  assign c142 = (a141 & b141) | (a141 & c141) | (b141 & c141);
  wire c_sub142;
  assign c_sub142 = (a141 & b_inv141) | (a141 & c141) | (b_inv141 & c141);
  wire s142, sub142, and142, or142;
  wire b_inv142;
  assign b_inv142 = ~b142;
  assign s142  = a142 ^ b142 ^ c142;
  assign sub142 = a142 ^ b_inv142 ^ c142;
  assign and142 = a142 & b142;
  assign or142  = a142 | b142;
  assign c143 = (a142 & b142) | (a142 & c142) | (b142 & c142);
  wire c_sub143;
  assign c_sub143 = (a142 & b_inv142) | (a142 & c142) | (b_inv142 & c142);
  wire s143, sub143, and143, or143;
  wire b_inv143;
  assign b_inv143 = ~b143;
  assign s143  = a143 ^ b143 ^ c143;
  assign sub143 = a143 ^ b_inv143 ^ c143;
  assign and143 = a143 & b143;
  assign or143  = a143 | b143;
  assign c144 = (a143 & b143) | (a143 & c143) | (b143 & c143);
  wire c_sub144;
  assign c_sub144 = (a143 & b_inv143) | (a143 & c143) | (b_inv143 & c143);
  wire s144, sub144, and144, or144;
  wire b_inv144;
  assign b_inv144 = ~b144;
  assign s144  = a144 ^ b144 ^ c144;
  assign sub144 = a144 ^ b_inv144 ^ c144;
  assign and144 = a144 & b144;
  assign or144  = a144 | b144;
  assign c145 = (a144 & b144) | (a144 & c144) | (b144 & c144);
  wire c_sub145;
  assign c_sub145 = (a144 & b_inv144) | (a144 & c144) | (b_inv144 & c144);
  wire s145, sub145, and145, or145;
  wire b_inv145;
  assign b_inv145 = ~b145;
  assign s145  = a145 ^ b145 ^ c145;
  assign sub145 = a145 ^ b_inv145 ^ c145;
  assign and145 = a145 & b145;
  assign or145  = a145 | b145;
  assign c146 = (a145 & b145) | (a145 & c145) | (b145 & c145);
  wire c_sub146;
  assign c_sub146 = (a145 & b_inv145) | (a145 & c145) | (b_inv145 & c145);
  wire s146, sub146, and146, or146;
  wire b_inv146;
  assign b_inv146 = ~b146;
  assign s146  = a146 ^ b146 ^ c146;
  assign sub146 = a146 ^ b_inv146 ^ c146;
  assign and146 = a146 & b146;
  assign or146  = a146 | b146;
  assign c147 = (a146 & b146) | (a146 & c146) | (b146 & c146);
  wire c_sub147;
  assign c_sub147 = (a146 & b_inv146) | (a146 & c146) | (b_inv146 & c146);
  wire s147, sub147, and147, or147;
  wire b_inv147;
  assign b_inv147 = ~b147;
  assign s147  = a147 ^ b147 ^ c147;
  assign sub147 = a147 ^ b_inv147 ^ c147;
  assign and147 = a147 & b147;
  assign or147  = a147 | b147;
  assign c148 = (a147 & b147) | (a147 & c147) | (b147 & c147);
  wire c_sub148;
  assign c_sub148 = (a147 & b_inv147) | (a147 & c147) | (b_inv147 & c147);
  wire s148, sub148, and148, or148;
  wire b_inv148;
  assign b_inv148 = ~b148;
  assign s148  = a148 ^ b148 ^ c148;
  assign sub148 = a148 ^ b_inv148 ^ c148;
  assign and148 = a148 & b148;
  assign or148  = a148 | b148;
  assign c149 = (a148 & b148) | (a148 & c148) | (b148 & c148);
  wire c_sub149;
  assign c_sub149 = (a148 & b_inv148) | (a148 & c148) | (b_inv148 & c148);
  wire s149, sub149, and149, or149;
  wire b_inv149;
  assign b_inv149 = ~b149;
  assign s149  = a149 ^ b149 ^ c149;
  assign sub149 = a149 ^ b_inv149 ^ c149;
  assign and149 = a149 & b149;
  assign or149  = a149 | b149;
  assign c150 = (a149 & b149) | (a149 & c149) | (b149 & c149);
  wire c_sub150;
  assign c_sub150 = (a149 & b_inv149) | (a149 & c149) | (b_inv149 & c149);
  wire s150, sub150, and150, or150;
  wire b_inv150;
  assign b_inv150 = ~b150;
  assign s150  = a150 ^ b150 ^ c150;
  assign sub150 = a150 ^ b_inv150 ^ c150;
  assign and150 = a150 & b150;
  assign or150  = a150 | b150;
  assign c151 = (a150 & b150) | (a150 & c150) | (b150 & c150);
  wire c_sub151;
  assign c_sub151 = (a150 & b_inv150) | (a150 & c150) | (b_inv150 & c150);
  wire s151, sub151, and151, or151;
  wire b_inv151;
  assign b_inv151 = ~b151;
  assign s151  = a151 ^ b151 ^ c151;
  assign sub151 = a151 ^ b_inv151 ^ c151;
  assign and151 = a151 & b151;
  assign or151  = a151 | b151;
  assign c152 = (a151 & b151) | (a151 & c151) | (b151 & c151);
  wire c_sub152;
  assign c_sub152 = (a151 & b_inv151) | (a151 & c151) | (b_inv151 & c151);
  wire s152, sub152, and152, or152;
  wire b_inv152;
  assign b_inv152 = ~b152;
  assign s152  = a152 ^ b152 ^ c152;
  assign sub152 = a152 ^ b_inv152 ^ c152;
  assign and152 = a152 & b152;
  assign or152  = a152 | b152;
  assign c153 = (a152 & b152) | (a152 & c152) | (b152 & c152);
  wire c_sub153;
  assign c_sub153 = (a152 & b_inv152) | (a152 & c152) | (b_inv152 & c152);
  wire s153, sub153, and153, or153;
  wire b_inv153;
  assign b_inv153 = ~b153;
  assign s153  = a153 ^ b153 ^ c153;
  assign sub153 = a153 ^ b_inv153 ^ c153;
  assign and153 = a153 & b153;
  assign or153  = a153 | b153;
  assign c154 = (a153 & b153) | (a153 & c153) | (b153 & c153);
  wire c_sub154;
  assign c_sub154 = (a153 & b_inv153) | (a153 & c153) | (b_inv153 & c153);
  wire s154, sub154, and154, or154;
  wire b_inv154;
  assign b_inv154 = ~b154;
  assign s154  = a154 ^ b154 ^ c154;
  assign sub154 = a154 ^ b_inv154 ^ c154;
  assign and154 = a154 & b154;
  assign or154  = a154 | b154;
  assign c155 = (a154 & b154) | (a154 & c154) | (b154 & c154);
  wire c_sub155;
  assign c_sub155 = (a154 & b_inv154) | (a154 & c154) | (b_inv154 & c154);
  wire s155, sub155, and155, or155;
  wire b_inv155;
  assign b_inv155 = ~b155;
  assign s155  = a155 ^ b155 ^ c155;
  assign sub155 = a155 ^ b_inv155 ^ c155;
  assign and155 = a155 & b155;
  assign or155  = a155 | b155;
  assign c156 = (a155 & b155) | (a155 & c155) | (b155 & c155);
  wire c_sub156;
  assign c_sub156 = (a155 & b_inv155) | (a155 & c155) | (b_inv155 & c155);
  wire s156, sub156, and156, or156;
  wire b_inv156;
  assign b_inv156 = ~b156;
  assign s156  = a156 ^ b156 ^ c156;
  assign sub156 = a156 ^ b_inv156 ^ c156;
  assign and156 = a156 & b156;
  assign or156  = a156 | b156;
  assign c157 = (a156 & b156) | (a156 & c156) | (b156 & c156);
  wire c_sub157;
  assign c_sub157 = (a156 & b_inv156) | (a156 & c156) | (b_inv156 & c156);
  wire s157, sub157, and157, or157;
  wire b_inv157;
  assign b_inv157 = ~b157;
  assign s157  = a157 ^ b157 ^ c157;
  assign sub157 = a157 ^ b_inv157 ^ c157;
  assign and157 = a157 & b157;
  assign or157  = a157 | b157;
  assign c158 = (a157 & b157) | (a157 & c157) | (b157 & c157);
  wire c_sub158;
  assign c_sub158 = (a157 & b_inv157) | (a157 & c157) | (b_inv157 & c157);
  wire s158, sub158, and158, or158;
  wire b_inv158;
  assign b_inv158 = ~b158;
  assign s158  = a158 ^ b158 ^ c158;
  assign sub158 = a158 ^ b_inv158 ^ c158;
  assign and158 = a158 & b158;
  assign or158  = a158 | b158;
  assign c159 = (a158 & b158) | (a158 & c158) | (b158 & c158);
  wire c_sub159;
  assign c_sub159 = (a158 & b_inv158) | (a158 & c158) | (b_inv158 & c158);
  wire s159, sub159, and159, or159;
  wire b_inv159;
  assign b_inv159 = ~b159;
  assign s159  = a159 ^ b159 ^ c159;
  assign sub159 = a159 ^ b_inv159 ^ c159;
  assign and159 = a159 & b159;
  assign or159  = a159 | b159;
  assign c160 = (a159 & b159) | (a159 & c159) | (b159 & c159);
  wire c_sub160;
  assign c_sub160 = (a159 & b_inv159) | (a159 & c159) | (b_inv159 & c159);
  wire s160, sub160, and160, or160;
  wire b_inv160;
  assign b_inv160 = ~b160;
  assign s160  = a160 ^ b160 ^ c160;
  assign sub160 = a160 ^ b_inv160 ^ c160;
  assign and160 = a160 & b160;
  assign or160  = a160 | b160;
  assign c161 = (a160 & b160) | (a160 & c160) | (b160 & c160);
  wire c_sub161;
  assign c_sub161 = (a160 & b_inv160) | (a160 & c160) | (b_inv160 & c160);
  wire s161, sub161, and161, or161;
  wire b_inv161;
  assign b_inv161 = ~b161;
  assign s161  = a161 ^ b161 ^ c161;
  assign sub161 = a161 ^ b_inv161 ^ c161;
  assign and161 = a161 & b161;
  assign or161  = a161 | b161;
  assign c162 = (a161 & b161) | (a161 & c161) | (b161 & c161);
  wire c_sub162;
  assign c_sub162 = (a161 & b_inv161) | (a161 & c161) | (b_inv161 & c161);
  wire s162, sub162, and162, or162;
  wire b_inv162;
  assign b_inv162 = ~b162;
  assign s162  = a162 ^ b162 ^ c162;
  assign sub162 = a162 ^ b_inv162 ^ c162;
  assign and162 = a162 & b162;
  assign or162  = a162 | b162;
  assign c163 = (a162 & b162) | (a162 & c162) | (b162 & c162);
  wire c_sub163;
  assign c_sub163 = (a162 & b_inv162) | (a162 & c162) | (b_inv162 & c162);
  wire s163, sub163, and163, or163;
  wire b_inv163;
  assign b_inv163 = ~b163;
  assign s163  = a163 ^ b163 ^ c163;
  assign sub163 = a163 ^ b_inv163 ^ c163;
  assign and163 = a163 & b163;
  assign or163  = a163 | b163;
  assign c164 = (a163 & b163) | (a163 & c163) | (b163 & c163);
  wire c_sub164;
  assign c_sub164 = (a163 & b_inv163) | (a163 & c163) | (b_inv163 & c163);
  wire s164, sub164, and164, or164;
  wire b_inv164;
  assign b_inv164 = ~b164;
  assign s164  = a164 ^ b164 ^ c164;
  assign sub164 = a164 ^ b_inv164 ^ c164;
  assign and164 = a164 & b164;
  assign or164  = a164 | b164;
  assign c165 = (a164 & b164) | (a164 & c164) | (b164 & c164);
  wire c_sub165;
  assign c_sub165 = (a164 & b_inv164) | (a164 & c164) | (b_inv164 & c164);
  wire s165, sub165, and165, or165;
  wire b_inv165;
  assign b_inv165 = ~b165;
  assign s165  = a165 ^ b165 ^ c165;
  assign sub165 = a165 ^ b_inv165 ^ c165;
  assign and165 = a165 & b165;
  assign or165  = a165 | b165;
  assign c166 = (a165 & b165) | (a165 & c165) | (b165 & c165);
  wire c_sub166;
  assign c_sub166 = (a165 & b_inv165) | (a165 & c165) | (b_inv165 & c165);
  wire s166, sub166, and166, or166;
  wire b_inv166;
  assign b_inv166 = ~b166;
  assign s166  = a166 ^ b166 ^ c166;
  assign sub166 = a166 ^ b_inv166 ^ c166;
  assign and166 = a166 & b166;
  assign or166  = a166 | b166;
  assign c167 = (a166 & b166) | (a166 & c166) | (b166 & c166);
  wire c_sub167;
  assign c_sub167 = (a166 & b_inv166) | (a166 & c166) | (b_inv166 & c166);
  wire s167, sub167, and167, or167;
  wire b_inv167;
  assign b_inv167 = ~b167;
  assign s167  = a167 ^ b167 ^ c167;
  assign sub167 = a167 ^ b_inv167 ^ c167;
  assign and167 = a167 & b167;
  assign or167  = a167 | b167;
  assign c168 = (a167 & b167) | (a167 & c167) | (b167 & c167);
  wire c_sub168;
  assign c_sub168 = (a167 & b_inv167) | (a167 & c167) | (b_inv167 & c167);
  wire s168, sub168, and168, or168;
  wire b_inv168;
  assign b_inv168 = ~b168;
  assign s168  = a168 ^ b168 ^ c168;
  assign sub168 = a168 ^ b_inv168 ^ c168;
  assign and168 = a168 & b168;
  assign or168  = a168 | b168;
  assign c169 = (a168 & b168) | (a168 & c168) | (b168 & c168);
  wire c_sub169;
  assign c_sub169 = (a168 & b_inv168) | (a168 & c168) | (b_inv168 & c168);
  wire s169, sub169, and169, or169;
  wire b_inv169;
  assign b_inv169 = ~b169;
  assign s169  = a169 ^ b169 ^ c169;
  assign sub169 = a169 ^ b_inv169 ^ c169;
  assign and169 = a169 & b169;
  assign or169  = a169 | b169;
  assign c170 = (a169 & b169) | (a169 & c169) | (b169 & c169);
  wire c_sub170;
  assign c_sub170 = (a169 & b_inv169) | (a169 & c169) | (b_inv169 & c169);
  wire s170, sub170, and170, or170;
  wire b_inv170;
  assign b_inv170 = ~b170;
  assign s170  = a170 ^ b170 ^ c170;
  assign sub170 = a170 ^ b_inv170 ^ c170;
  assign and170 = a170 & b170;
  assign or170  = a170 | b170;
  assign c171 = (a170 & b170) | (a170 & c170) | (b170 & c170);
  wire c_sub171;
  assign c_sub171 = (a170 & b_inv170) | (a170 & c170) | (b_inv170 & c170);
  wire s171, sub171, and171, or171;
  wire b_inv171;
  assign b_inv171 = ~b171;
  assign s171  = a171 ^ b171 ^ c171;
  assign sub171 = a171 ^ b_inv171 ^ c171;
  assign and171 = a171 & b171;
  assign or171  = a171 | b171;
  assign c172 = (a171 & b171) | (a171 & c171) | (b171 & c171);
  wire c_sub172;
  assign c_sub172 = (a171 & b_inv171) | (a171 & c171) | (b_inv171 & c171);
  wire s172, sub172, and172, or172;
  wire b_inv172;
  assign b_inv172 = ~b172;
  assign s172  = a172 ^ b172 ^ c172;
  assign sub172 = a172 ^ b_inv172 ^ c172;
  assign and172 = a172 & b172;
  assign or172  = a172 | b172;
  assign c173 = (a172 & b172) | (a172 & c172) | (b172 & c172);
  wire c_sub173;
  assign c_sub173 = (a172 & b_inv172) | (a172 & c172) | (b_inv172 & c172);
  wire s173, sub173, and173, or173;
  wire b_inv173;
  assign b_inv173 = ~b173;
  assign s173  = a173 ^ b173 ^ c173;
  assign sub173 = a173 ^ b_inv173 ^ c173;
  assign and173 = a173 & b173;
  assign or173  = a173 | b173;
  assign c174 = (a173 & b173) | (a173 & c173) | (b173 & c173);
  wire c_sub174;
  assign c_sub174 = (a173 & b_inv173) | (a173 & c173) | (b_inv173 & c173);
  wire s174, sub174, and174, or174;
  wire b_inv174;
  assign b_inv174 = ~b174;
  assign s174  = a174 ^ b174 ^ c174;
  assign sub174 = a174 ^ b_inv174 ^ c174;
  assign and174 = a174 & b174;
  assign or174  = a174 | b174;
  assign c175 = (a174 & b174) | (a174 & c174) | (b174 & c174);
  wire c_sub175;
  assign c_sub175 = (a174 & b_inv174) | (a174 & c174) | (b_inv174 & c174);
  wire s175, sub175, and175, or175;
  wire b_inv175;
  assign b_inv175 = ~b175;
  assign s175  = a175 ^ b175 ^ c175;
  assign sub175 = a175 ^ b_inv175 ^ c175;
  assign and175 = a175 & b175;
  assign or175  = a175 | b175;
  assign c176 = (a175 & b175) | (a175 & c175) | (b175 & c175);
  wire c_sub176;
  assign c_sub176 = (a175 & b_inv175) | (a175 & c175) | (b_inv175 & c175);
  wire s176, sub176, and176, or176;
  wire b_inv176;
  assign b_inv176 = ~b176;
  assign s176  = a176 ^ b176 ^ c176;
  assign sub176 = a176 ^ b_inv176 ^ c176;
  assign and176 = a176 & b176;
  assign or176  = a176 | b176;
  assign c177 = (a176 & b176) | (a176 & c176) | (b176 & c176);
  wire c_sub177;
  assign c_sub177 = (a176 & b_inv176) | (a176 & c176) | (b_inv176 & c176);
  wire s177, sub177, and177, or177;
  wire b_inv177;
  assign b_inv177 = ~b177;
  assign s177  = a177 ^ b177 ^ c177;
  assign sub177 = a177 ^ b_inv177 ^ c177;
  assign and177 = a177 & b177;
  assign or177  = a177 | b177;
  assign c178 = (a177 & b177) | (a177 & c177) | (b177 & c177);
  wire c_sub178;
  assign c_sub178 = (a177 & b_inv177) | (a177 & c177) | (b_inv177 & c177);
  wire s178, sub178, and178, or178;
  wire b_inv178;
  assign b_inv178 = ~b178;
  assign s178  = a178 ^ b178 ^ c178;
  assign sub178 = a178 ^ b_inv178 ^ c178;
  assign and178 = a178 & b178;
  assign or178  = a178 | b178;
  assign c179 = (a178 & b178) | (a178 & c178) | (b178 & c178);
  wire c_sub179;
  assign c_sub179 = (a178 & b_inv178) | (a178 & c178) | (b_inv178 & c178);
  wire s179, sub179, and179, or179;
  wire b_inv179;
  assign b_inv179 = ~b179;
  assign s179  = a179 ^ b179 ^ c179;
  assign sub179 = a179 ^ b_inv179 ^ c179;
  assign and179 = a179 & b179;
  assign or179  = a179 | b179;
  assign c180 = (a179 & b179) | (a179 & c179) | (b179 & c179);
  wire c_sub180;
  assign c_sub180 = (a179 & b_inv179) | (a179 & c179) | (b_inv179 & c179);
  wire s180, sub180, and180, or180;
  wire b_inv180;
  assign b_inv180 = ~b180;
  assign s180  = a180 ^ b180 ^ c180;
  assign sub180 = a180 ^ b_inv180 ^ c180;
  assign and180 = a180 & b180;
  assign or180  = a180 | b180;
  assign c181 = (a180 & b180) | (a180 & c180) | (b180 & c180);
  wire c_sub181;
  assign c_sub181 = (a180 & b_inv180) | (a180 & c180) | (b_inv180 & c180);
  wire s181, sub181, and181, or181;
  wire b_inv181;
  assign b_inv181 = ~b181;
  assign s181  = a181 ^ b181 ^ c181;
  assign sub181 = a181 ^ b_inv181 ^ c181;
  assign and181 = a181 & b181;
  assign or181  = a181 | b181;
  assign c182 = (a181 & b181) | (a181 & c181) | (b181 & c181);
  wire c_sub182;
  assign c_sub182 = (a181 & b_inv181) | (a181 & c181) | (b_inv181 & c181);
  wire s182, sub182, and182, or182;
  wire b_inv182;
  assign b_inv182 = ~b182;
  assign s182  = a182 ^ b182 ^ c182;
  assign sub182 = a182 ^ b_inv182 ^ c182;
  assign and182 = a182 & b182;
  assign or182  = a182 | b182;
  assign c183 = (a182 & b182) | (a182 & c182) | (b182 & c182);
  wire c_sub183;
  assign c_sub183 = (a182 & b_inv182) | (a182 & c182) | (b_inv182 & c182);
  wire s183, sub183, and183, or183;
  wire b_inv183;
  assign b_inv183 = ~b183;
  assign s183  = a183 ^ b183 ^ c183;
  assign sub183 = a183 ^ b_inv183 ^ c183;
  assign and183 = a183 & b183;
  assign or183  = a183 | b183;
  assign c184 = (a183 & b183) | (a183 & c183) | (b183 & c183);
  wire c_sub184;
  assign c_sub184 = (a183 & b_inv183) | (a183 & c183) | (b_inv183 & c183);
  wire s184, sub184, and184, or184;
  wire b_inv184;
  assign b_inv184 = ~b184;
  assign s184  = a184 ^ b184 ^ c184;
  assign sub184 = a184 ^ b_inv184 ^ c184;
  assign and184 = a184 & b184;
  assign or184  = a184 | b184;
  assign c185 = (a184 & b184) | (a184 & c184) | (b184 & c184);
  wire c_sub185;
  assign c_sub185 = (a184 & b_inv184) | (a184 & c184) | (b_inv184 & c184);
  wire s185, sub185, and185, or185;
  wire b_inv185;
  assign b_inv185 = ~b185;
  assign s185  = a185 ^ b185 ^ c185;
  assign sub185 = a185 ^ b_inv185 ^ c185;
  assign and185 = a185 & b185;
  assign or185  = a185 | b185;
  assign c186 = (a185 & b185) | (a185 & c185) | (b185 & c185);
  wire c_sub186;
  assign c_sub186 = (a185 & b_inv185) | (a185 & c185) | (b_inv185 & c185);
  wire s186, sub186, and186, or186;
  wire b_inv186;
  assign b_inv186 = ~b186;
  assign s186  = a186 ^ b186 ^ c186;
  assign sub186 = a186 ^ b_inv186 ^ c186;
  assign and186 = a186 & b186;
  assign or186  = a186 | b186;
  assign c187 = (a186 & b186) | (a186 & c186) | (b186 & c186);
  wire c_sub187;
  assign c_sub187 = (a186 & b_inv186) | (a186 & c186) | (b_inv186 & c186);
  wire s187, sub187, and187, or187;
  wire b_inv187;
  assign b_inv187 = ~b187;
  assign s187  = a187 ^ b187 ^ c187;
  assign sub187 = a187 ^ b_inv187 ^ c187;
  assign and187 = a187 & b187;
  assign or187  = a187 | b187;
  assign c188 = (a187 & b187) | (a187 & c187) | (b187 & c187);
  wire c_sub188;
  assign c_sub188 = (a187 & b_inv187) | (a187 & c187) | (b_inv187 & c187);
  wire s188, sub188, and188, or188;
  wire b_inv188;
  assign b_inv188 = ~b188;
  assign s188  = a188 ^ b188 ^ c188;
  assign sub188 = a188 ^ b_inv188 ^ c188;
  assign and188 = a188 & b188;
  assign or188  = a188 | b188;
  assign c189 = (a188 & b188) | (a188 & c188) | (b188 & c188);
  wire c_sub189;
  assign c_sub189 = (a188 & b_inv188) | (a188 & c188) | (b_inv188 & c188);
  wire s189, sub189, and189, or189;
  wire b_inv189;
  assign b_inv189 = ~b189;
  assign s189  = a189 ^ b189 ^ c189;
  assign sub189 = a189 ^ b_inv189 ^ c189;
  assign and189 = a189 & b189;
  assign or189  = a189 | b189;
  assign c190 = (a189 & b189) | (a189 & c189) | (b189 & c189);
  wire c_sub190;
  assign c_sub190 = (a189 & b_inv189) | (a189 & c189) | (b_inv189 & c189);
  wire s190, sub190, and190, or190;
  wire b_inv190;
  assign b_inv190 = ~b190;
  assign s190  = a190 ^ b190 ^ c190;
  assign sub190 = a190 ^ b_inv190 ^ c190;
  assign and190 = a190 & b190;
  assign or190  = a190 | b190;
  assign c191 = (a190 & b190) | (a190 & c190) | (b190 & c190);
  wire c_sub191;
  assign c_sub191 = (a190 & b_inv190) | (a190 & c190) | (b_inv190 & c190);
  wire s191, sub191, and191, or191;
  wire b_inv191;
  assign b_inv191 = ~b191;
  assign s191  = a191 ^ b191 ^ c191;
  assign sub191 = a191 ^ b_inv191 ^ c191;
  assign and191 = a191 & b191;
  assign or191  = a191 | b191;
  assign c192 = (a191 & b191) | (a191 & c191) | (b191 & c191);
  wire c_sub192;
  assign c_sub192 = (a191 & b_inv191) | (a191 & c191) | (b_inv191 & c191);
  wire s192, sub192, and192, or192;
  wire b_inv192;
  assign b_inv192 = ~b192;
  assign s192  = a192 ^ b192 ^ c192;
  assign sub192 = a192 ^ b_inv192 ^ c192;
  assign and192 = a192 & b192;
  assign or192  = a192 | b192;
  assign c193 = (a192 & b192) | (a192 & c192) | (b192 & c192);
  wire c_sub193;
  assign c_sub193 = (a192 & b_inv192) | (a192 & c192) | (b_inv192 & c192);
  wire s193, sub193, and193, or193;
  wire b_inv193;
  assign b_inv193 = ~b193;
  assign s193  = a193 ^ b193 ^ c193;
  assign sub193 = a193 ^ b_inv193 ^ c193;
  assign and193 = a193 & b193;
  assign or193  = a193 | b193;
  assign c194 = (a193 & b193) | (a193 & c193) | (b193 & c193);
  wire c_sub194;
  assign c_sub194 = (a193 & b_inv193) | (a193 & c193) | (b_inv193 & c193);
  wire s194, sub194, and194, or194;
  wire b_inv194;
  assign b_inv194 = ~b194;
  assign s194  = a194 ^ b194 ^ c194;
  assign sub194 = a194 ^ b_inv194 ^ c194;
  assign and194 = a194 & b194;
  assign or194  = a194 | b194;
  assign c195 = (a194 & b194) | (a194 & c194) | (b194 & c194);
  wire c_sub195;
  assign c_sub195 = (a194 & b_inv194) | (a194 & c194) | (b_inv194 & c194);
  wire s195, sub195, and195, or195;
  wire b_inv195;
  assign b_inv195 = ~b195;
  assign s195  = a195 ^ b195 ^ c195;
  assign sub195 = a195 ^ b_inv195 ^ c195;
  assign and195 = a195 & b195;
  assign or195  = a195 | b195;
  assign c196 = (a195 & b195) | (a195 & c195) | (b195 & c195);
  wire c_sub196;
  assign c_sub196 = (a195 & b_inv195) | (a195 & c195) | (b_inv195 & c195);
  wire s196, sub196, and196, or196;
  wire b_inv196;
  assign b_inv196 = ~b196;
  assign s196  = a196 ^ b196 ^ c196;
  assign sub196 = a196 ^ b_inv196 ^ c196;
  assign and196 = a196 & b196;
  assign or196  = a196 | b196;
  assign c197 = (a196 & b196) | (a196 & c196) | (b196 & c196);
  wire c_sub197;
  assign c_sub197 = (a196 & b_inv196) | (a196 & c196) | (b_inv196 & c196);
  wire s197, sub197, and197, or197;
  wire b_inv197;
  assign b_inv197 = ~b197;
  assign s197  = a197 ^ b197 ^ c197;
  assign sub197 = a197 ^ b_inv197 ^ c197;
  assign and197 = a197 & b197;
  assign or197  = a197 | b197;
  assign c198 = (a197 & b197) | (a197 & c197) | (b197 & c197);
  wire c_sub198;
  assign c_sub198 = (a197 & b_inv197) | (a197 & c197) | (b_inv197 & c197);
  wire s198, sub198, and198, or198;
  wire b_inv198;
  assign b_inv198 = ~b198;
  assign s198  = a198 ^ b198 ^ c198;
  assign sub198 = a198 ^ b_inv198 ^ c198;
  assign and198 = a198 & b198;
  assign or198  = a198 | b198;
  assign c199 = (a198 & b198) | (a198 & c198) | (b198 & c198);
  wire c_sub199;
  assign c_sub199 = (a198 & b_inv198) | (a198 & c198) | (b_inv198 & c198);
  wire s199, sub199, and199, or199;
  wire b_inv199;
  assign b_inv199 = ~b199;
  assign s199  = a199 ^ b199 ^ c199;
  assign sub199 = a199 ^ b_inv199 ^ c199;
  assign and199 = a199 & b199;
  assign or199  = a199 | b199;
  assign c200 = (a199 & b199) | (a199 & c199) | (b199 & c199);
  wire c_sub200;
  assign c_sub200 = (a199 & b_inv199) | (a199 & c199) | (b_inv199 & c199);
  wire s200, sub200, and200, or200;
  wire b_inv200;
  assign b_inv200 = ~b200;
  assign s200  = a200 ^ b200 ^ c200;
  assign sub200 = a200 ^ b_inv200 ^ c200;
  assign and200 = a200 & b200;
  assign or200  = a200 | b200;
  assign c201 = (a200 & b200) | (a200 & c200) | (b200 & c200);
  wire c_sub201;
  assign c_sub201 = (a200 & b_inv200) | (a200 & c200) | (b_inv200 & c200);
  wire s201, sub201, and201, or201;
  wire b_inv201;
  assign b_inv201 = ~b201;
  assign s201  = a201 ^ b201 ^ c201;
  assign sub201 = a201 ^ b_inv201 ^ c201;
  assign and201 = a201 & b201;
  assign or201  = a201 | b201;
  assign c202 = (a201 & b201) | (a201 & c201) | (b201 & c201);
  wire c_sub202;
  assign c_sub202 = (a201 & b_inv201) | (a201 & c201) | (b_inv201 & c201);
  wire s202, sub202, and202, or202;
  wire b_inv202;
  assign b_inv202 = ~b202;
  assign s202  = a202 ^ b202 ^ c202;
  assign sub202 = a202 ^ b_inv202 ^ c202;
  assign and202 = a202 & b202;
  assign or202  = a202 | b202;
  assign c203 = (a202 & b202) | (a202 & c202) | (b202 & c202);
  wire c_sub203;
  assign c_sub203 = (a202 & b_inv202) | (a202 & c202) | (b_inv202 & c202);
  wire s203, sub203, and203, or203;
  wire b_inv203;
  assign b_inv203 = ~b203;
  assign s203  = a203 ^ b203 ^ c203;
  assign sub203 = a203 ^ b_inv203 ^ c203;
  assign and203 = a203 & b203;
  assign or203  = a203 | b203;
  assign c204 = (a203 & b203) | (a203 & c203) | (b203 & c203);
  wire c_sub204;
  assign c_sub204 = (a203 & b_inv203) | (a203 & c203) | (b_inv203 & c203);
  wire s204, sub204, and204, or204;
  wire b_inv204;
  assign b_inv204 = ~b204;
  assign s204  = a204 ^ b204 ^ c204;
  assign sub204 = a204 ^ b_inv204 ^ c204;
  assign and204 = a204 & b204;
  assign or204  = a204 | b204;
  assign c205 = (a204 & b204) | (a204 & c204) | (b204 & c204);
  wire c_sub205;
  assign c_sub205 = (a204 & b_inv204) | (a204 & c204) | (b_inv204 & c204);
  wire s205, sub205, and205, or205;
  wire b_inv205;
  assign b_inv205 = ~b205;
  assign s205  = a205 ^ b205 ^ c205;
  assign sub205 = a205 ^ b_inv205 ^ c205;
  assign and205 = a205 & b205;
  assign or205  = a205 | b205;
  assign c206 = (a205 & b205) | (a205 & c205) | (b205 & c205);
  wire c_sub206;
  assign c_sub206 = (a205 & b_inv205) | (a205 & c205) | (b_inv205 & c205);
  wire s206, sub206, and206, or206;
  wire b_inv206;
  assign b_inv206 = ~b206;
  assign s206  = a206 ^ b206 ^ c206;
  assign sub206 = a206 ^ b_inv206 ^ c206;
  assign and206 = a206 & b206;
  assign or206  = a206 | b206;
  assign c207 = (a206 & b206) | (a206 & c206) | (b206 & c206);
  wire c_sub207;
  assign c_sub207 = (a206 & b_inv206) | (a206 & c206) | (b_inv206 & c206);
  wire s207, sub207, and207, or207;
  wire b_inv207;
  assign b_inv207 = ~b207;
  assign s207  = a207 ^ b207 ^ c207;
  assign sub207 = a207 ^ b_inv207 ^ c207;
  assign and207 = a207 & b207;
  assign or207  = a207 | b207;
  assign c208 = (a207 & b207) | (a207 & c207) | (b207 & c207);
  wire c_sub208;
  assign c_sub208 = (a207 & b_inv207) | (a207 & c207) | (b_inv207 & c207);
  wire s208, sub208, and208, or208;
  wire b_inv208;
  assign b_inv208 = ~b208;
  assign s208  = a208 ^ b208 ^ c208;
  assign sub208 = a208 ^ b_inv208 ^ c208;
  assign and208 = a208 & b208;
  assign or208  = a208 | b208;
  assign c209 = (a208 & b208) | (a208 & c208) | (b208 & c208);
  wire c_sub209;
  assign c_sub209 = (a208 & b_inv208) | (a208 & c208) | (b_inv208 & c208);
  wire s209, sub209, and209, or209;
  wire b_inv209;
  assign b_inv209 = ~b209;
  assign s209  = a209 ^ b209 ^ c209;
  assign sub209 = a209 ^ b_inv209 ^ c209;
  assign and209 = a209 & b209;
  assign or209  = a209 | b209;
  assign c210 = (a209 & b209) | (a209 & c209) | (b209 & c209);
  wire c_sub210;
  assign c_sub210 = (a209 & b_inv209) | (a209 & c209) | (b_inv209 & c209);
  wire s210, sub210, and210, or210;
  wire b_inv210;
  assign b_inv210 = ~b210;
  assign s210  = a210 ^ b210 ^ c210;
  assign sub210 = a210 ^ b_inv210 ^ c210;
  assign and210 = a210 & b210;
  assign or210  = a210 | b210;
  assign c211 = (a210 & b210) | (a210 & c210) | (b210 & c210);
  wire c_sub211;
  assign c_sub211 = (a210 & b_inv210) | (a210 & c210) | (b_inv210 & c210);
  wire s211, sub211, and211, or211;
  wire b_inv211;
  assign b_inv211 = ~b211;
  assign s211  = a211 ^ b211 ^ c211;
  assign sub211 = a211 ^ b_inv211 ^ c211;
  assign and211 = a211 & b211;
  assign or211  = a211 | b211;
  assign c212 = (a211 & b211) | (a211 & c211) | (b211 & c211);
  wire c_sub212;
  assign c_sub212 = (a211 & b_inv211) | (a211 & c211) | (b_inv211 & c211);
  wire s212, sub212, and212, or212;
  wire b_inv212;
  assign b_inv212 = ~b212;
  assign s212  = a212 ^ b212 ^ c212;
  assign sub212 = a212 ^ b_inv212 ^ c212;
  assign and212 = a212 & b212;
  assign or212  = a212 | b212;
  assign c213 = (a212 & b212) | (a212 & c212) | (b212 & c212);
  wire c_sub213;
  assign c_sub213 = (a212 & b_inv212) | (a212 & c212) | (b_inv212 & c212);
  wire s213, sub213, and213, or213;
  wire b_inv213;
  assign b_inv213 = ~b213;
  assign s213  = a213 ^ b213 ^ c213;
  assign sub213 = a213 ^ b_inv213 ^ c213;
  assign and213 = a213 & b213;
  assign or213  = a213 | b213;
  assign c214 = (a213 & b213) | (a213 & c213) | (b213 & c213);
  wire c_sub214;
  assign c_sub214 = (a213 & b_inv213) | (a213 & c213) | (b_inv213 & c213);
  wire s214, sub214, and214, or214;
  wire b_inv214;
  assign b_inv214 = ~b214;
  assign s214  = a214 ^ b214 ^ c214;
  assign sub214 = a214 ^ b_inv214 ^ c214;
  assign and214 = a214 & b214;
  assign or214  = a214 | b214;
  assign c215 = (a214 & b214) | (a214 & c214) | (b214 & c214);
  wire c_sub215;
  assign c_sub215 = (a214 & b_inv214) | (a214 & c214) | (b_inv214 & c214);
  wire s215, sub215, and215, or215;
  wire b_inv215;
  assign b_inv215 = ~b215;
  assign s215  = a215 ^ b215 ^ c215;
  assign sub215 = a215 ^ b_inv215 ^ c215;
  assign and215 = a215 & b215;
  assign or215  = a215 | b215;
  assign c216 = (a215 & b215) | (a215 & c215) | (b215 & c215);
  wire c_sub216;
  assign c_sub216 = (a215 & b_inv215) | (a215 & c215) | (b_inv215 & c215);
  wire s216, sub216, and216, or216;
  wire b_inv216;
  assign b_inv216 = ~b216;
  assign s216  = a216 ^ b216 ^ c216;
  assign sub216 = a216 ^ b_inv216 ^ c216;
  assign and216 = a216 & b216;
  assign or216  = a216 | b216;
  assign c217 = (a216 & b216) | (a216 & c216) | (b216 & c216);
  wire c_sub217;
  assign c_sub217 = (a216 & b_inv216) | (a216 & c216) | (b_inv216 & c216);
  wire s217, sub217, and217, or217;
  wire b_inv217;
  assign b_inv217 = ~b217;
  assign s217  = a217 ^ b217 ^ c217;
  assign sub217 = a217 ^ b_inv217 ^ c217;
  assign and217 = a217 & b217;
  assign or217  = a217 | b217;
  assign c218 = (a217 & b217) | (a217 & c217) | (b217 & c217);
  wire c_sub218;
  assign c_sub218 = (a217 & b_inv217) | (a217 & c217) | (b_inv217 & c217);
  wire s218, sub218, and218, or218;
  wire b_inv218;
  assign b_inv218 = ~b218;
  assign s218  = a218 ^ b218 ^ c218;
  assign sub218 = a218 ^ b_inv218 ^ c218;
  assign and218 = a218 & b218;
  assign or218  = a218 | b218;
  assign c219 = (a218 & b218) | (a218 & c218) | (b218 & c218);
  wire c_sub219;
  assign c_sub219 = (a218 & b_inv218) | (a218 & c218) | (b_inv218 & c218);
  wire s219, sub219, and219, or219;
  wire b_inv219;
  assign b_inv219 = ~b219;
  assign s219  = a219 ^ b219 ^ c219;
  assign sub219 = a219 ^ b_inv219 ^ c219;
  assign and219 = a219 & b219;
  assign or219  = a219 | b219;
  assign c220 = (a219 & b219) | (a219 & c219) | (b219 & c219);
  wire c_sub220;
  assign c_sub220 = (a219 & b_inv219) | (a219 & c219) | (b_inv219 & c219);
  wire s220, sub220, and220, or220;
  wire b_inv220;
  assign b_inv220 = ~b220;
  assign s220  = a220 ^ b220 ^ c220;
  assign sub220 = a220 ^ b_inv220 ^ c220;
  assign and220 = a220 & b220;
  assign or220  = a220 | b220;
  assign c221 = (a220 & b220) | (a220 & c220) | (b220 & c220);
  wire c_sub221;
  assign c_sub221 = (a220 & b_inv220) | (a220 & c220) | (b_inv220 & c220);
  wire s221, sub221, and221, or221;
  wire b_inv221;
  assign b_inv221 = ~b221;
  assign s221  = a221 ^ b221 ^ c221;
  assign sub221 = a221 ^ b_inv221 ^ c221;
  assign and221 = a221 & b221;
  assign or221  = a221 | b221;
  assign c222 = (a221 & b221) | (a221 & c221) | (b221 & c221);
  wire c_sub222;
  assign c_sub222 = (a221 & b_inv221) | (a221 & c221) | (b_inv221 & c221);
  wire s222, sub222, and222, or222;
  wire b_inv222;
  assign b_inv222 = ~b222;
  assign s222  = a222 ^ b222 ^ c222;
  assign sub222 = a222 ^ b_inv222 ^ c222;
  assign and222 = a222 & b222;
  assign or222  = a222 | b222;
  assign c223 = (a222 & b222) | (a222 & c222) | (b222 & c222);
  wire c_sub223;
  assign c_sub223 = (a222 & b_inv222) | (a222 & c222) | (b_inv222 & c222);
  wire s223, sub223, and223, or223;
  wire b_inv223;
  assign b_inv223 = ~b223;
  assign s223  = a223 ^ b223 ^ c223;
  assign sub223 = a223 ^ b_inv223 ^ c223;
  assign and223 = a223 & b223;
  assign or223  = a223 | b223;
  assign c224 = (a223 & b223) | (a223 & c223) | (b223 & c223);
  wire c_sub224;
  assign c_sub224 = (a223 & b_inv223) | (a223 & c223) | (b_inv223 & c223);
  wire s224, sub224, and224, or224;
  wire b_inv224;
  assign b_inv224 = ~b224;
  assign s224  = a224 ^ b224 ^ c224;
  assign sub224 = a224 ^ b_inv224 ^ c224;
  assign and224 = a224 & b224;
  assign or224  = a224 | b224;
  assign c225 = (a224 & b224) | (a224 & c224) | (b224 & c224);
  wire c_sub225;
  assign c_sub225 = (a224 & b_inv224) | (a224 & c224) | (b_inv224 & c224);
  wire s225, sub225, and225, or225;
  wire b_inv225;
  assign b_inv225 = ~b225;
  assign s225  = a225 ^ b225 ^ c225;
  assign sub225 = a225 ^ b_inv225 ^ c225;
  assign and225 = a225 & b225;
  assign or225  = a225 | b225;
  assign c226 = (a225 & b225) | (a225 & c225) | (b225 & c225);
  wire c_sub226;
  assign c_sub226 = (a225 & b_inv225) | (a225 & c225) | (b_inv225 & c225);
  wire s226, sub226, and226, or226;
  wire b_inv226;
  assign b_inv226 = ~b226;
  assign s226  = a226 ^ b226 ^ c226;
  assign sub226 = a226 ^ b_inv226 ^ c226;
  assign and226 = a226 & b226;
  assign or226  = a226 | b226;
  assign c227 = (a226 & b226) | (a226 & c226) | (b226 & c226);
  wire c_sub227;
  assign c_sub227 = (a226 & b_inv226) | (a226 & c226) | (b_inv226 & c226);
  wire s227, sub227, and227, or227;
  wire b_inv227;
  assign b_inv227 = ~b227;
  assign s227  = a227 ^ b227 ^ c227;
  assign sub227 = a227 ^ b_inv227 ^ c227;
  assign and227 = a227 & b227;
  assign or227  = a227 | b227;
  assign c228 = (a227 & b227) | (a227 & c227) | (b227 & c227);
  wire c_sub228;
  assign c_sub228 = (a227 & b_inv227) | (a227 & c227) | (b_inv227 & c227);
  wire s228, sub228, and228, or228;
  wire b_inv228;
  assign b_inv228 = ~b228;
  assign s228  = a228 ^ b228 ^ c228;
  assign sub228 = a228 ^ b_inv228 ^ c228;
  assign and228 = a228 & b228;
  assign or228  = a228 | b228;
  assign c229 = (a228 & b228) | (a228 & c228) | (b228 & c228);
  wire c_sub229;
  assign c_sub229 = (a228 & b_inv228) | (a228 & c228) | (b_inv228 & c228);
  wire s229, sub229, and229, or229;
  wire b_inv229;
  assign b_inv229 = ~b229;
  assign s229  = a229 ^ b229 ^ c229;
  assign sub229 = a229 ^ b_inv229 ^ c229;
  assign and229 = a229 & b229;
  assign or229  = a229 | b229;
  assign c230 = (a229 & b229) | (a229 & c229) | (b229 & c229);
  wire c_sub230;
  assign c_sub230 = (a229 & b_inv229) | (a229 & c229) | (b_inv229 & c229);
  wire s230, sub230, and230, or230;
  wire b_inv230;
  assign b_inv230 = ~b230;
  assign s230  = a230 ^ b230 ^ c230;
  assign sub230 = a230 ^ b_inv230 ^ c230;
  assign and230 = a230 & b230;
  assign or230  = a230 | b230;
  assign c231 = (a230 & b230) | (a230 & c230) | (b230 & c230);
  wire c_sub231;
  assign c_sub231 = (a230 & b_inv230) | (a230 & c230) | (b_inv230 & c230);
  wire s231, sub231, and231, or231;
  wire b_inv231;
  assign b_inv231 = ~b231;
  assign s231  = a231 ^ b231 ^ c231;
  assign sub231 = a231 ^ b_inv231 ^ c231;
  assign and231 = a231 & b231;
  assign or231  = a231 | b231;
  assign c232 = (a231 & b231) | (a231 & c231) | (b231 & c231);
  wire c_sub232;
  assign c_sub232 = (a231 & b_inv231) | (a231 & c231) | (b_inv231 & c231);
  wire s232, sub232, and232, or232;
  wire b_inv232;
  assign b_inv232 = ~b232;
  assign s232  = a232 ^ b232 ^ c232;
  assign sub232 = a232 ^ b_inv232 ^ c232;
  assign and232 = a232 & b232;
  assign or232  = a232 | b232;
  assign c233 = (a232 & b232) | (a232 & c232) | (b232 & c232);
  wire c_sub233;
  assign c_sub233 = (a232 & b_inv232) | (a232 & c232) | (b_inv232 & c232);
  wire s233, sub233, and233, or233;
  wire b_inv233;
  assign b_inv233 = ~b233;
  assign s233  = a233 ^ b233 ^ c233;
  assign sub233 = a233 ^ b_inv233 ^ c233;
  assign and233 = a233 & b233;
  assign or233  = a233 | b233;
  assign c234 = (a233 & b233) | (a233 & c233) | (b233 & c233);
  wire c_sub234;
  assign c_sub234 = (a233 & b_inv233) | (a233 & c233) | (b_inv233 & c233);
  wire s234, sub234, and234, or234;
  wire b_inv234;
  assign b_inv234 = ~b234;
  assign s234  = a234 ^ b234 ^ c234;
  assign sub234 = a234 ^ b_inv234 ^ c234;
  assign and234 = a234 & b234;
  assign or234  = a234 | b234;
  assign c235 = (a234 & b234) | (a234 & c234) | (b234 & c234);
  wire c_sub235;
  assign c_sub235 = (a234 & b_inv234) | (a234 & c234) | (b_inv234 & c234);
  wire s235, sub235, and235, or235;
  wire b_inv235;
  assign b_inv235 = ~b235;
  assign s235  = a235 ^ b235 ^ c235;
  assign sub235 = a235 ^ b_inv235 ^ c235;
  assign and235 = a235 & b235;
  assign or235  = a235 | b235;
  assign c236 = (a235 & b235) | (a235 & c235) | (b235 & c235);
  wire c_sub236;
  assign c_sub236 = (a235 & b_inv235) | (a235 & c235) | (b_inv235 & c235);
  wire s236, sub236, and236, or236;
  wire b_inv236;
  assign b_inv236 = ~b236;
  assign s236  = a236 ^ b236 ^ c236;
  assign sub236 = a236 ^ b_inv236 ^ c236;
  assign and236 = a236 & b236;
  assign or236  = a236 | b236;
  assign c237 = (a236 & b236) | (a236 & c236) | (b236 & c236);
  wire c_sub237;
  assign c_sub237 = (a236 & b_inv236) | (a236 & c236) | (b_inv236 & c236);
  wire s237, sub237, and237, or237;
  wire b_inv237;
  assign b_inv237 = ~b237;
  assign s237  = a237 ^ b237 ^ c237;
  assign sub237 = a237 ^ b_inv237 ^ c237;
  assign and237 = a237 & b237;
  assign or237  = a237 | b237;
  assign c238 = (a237 & b237) | (a237 & c237) | (b237 & c237);
  wire c_sub238;
  assign c_sub238 = (a237 & b_inv237) | (a237 & c237) | (b_inv237 & c237);
  wire s238, sub238, and238, or238;
  wire b_inv238;
  assign b_inv238 = ~b238;
  assign s238  = a238 ^ b238 ^ c238;
  assign sub238 = a238 ^ b_inv238 ^ c238;
  assign and238 = a238 & b238;
  assign or238  = a238 | b238;
  assign c239 = (a238 & b238) | (a238 & c238) | (b238 & c238);
  wire c_sub239;
  assign c_sub239 = (a238 & b_inv238) | (a238 & c238) | (b_inv238 & c238);
  wire s239, sub239, and239, or239;
  wire b_inv239;
  assign b_inv239 = ~b239;
  assign s239  = a239 ^ b239 ^ c239;
  assign sub239 = a239 ^ b_inv239 ^ c239;
  assign and239 = a239 & b239;
  assign or239  = a239 | b239;
  assign c240 = (a239 & b239) | (a239 & c239) | (b239 & c239);
  wire c_sub240;
  assign c_sub240 = (a239 & b_inv239) | (a239 & c239) | (b_inv239 & c239);
  wire s240, sub240, and240, or240;
  wire b_inv240;
  assign b_inv240 = ~b240;
  assign s240  = a240 ^ b240 ^ c240;
  assign sub240 = a240 ^ b_inv240 ^ c240;
  assign and240 = a240 & b240;
  assign or240  = a240 | b240;
  assign c241 = (a240 & b240) | (a240 & c240) | (b240 & c240);
  wire c_sub241;
  assign c_sub241 = (a240 & b_inv240) | (a240 & c240) | (b_inv240 & c240);
  wire s241, sub241, and241, or241;
  wire b_inv241;
  assign b_inv241 = ~b241;
  assign s241  = a241 ^ b241 ^ c241;
  assign sub241 = a241 ^ b_inv241 ^ c241;
  assign and241 = a241 & b241;
  assign or241  = a241 | b241;
  assign c242 = (a241 & b241) | (a241 & c241) | (b241 & c241);
  wire c_sub242;
  assign c_sub242 = (a241 & b_inv241) | (a241 & c241) | (b_inv241 & c241);
  wire s242, sub242, and242, or242;
  wire b_inv242;
  assign b_inv242 = ~b242;
  assign s242  = a242 ^ b242 ^ c242;
  assign sub242 = a242 ^ b_inv242 ^ c242;
  assign and242 = a242 & b242;
  assign or242  = a242 | b242;
  assign c243 = (a242 & b242) | (a242 & c242) | (b242 & c242);
  wire c_sub243;
  assign c_sub243 = (a242 & b_inv242) | (a242 & c242) | (b_inv242 & c242);
  wire s243, sub243, and243, or243;
  wire b_inv243;
  assign b_inv243 = ~b243;
  assign s243  = a243 ^ b243 ^ c243;
  assign sub243 = a243 ^ b_inv243 ^ c243;
  assign and243 = a243 & b243;
  assign or243  = a243 | b243;
  assign c244 = (a243 & b243) | (a243 & c243) | (b243 & c243);
  wire c_sub244;
  assign c_sub244 = (a243 & b_inv243) | (a243 & c243) | (b_inv243 & c243);
  wire s244, sub244, and244, or244;
  wire b_inv244;
  assign b_inv244 = ~b244;
  assign s244  = a244 ^ b244 ^ c244;
  assign sub244 = a244 ^ b_inv244 ^ c244;
  assign and244 = a244 & b244;
  assign or244  = a244 | b244;
  assign c245 = (a244 & b244) | (a244 & c244) | (b244 & c244);
  wire c_sub245;
  assign c_sub245 = (a244 & b_inv244) | (a244 & c244) | (b_inv244 & c244);
  wire s245, sub245, and245, or245;
  wire b_inv245;
  assign b_inv245 = ~b245;
  assign s245  = a245 ^ b245 ^ c245;
  assign sub245 = a245 ^ b_inv245 ^ c245;
  assign and245 = a245 & b245;
  assign or245  = a245 | b245;
  assign c246 = (a245 & b245) | (a245 & c245) | (b245 & c245);
  wire c_sub246;
  assign c_sub246 = (a245 & b_inv245) | (a245 & c245) | (b_inv245 & c245);
  wire s246, sub246, and246, or246;
  wire b_inv246;
  assign b_inv246 = ~b246;
  assign s246  = a246 ^ b246 ^ c246;
  assign sub246 = a246 ^ b_inv246 ^ c246;
  assign and246 = a246 & b246;
  assign or246  = a246 | b246;
  assign c247 = (a246 & b246) | (a246 & c246) | (b246 & c246);
  wire c_sub247;
  assign c_sub247 = (a246 & b_inv246) | (a246 & c246) | (b_inv246 & c246);
  wire s247, sub247, and247, or247;
  wire b_inv247;
  assign b_inv247 = ~b247;
  assign s247  = a247 ^ b247 ^ c247;
  assign sub247 = a247 ^ b_inv247 ^ c247;
  assign and247 = a247 & b247;
  assign or247  = a247 | b247;
  assign c248 = (a247 & b247) | (a247 & c247) | (b247 & c247);
  wire c_sub248;
  assign c_sub248 = (a247 & b_inv247) | (a247 & c247) | (b_inv247 & c247);
  wire s248, sub248, and248, or248;
  wire b_inv248;
  assign b_inv248 = ~b248;
  assign s248  = a248 ^ b248 ^ c248;
  assign sub248 = a248 ^ b_inv248 ^ c248;
  assign and248 = a248 & b248;
  assign or248  = a248 | b248;
  assign c249 = (a248 & b248) | (a248 & c248) | (b248 & c248);
  wire c_sub249;
  assign c_sub249 = (a248 & b_inv248) | (a248 & c248) | (b_inv248 & c248);
  wire s249, sub249, and249, or249;
  wire b_inv249;
  assign b_inv249 = ~b249;
  assign s249  = a249 ^ b249 ^ c249;
  assign sub249 = a249 ^ b_inv249 ^ c249;
  assign and249 = a249 & b249;
  assign or249  = a249 | b249;
  assign c250 = (a249 & b249) | (a249 & c249) | (b249 & c249);
  wire c_sub250;
  assign c_sub250 = (a249 & b_inv249) | (a249 & c249) | (b_inv249 & c249);
  wire s250, sub250, and250, or250;
  wire b_inv250;
  assign b_inv250 = ~b250;
  assign s250  = a250 ^ b250 ^ c250;
  assign sub250 = a250 ^ b_inv250 ^ c250;
  assign and250 = a250 & b250;
  assign or250  = a250 | b250;
  assign c251 = (a250 & b250) | (a250 & c250) | (b250 & c250);
  wire c_sub251;
  assign c_sub251 = (a250 & b_inv250) | (a250 & c250) | (b_inv250 & c250);
  wire s251, sub251, and251, or251;
  wire b_inv251;
  assign b_inv251 = ~b251;
  assign s251  = a251 ^ b251 ^ c251;
  assign sub251 = a251 ^ b_inv251 ^ c251;
  assign and251 = a251 & b251;
  assign or251  = a251 | b251;
  assign c252 = (a251 & b251) | (a251 & c251) | (b251 & c251);
  wire c_sub252;
  assign c_sub252 = (a251 & b_inv251) | (a251 & c251) | (b_inv251 & c251);
  wire s252, sub252, and252, or252;
  wire b_inv252;
  assign b_inv252 = ~b252;
  assign s252  = a252 ^ b252 ^ c252;
  assign sub252 = a252 ^ b_inv252 ^ c252;
  assign and252 = a252 & b252;
  assign or252  = a252 | b252;
  assign c253 = (a252 & b252) | (a252 & c252) | (b252 & c252);
  wire c_sub253;
  assign c_sub253 = (a252 & b_inv252) | (a252 & c252) | (b_inv252 & c252);
  wire s253, sub253, and253, or253;
  wire b_inv253;
  assign b_inv253 = ~b253;
  assign s253  = a253 ^ b253 ^ c253;
  assign sub253 = a253 ^ b_inv253 ^ c253;
  assign and253 = a253 & b253;
  assign or253  = a253 | b253;
  assign c254 = (a253 & b253) | (a253 & c253) | (b253 & c253);
  wire c_sub254;
  assign c_sub254 = (a253 & b_inv253) | (a253 & c253) | (b_inv253 & c253);
  wire s254, sub254, and254, or254;
  wire b_inv254;
  assign b_inv254 = ~b254;
  assign s254  = a254 ^ b254 ^ c254;
  assign sub254 = a254 ^ b_inv254 ^ c254;
  assign and254 = a254 & b254;
  assign or254  = a254 | b254;
  assign c255 = (a254 & b254) | (a254 & c254) | (b254 & c254);
  wire c_sub255;
  assign c_sub255 = (a254 & b_inv254) | (a254 & c254) | (b_inv254 & c254);
  wire s255, sub255, and255, or255;
  wire b_inv255;
  assign b_inv255 = ~b255;
  assign s255  = a255 ^ b255 ^ c255;
  assign sub255 = a255 ^ b_inv255 ^ c255;
  assign and255 = a255 & b255;
  assign or255  = a255 | b255;
  assign c256 = (a255 & b255) | (a255 & c255) | (b255 & c255);
  wire c_sub256;
  assign c_sub256 = (a255 & b_inv255) | (a255 & c255) | (b_inv255 & c255);
  wire s256, sub256, and256, or256;
  wire b_inv256;
  assign b_inv256 = ~b256;
  assign s256  = a256 ^ b256 ^ c256;
  assign sub256 = a256 ^ b_inv256 ^ c256;
  assign and256 = a256 & b256;
  assign or256  = a256 | b256;
  assign c257 = (a256 & b256) | (a256 & c256) | (b256 & c256);
  wire c_sub257;
  assign c_sub257 = (a256 & b_inv256) | (a256 & c256) | (b_inv256 & c256);
  wire s257, sub257, and257, or257;
  wire b_inv257;
  assign b_inv257 = ~b257;
  assign s257  = a257 ^ b257 ^ c257;
  assign sub257 = a257 ^ b_inv257 ^ c257;
  assign and257 = a257 & b257;
  assign or257  = a257 | b257;
  assign c258 = (a257 & b257) | (a257 & c257) | (b257 & c257);
  wire c_sub258;
  assign c_sub258 = (a257 & b_inv257) | (a257 & c257) | (b_inv257 & c257);
  wire s258, sub258, and258, or258;
  wire b_inv258;
  assign b_inv258 = ~b258;
  assign s258  = a258 ^ b258 ^ c258;
  assign sub258 = a258 ^ b_inv258 ^ c258;
  assign and258 = a258 & b258;
  assign or258  = a258 | b258;
  assign c259 = (a258 & b258) | (a258 & c258) | (b258 & c258);
  wire c_sub259;
  assign c_sub259 = (a258 & b_inv258) | (a258 & c258) | (b_inv258 & c258);
  wire s259, sub259, and259, or259;
  wire b_inv259;
  assign b_inv259 = ~b259;
  assign s259  = a259 ^ b259 ^ c259;
  assign sub259 = a259 ^ b_inv259 ^ c259;
  assign and259 = a259 & b259;
  assign or259  = a259 | b259;
  assign c260 = (a259 & b259) | (a259 & c259) | (b259 & c259);
  wire c_sub260;
  assign c_sub260 = (a259 & b_inv259) | (a259 & c259) | (b_inv259 & c259);
  wire s260, sub260, and260, or260;
  wire b_inv260;
  assign b_inv260 = ~b260;
  assign s260  = a260 ^ b260 ^ c260;
  assign sub260 = a260 ^ b_inv260 ^ c260;
  assign and260 = a260 & b260;
  assign or260  = a260 | b260;
  assign c261 = (a260 & b260) | (a260 & c260) | (b260 & c260);
  wire c_sub261;
  assign c_sub261 = (a260 & b_inv260) | (a260 & c260) | (b_inv260 & c260);
  wire s261, sub261, and261, or261;
  wire b_inv261;
  assign b_inv261 = ~b261;
  assign s261  = a261 ^ b261 ^ c261;
  assign sub261 = a261 ^ b_inv261 ^ c261;
  assign and261 = a261 & b261;
  assign or261  = a261 | b261;
  assign c262 = (a261 & b261) | (a261 & c261) | (b261 & c261);
  wire c_sub262;
  assign c_sub262 = (a261 & b_inv261) | (a261 & c261) | (b_inv261 & c261);
  wire s262, sub262, and262, or262;
  wire b_inv262;
  assign b_inv262 = ~b262;
  assign s262  = a262 ^ b262 ^ c262;
  assign sub262 = a262 ^ b_inv262 ^ c262;
  assign and262 = a262 & b262;
  assign or262  = a262 | b262;
  assign c263 = (a262 & b262) | (a262 & c262) | (b262 & c262);
  wire c_sub263;
  assign c_sub263 = (a262 & b_inv262) | (a262 & c262) | (b_inv262 & c262);
  wire s263, sub263, and263, or263;
  wire b_inv263;
  assign b_inv263 = ~b263;
  assign s263  = a263 ^ b263 ^ c263;
  assign sub263 = a263 ^ b_inv263 ^ c263;
  assign and263 = a263 & b263;
  assign or263  = a263 | b263;
  assign c264 = (a263 & b263) | (a263 & c263) | (b263 & c263);
  wire c_sub264;
  assign c_sub264 = (a263 & b_inv263) | (a263 & c263) | (b_inv263 & c263);
  wire s264, sub264, and264, or264;
  wire b_inv264;
  assign b_inv264 = ~b264;
  assign s264  = a264 ^ b264 ^ c264;
  assign sub264 = a264 ^ b_inv264 ^ c264;
  assign and264 = a264 & b264;
  assign or264  = a264 | b264;
  assign c265 = (a264 & b264) | (a264 & c264) | (b264 & c264);
  wire c_sub265;
  assign c_sub265 = (a264 & b_inv264) | (a264 & c264) | (b_inv264 & c264);
  wire s265, sub265, and265, or265;
  wire b_inv265;
  assign b_inv265 = ~b265;
  assign s265  = a265 ^ b265 ^ c265;
  assign sub265 = a265 ^ b_inv265 ^ c265;
  assign and265 = a265 & b265;
  assign or265  = a265 | b265;
  assign c266 = (a265 & b265) | (a265 & c265) | (b265 & c265);
  wire c_sub266;
  assign c_sub266 = (a265 & b_inv265) | (a265 & c265) | (b_inv265 & c265);
  wire s266, sub266, and266, or266;
  wire b_inv266;
  assign b_inv266 = ~b266;
  assign s266  = a266 ^ b266 ^ c266;
  assign sub266 = a266 ^ b_inv266 ^ c266;
  assign and266 = a266 & b266;
  assign or266  = a266 | b266;
  assign c267 = (a266 & b266) | (a266 & c266) | (b266 & c266);
  wire c_sub267;
  assign c_sub267 = (a266 & b_inv266) | (a266 & c266) | (b_inv266 & c266);
  wire s267, sub267, and267, or267;
  wire b_inv267;
  assign b_inv267 = ~b267;
  assign s267  = a267 ^ b267 ^ c267;
  assign sub267 = a267 ^ b_inv267 ^ c267;
  assign and267 = a267 & b267;
  assign or267  = a267 | b267;
  assign c268 = (a267 & b267) | (a267 & c267) | (b267 & c267);
  wire c_sub268;
  assign c_sub268 = (a267 & b_inv267) | (a267 & c267) | (b_inv267 & c267);
  wire s268, sub268, and268, or268;
  wire b_inv268;
  assign b_inv268 = ~b268;
  assign s268  = a268 ^ b268 ^ c268;
  assign sub268 = a268 ^ b_inv268 ^ c268;
  assign and268 = a268 & b268;
  assign or268  = a268 | b268;
  assign c269 = (a268 & b268) | (a268 & c268) | (b268 & c268);
  wire c_sub269;
  assign c_sub269 = (a268 & b_inv268) | (a268 & c268) | (b_inv268 & c268);
  wire s269, sub269, and269, or269;
  wire b_inv269;
  assign b_inv269 = ~b269;
  assign s269  = a269 ^ b269 ^ c269;
  assign sub269 = a269 ^ b_inv269 ^ c269;
  assign and269 = a269 & b269;
  assign or269  = a269 | b269;
  assign c270 = (a269 & b269) | (a269 & c269) | (b269 & c269);
  wire c_sub270;
  assign c_sub270 = (a269 & b_inv269) | (a269 & c269) | (b_inv269 & c269);
  wire s270, sub270, and270, or270;
  wire b_inv270;
  assign b_inv270 = ~b270;
  assign s270  = a270 ^ b270 ^ c270;
  assign sub270 = a270 ^ b_inv270 ^ c270;
  assign and270 = a270 & b270;
  assign or270  = a270 | b270;
  assign c271 = (a270 & b270) | (a270 & c270) | (b270 & c270);
  wire c_sub271;
  assign c_sub271 = (a270 & b_inv270) | (a270 & c270) | (b_inv270 & c270);
  wire s271, sub271, and271, or271;
  wire b_inv271;
  assign b_inv271 = ~b271;
  assign s271  = a271 ^ b271 ^ c271;
  assign sub271 = a271 ^ b_inv271 ^ c271;
  assign and271 = a271 & b271;
  assign or271  = a271 | b271;
  assign c272 = (a271 & b271) | (a271 & c271) | (b271 & c271);
  wire c_sub272;
  assign c_sub272 = (a271 & b_inv271) | (a271 & c271) | (b_inv271 & c271);
  wire s272, sub272, and272, or272;
  wire b_inv272;
  assign b_inv272 = ~b272;
  assign s272  = a272 ^ b272 ^ c272;
  assign sub272 = a272 ^ b_inv272 ^ c272;
  assign and272 = a272 & b272;
  assign or272  = a272 | b272;
  assign c273 = (a272 & b272) | (a272 & c272) | (b272 & c272);
  wire c_sub273;
  assign c_sub273 = (a272 & b_inv272) | (a272 & c272) | (b_inv272 & c272);
  wire s273, sub273, and273, or273;
  wire b_inv273;
  assign b_inv273 = ~b273;
  assign s273  = a273 ^ b273 ^ c273;
  assign sub273 = a273 ^ b_inv273 ^ c273;
  assign and273 = a273 & b273;
  assign or273  = a273 | b273;
  assign c274 = (a273 & b273) | (a273 & c273) | (b273 & c273);
  wire c_sub274;
  assign c_sub274 = (a273 & b_inv273) | (a273 & c273) | (b_inv273 & c273);
  wire s274, sub274, and274, or274;
  wire b_inv274;
  assign b_inv274 = ~b274;
  assign s274  = a274 ^ b274 ^ c274;
  assign sub274 = a274 ^ b_inv274 ^ c274;
  assign and274 = a274 & b274;
  assign or274  = a274 | b274;
  assign c275 = (a274 & b274) | (a274 & c274) | (b274 & c274);
  wire c_sub275;
  assign c_sub275 = (a274 & b_inv274) | (a274 & c274) | (b_inv274 & c274);
  wire s275, sub275, and275, or275;
  wire b_inv275;
  assign b_inv275 = ~b275;
  assign s275  = a275 ^ b275 ^ c275;
  assign sub275 = a275 ^ b_inv275 ^ c275;
  assign and275 = a275 & b275;
  assign or275  = a275 | b275;
  assign c276 = (a275 & b275) | (a275 & c275) | (b275 & c275);
  wire c_sub276;
  assign c_sub276 = (a275 & b_inv275) | (a275 & c275) | (b_inv275 & c275);
  wire s276, sub276, and276, or276;
  wire b_inv276;
  assign b_inv276 = ~b276;
  assign s276  = a276 ^ b276 ^ c276;
  assign sub276 = a276 ^ b_inv276 ^ c276;
  assign and276 = a276 & b276;
  assign or276  = a276 | b276;
  assign c277 = (a276 & b276) | (a276 & c276) | (b276 & c276);
  wire c_sub277;
  assign c_sub277 = (a276 & b_inv276) | (a276 & c276) | (b_inv276 & c276);
  wire s277, sub277, and277, or277;
  wire b_inv277;
  assign b_inv277 = ~b277;
  assign s277  = a277 ^ b277 ^ c277;
  assign sub277 = a277 ^ b_inv277 ^ c277;
  assign and277 = a277 & b277;
  assign or277  = a277 | b277;
  assign c278 = (a277 & b277) | (a277 & c277) | (b277 & c277);
  wire c_sub278;
  assign c_sub278 = (a277 & b_inv277) | (a277 & c277) | (b_inv277 & c277);
  wire s278, sub278, and278, or278;
  wire b_inv278;
  assign b_inv278 = ~b278;
  assign s278  = a278 ^ b278 ^ c278;
  assign sub278 = a278 ^ b_inv278 ^ c278;
  assign and278 = a278 & b278;
  assign or278  = a278 | b278;
  assign c279 = (a278 & b278) | (a278 & c278) | (b278 & c278);
  wire c_sub279;
  assign c_sub279 = (a278 & b_inv278) | (a278 & c278) | (b_inv278 & c278);
  wire s279, sub279, and279, or279;
  wire b_inv279;
  assign b_inv279 = ~b279;
  assign s279  = a279 ^ b279 ^ c279;
  assign sub279 = a279 ^ b_inv279 ^ c279;
  assign and279 = a279 & b279;
  assign or279  = a279 | b279;
  assign c280 = (a279 & b279) | (a279 & c279) | (b279 & c279);
  wire c_sub280;
  assign c_sub280 = (a279 & b_inv279) | (a279 & c279) | (b_inv279 & c279);
  wire s280, sub280, and280, or280;
  wire b_inv280;
  assign b_inv280 = ~b280;
  assign s280  = a280 ^ b280 ^ c280;
  assign sub280 = a280 ^ b_inv280 ^ c280;
  assign and280 = a280 & b280;
  assign or280  = a280 | b280;
  assign c281 = (a280 & b280) | (a280 & c280) | (b280 & c280);
  wire c_sub281;
  assign c_sub281 = (a280 & b_inv280) | (a280 & c280) | (b_inv280 & c280);
  wire s281, sub281, and281, or281;
  wire b_inv281;
  assign b_inv281 = ~b281;
  assign s281  = a281 ^ b281 ^ c281;
  assign sub281 = a281 ^ b_inv281 ^ c281;
  assign and281 = a281 & b281;
  assign or281  = a281 | b281;
  assign c282 = (a281 & b281) | (a281 & c281) | (b281 & c281);
  wire c_sub282;
  assign c_sub282 = (a281 & b_inv281) | (a281 & c281) | (b_inv281 & c281);
  wire s282, sub282, and282, or282;
  wire b_inv282;
  assign b_inv282 = ~b282;
  assign s282  = a282 ^ b282 ^ c282;
  assign sub282 = a282 ^ b_inv282 ^ c282;
  assign and282 = a282 & b282;
  assign or282  = a282 | b282;
  assign c283 = (a282 & b282) | (a282 & c282) | (b282 & c282);
  wire c_sub283;
  assign c_sub283 = (a282 & b_inv282) | (a282 & c282) | (b_inv282 & c282);
  wire s283, sub283, and283, or283;
  wire b_inv283;
  assign b_inv283 = ~b283;
  assign s283  = a283 ^ b283 ^ c283;
  assign sub283 = a283 ^ b_inv283 ^ c283;
  assign and283 = a283 & b283;
  assign or283  = a283 | b283;
  assign c284 = (a283 & b283) | (a283 & c283) | (b283 & c283);
  wire c_sub284;
  assign c_sub284 = (a283 & b_inv283) | (a283 & c283) | (b_inv283 & c283);
  wire s284, sub284, and284, or284;
  wire b_inv284;
  assign b_inv284 = ~b284;
  assign s284  = a284 ^ b284 ^ c284;
  assign sub284 = a284 ^ b_inv284 ^ c284;
  assign and284 = a284 & b284;
  assign or284  = a284 | b284;
  assign c285 = (a284 & b284) | (a284 & c284) | (b284 & c284);
  wire c_sub285;
  assign c_sub285 = (a284 & b_inv284) | (a284 & c284) | (b_inv284 & c284);
  wire s285, sub285, and285, or285;
  wire b_inv285;
  assign b_inv285 = ~b285;
  assign s285  = a285 ^ b285 ^ c285;
  assign sub285 = a285 ^ b_inv285 ^ c285;
  assign and285 = a285 & b285;
  assign or285  = a285 | b285;
  assign c286 = (a285 & b285) | (a285 & c285) | (b285 & c285);
  wire c_sub286;
  assign c_sub286 = (a285 & b_inv285) | (a285 & c285) | (b_inv285 & c285);
  wire s286, sub286, and286, or286;
  wire b_inv286;
  assign b_inv286 = ~b286;
  assign s286  = a286 ^ b286 ^ c286;
  assign sub286 = a286 ^ b_inv286 ^ c286;
  assign and286 = a286 & b286;
  assign or286  = a286 | b286;
  assign c287 = (a286 & b286) | (a286 & c286) | (b286 & c286);
  wire c_sub287;
  assign c_sub287 = (a286 & b_inv286) | (a286 & c286) | (b_inv286 & c286);
  wire s287, sub287, and287, or287;
  wire b_inv287;
  assign b_inv287 = ~b287;
  assign s287  = a287 ^ b287 ^ c287;
  assign sub287 = a287 ^ b_inv287 ^ c287;
  assign and287 = a287 & b287;
  assign or287  = a287 | b287;
  assign c288 = (a287 & b287) | (a287 & c287) | (b287 & c287);
  wire c_sub288;
  assign c_sub288 = (a287 & b_inv287) | (a287 & c287) | (b_inv287 & c287);
  wire s288, sub288, and288, or288;
  wire b_inv288;
  assign b_inv288 = ~b288;
  assign s288  = a288 ^ b288 ^ c288;
  assign sub288 = a288 ^ b_inv288 ^ c288;
  assign and288 = a288 & b288;
  assign or288  = a288 | b288;
  assign c289 = (a288 & b288) | (a288 & c288) | (b288 & c288);
  wire c_sub289;
  assign c_sub289 = (a288 & b_inv288) | (a288 & c288) | (b_inv288 & c288);
  wire s289, sub289, and289, or289;
  wire b_inv289;
  assign b_inv289 = ~b289;
  assign s289  = a289 ^ b289 ^ c289;
  assign sub289 = a289 ^ b_inv289 ^ c289;
  assign and289 = a289 & b289;
  assign or289  = a289 | b289;
  assign c290 = (a289 & b289) | (a289 & c289) | (b289 & c289);
  wire c_sub290;
  assign c_sub290 = (a289 & b_inv289) | (a289 & c289) | (b_inv289 & c289);
  wire s290, sub290, and290, or290;
  wire b_inv290;
  assign b_inv290 = ~b290;
  assign s290  = a290 ^ b290 ^ c290;
  assign sub290 = a290 ^ b_inv290 ^ c290;
  assign and290 = a290 & b290;
  assign or290  = a290 | b290;
  assign c291 = (a290 & b290) | (a290 & c290) | (b290 & c290);
  wire c_sub291;
  assign c_sub291 = (a290 & b_inv290) | (a290 & c290) | (b_inv290 & c290);
  wire s291, sub291, and291, or291;
  wire b_inv291;
  assign b_inv291 = ~b291;
  assign s291  = a291 ^ b291 ^ c291;
  assign sub291 = a291 ^ b_inv291 ^ c291;
  assign and291 = a291 & b291;
  assign or291  = a291 | b291;
  assign c292 = (a291 & b291) | (a291 & c291) | (b291 & c291);
  wire c_sub292;
  assign c_sub292 = (a291 & b_inv291) | (a291 & c291) | (b_inv291 & c291);
  wire s292, sub292, and292, or292;
  wire b_inv292;
  assign b_inv292 = ~b292;
  assign s292  = a292 ^ b292 ^ c292;
  assign sub292 = a292 ^ b_inv292 ^ c292;
  assign and292 = a292 & b292;
  assign or292  = a292 | b292;
  assign c293 = (a292 & b292) | (a292 & c292) | (b292 & c292);
  wire c_sub293;
  assign c_sub293 = (a292 & b_inv292) | (a292 & c292) | (b_inv292 & c292);
  wire s293, sub293, and293, or293;
  wire b_inv293;
  assign b_inv293 = ~b293;
  assign s293  = a293 ^ b293 ^ c293;
  assign sub293 = a293 ^ b_inv293 ^ c293;
  assign and293 = a293 & b293;
  assign or293  = a293 | b293;
  assign c294 = (a293 & b293) | (a293 & c293) | (b293 & c293);
  wire c_sub294;
  assign c_sub294 = (a293 & b_inv293) | (a293 & c293) | (b_inv293 & c293);
  wire s294, sub294, and294, or294;
  wire b_inv294;
  assign b_inv294 = ~b294;
  assign s294  = a294 ^ b294 ^ c294;
  assign sub294 = a294 ^ b_inv294 ^ c294;
  assign and294 = a294 & b294;
  assign or294  = a294 | b294;
  assign c295 = (a294 & b294) | (a294 & c294) | (b294 & c294);
  wire c_sub295;
  assign c_sub295 = (a294 & b_inv294) | (a294 & c294) | (b_inv294 & c294);
  wire s295, sub295, and295, or295;
  wire b_inv295;
  assign b_inv295 = ~b295;
  assign s295  = a295 ^ b295 ^ c295;
  assign sub295 = a295 ^ b_inv295 ^ c295;
  assign and295 = a295 & b295;
  assign or295  = a295 | b295;
  assign c296 = (a295 & b295) | (a295 & c295) | (b295 & c295);
  wire c_sub296;
  assign c_sub296 = (a295 & b_inv295) | (a295 & c295) | (b_inv295 & c295);
  wire s296, sub296, and296, or296;
  wire b_inv296;
  assign b_inv296 = ~b296;
  assign s296  = a296 ^ b296 ^ c296;
  assign sub296 = a296 ^ b_inv296 ^ c296;
  assign and296 = a296 & b296;
  assign or296  = a296 | b296;
  assign c297 = (a296 & b296) | (a296 & c296) | (b296 & c296);
  wire c_sub297;
  assign c_sub297 = (a296 & b_inv296) | (a296 & c296) | (b_inv296 & c296);
  wire s297, sub297, and297, or297;
  wire b_inv297;
  assign b_inv297 = ~b297;
  assign s297  = a297 ^ b297 ^ c297;
  assign sub297 = a297 ^ b_inv297 ^ c297;
  assign and297 = a297 & b297;
  assign or297  = a297 | b297;
  assign c298 = (a297 & b297) | (a297 & c297) | (b297 & c297);
  wire c_sub298;
  assign c_sub298 = (a297 & b_inv297) | (a297 & c297) | (b_inv297 & c297);
  wire s298, sub298, and298, or298;
  wire b_inv298;
  assign b_inv298 = ~b298;
  assign s298  = a298 ^ b298 ^ c298;
  assign sub298 = a298 ^ b_inv298 ^ c298;
  assign and298 = a298 & b298;
  assign or298  = a298 | b298;
  assign c299 = (a298 & b298) | (a298 & c298) | (b298 & c298);
  wire c_sub299;
  assign c_sub299 = (a298 & b_inv298) | (a298 & c298) | (b_inv298 & c298);
  wire s299, sub299, and299, or299;
  wire b_inv299;
  assign b_inv299 = ~b299;
  assign s299  = a299 ^ b299 ^ c299;
  assign sub299 = a299 ^ b_inv299 ^ c299;
  assign and299 = a299 & b299;
  assign or299  = a299 | b299;
  assign c300 = (a299 & b299) | (a299 & c299) | (b299 & c299);
  wire c_sub300;
  assign c_sub300 = (a299 & b_inv299) | (a299 & c299) | (b_inv299 & c299);
  wire s300, sub300, and300, or300;
  wire b_inv300;
  assign b_inv300 = ~b300;
  assign s300  = a300 ^ b300 ^ c300;
  assign sub300 = a300 ^ b_inv300 ^ c300;
  assign and300 = a300 & b300;
  assign or300  = a300 | b300;
  assign c301 = (a300 & b300) | (a300 & c300) | (b300 & c300);
  wire c_sub301;
  assign c_sub301 = (a300 & b_inv300) | (a300 & c300) | (b_inv300 & c300);
  wire s301, sub301, and301, or301;
  wire b_inv301;
  assign b_inv301 = ~b301;
  assign s301  = a301 ^ b301 ^ c301;
  assign sub301 = a301 ^ b_inv301 ^ c301;
  assign and301 = a301 & b301;
  assign or301  = a301 | b301;
  assign c302 = (a301 & b301) | (a301 & c301) | (b301 & c301);
  wire c_sub302;
  assign c_sub302 = (a301 & b_inv301) | (a301 & c301) | (b_inv301 & c301);
  wire s302, sub302, and302, or302;
  wire b_inv302;
  assign b_inv302 = ~b302;
  assign s302  = a302 ^ b302 ^ c302;
  assign sub302 = a302 ^ b_inv302 ^ c302;
  assign and302 = a302 & b302;
  assign or302  = a302 | b302;
  assign c303 = (a302 & b302) | (a302 & c302) | (b302 & c302);
  wire c_sub303;
  assign c_sub303 = (a302 & b_inv302) | (a302 & c302) | (b_inv302 & c302);
  wire s303, sub303, and303, or303;
  wire b_inv303;
  assign b_inv303 = ~b303;
  assign s303  = a303 ^ b303 ^ c303;
  assign sub303 = a303 ^ b_inv303 ^ c303;
  assign and303 = a303 & b303;
  assign or303  = a303 | b303;
  assign c304 = (a303 & b303) | (a303 & c303) | (b303 & c303);
  wire c_sub304;
  assign c_sub304 = (a303 & b_inv303) | (a303 & c303) | (b_inv303 & c303);
  wire s304, sub304, and304, or304;
  wire b_inv304;
  assign b_inv304 = ~b304;
  assign s304  = a304 ^ b304 ^ c304;
  assign sub304 = a304 ^ b_inv304 ^ c304;
  assign and304 = a304 & b304;
  assign or304  = a304 | b304;
  assign c305 = (a304 & b304) | (a304 & c304) | (b304 & c304);
  wire c_sub305;
  assign c_sub305 = (a304 & b_inv304) | (a304 & c304) | (b_inv304 & c304);
  wire s305, sub305, and305, or305;
  wire b_inv305;
  assign b_inv305 = ~b305;
  assign s305  = a305 ^ b305 ^ c305;
  assign sub305 = a305 ^ b_inv305 ^ c305;
  assign and305 = a305 & b305;
  assign or305  = a305 | b305;
  assign c306 = (a305 & b305) | (a305 & c305) | (b305 & c305);
  wire c_sub306;
  assign c_sub306 = (a305 & b_inv305) | (a305 & c305) | (b_inv305 & c305);
  wire s306, sub306, and306, or306;
  wire b_inv306;
  assign b_inv306 = ~b306;
  assign s306  = a306 ^ b306 ^ c306;
  assign sub306 = a306 ^ b_inv306 ^ c306;
  assign and306 = a306 & b306;
  assign or306  = a306 | b306;
  assign c307 = (a306 & b306) | (a306 & c306) | (b306 & c306);
  wire c_sub307;
  assign c_sub307 = (a306 & b_inv306) | (a306 & c306) | (b_inv306 & c306);
  wire s307, sub307, and307, or307;
  wire b_inv307;
  assign b_inv307 = ~b307;
  assign s307  = a307 ^ b307 ^ c307;
  assign sub307 = a307 ^ b_inv307 ^ c307;
  assign and307 = a307 & b307;
  assign or307  = a307 | b307;
  assign c308 = (a307 & b307) | (a307 & c307) | (b307 & c307);
  wire c_sub308;
  assign c_sub308 = (a307 & b_inv307) | (a307 & c307) | (b_inv307 & c307);
  wire s308, sub308, and308, or308;
  wire b_inv308;
  assign b_inv308 = ~b308;
  assign s308  = a308 ^ b308 ^ c308;
  assign sub308 = a308 ^ b_inv308 ^ c308;
  assign and308 = a308 & b308;
  assign or308  = a308 | b308;
  assign c309 = (a308 & b308) | (a308 & c308) | (b308 & c308);
  wire c_sub309;
  assign c_sub309 = (a308 & b_inv308) | (a308 & c308) | (b_inv308 & c308);
  wire s309, sub309, and309, or309;
  wire b_inv309;
  assign b_inv309 = ~b309;
  assign s309  = a309 ^ b309 ^ c309;
  assign sub309 = a309 ^ b_inv309 ^ c309;
  assign and309 = a309 & b309;
  assign or309  = a309 | b309;
  assign c310 = (a309 & b309) | (a309 & c309) | (b309 & c309);
  wire c_sub310;
  assign c_sub310 = (a309 & b_inv309) | (a309 & c309) | (b_inv309 & c309);
  wire s310, sub310, and310, or310;
  wire b_inv310;
  assign b_inv310 = ~b310;
  assign s310  = a310 ^ b310 ^ c310;
  assign sub310 = a310 ^ b_inv310 ^ c310;
  assign and310 = a310 & b310;
  assign or310  = a310 | b310;
  assign c311 = (a310 & b310) | (a310 & c310) | (b310 & c310);
  wire c_sub311;
  assign c_sub311 = (a310 & b_inv310) | (a310 & c310) | (b_inv310 & c310);
  wire s311, sub311, and311, or311;
  wire b_inv311;
  assign b_inv311 = ~b311;
  assign s311  = a311 ^ b311 ^ c311;
  assign sub311 = a311 ^ b_inv311 ^ c311;
  assign and311 = a311 & b311;
  assign or311  = a311 | b311;
  assign c312 = (a311 & b311) | (a311 & c311) | (b311 & c311);
  wire c_sub312;
  assign c_sub312 = (a311 & b_inv311) | (a311 & c311) | (b_inv311 & c311);
  wire s312, sub312, and312, or312;
  wire b_inv312;
  assign b_inv312 = ~b312;
  assign s312  = a312 ^ b312 ^ c312;
  assign sub312 = a312 ^ b_inv312 ^ c312;
  assign and312 = a312 & b312;
  assign or312  = a312 | b312;
  assign c313 = (a312 & b312) | (a312 & c312) | (b312 & c312);
  wire c_sub313;
  assign c_sub313 = (a312 & b_inv312) | (a312 & c312) | (b_inv312 & c312);
  wire s313, sub313, and313, or313;
  wire b_inv313;
  assign b_inv313 = ~b313;
  assign s313  = a313 ^ b313 ^ c313;
  assign sub313 = a313 ^ b_inv313 ^ c313;
  assign and313 = a313 & b313;
  assign or313  = a313 | b313;
  assign c314 = (a313 & b313) | (a313 & c313) | (b313 & c313);
  wire c_sub314;
  assign c_sub314 = (a313 & b_inv313) | (a313 & c313) | (b_inv313 & c313);
  wire s314, sub314, and314, or314;
  wire b_inv314;
  assign b_inv314 = ~b314;
  assign s314  = a314 ^ b314 ^ c314;
  assign sub314 = a314 ^ b_inv314 ^ c314;
  assign and314 = a314 & b314;
  assign or314  = a314 | b314;
  assign c315 = (a314 & b314) | (a314 & c314) | (b314 & c314);
  wire c_sub315;
  assign c_sub315 = (a314 & b_inv314) | (a314 & c314) | (b_inv314 & c314);
  wire s315, sub315, and315, or315;
  wire b_inv315;
  assign b_inv315 = ~b315;
  assign s315  = a315 ^ b315 ^ c315;
  assign sub315 = a315 ^ b_inv315 ^ c315;
  assign and315 = a315 & b315;
  assign or315  = a315 | b315;
  assign c316 = (a315 & b315) | (a315 & c315) | (b315 & c315);
  wire c_sub316;
  assign c_sub316 = (a315 & b_inv315) | (a315 & c315) | (b_inv315 & c315);
  wire s316, sub316, and316, or316;
  wire b_inv316;
  assign b_inv316 = ~b316;
  assign s316  = a316 ^ b316 ^ c316;
  assign sub316 = a316 ^ b_inv316 ^ c316;
  assign and316 = a316 & b316;
  assign or316  = a316 | b316;
  assign c317 = (a316 & b316) | (a316 & c316) | (b316 & c316);
  wire c_sub317;
  assign c_sub317 = (a316 & b_inv316) | (a316 & c316) | (b_inv316 & c316);
  wire s317, sub317, and317, or317;
  wire b_inv317;
  assign b_inv317 = ~b317;
  assign s317  = a317 ^ b317 ^ c317;
  assign sub317 = a317 ^ b_inv317 ^ c317;
  assign and317 = a317 & b317;
  assign or317  = a317 | b317;
  assign c318 = (a317 & b317) | (a317 & c317) | (b317 & c317);
  wire c_sub318;
  assign c_sub318 = (a317 & b_inv317) | (a317 & c317) | (b_inv317 & c317);
  wire s318, sub318, and318, or318;
  wire b_inv318;
  assign b_inv318 = ~b318;
  assign s318  = a318 ^ b318 ^ c318;
  assign sub318 = a318 ^ b_inv318 ^ c318;
  assign and318 = a318 & b318;
  assign or318  = a318 | b318;
  assign c319 = (a318 & b318) | (a318 & c318) | (b318 & c318);
  wire c_sub319;
  assign c_sub319 = (a318 & b_inv318) | (a318 & c318) | (b_inv318 & c318);
  wire s319, sub319, and319, or319;
  wire b_inv319;
  assign b_inv319 = ~b319;
  assign s319  = a319 ^ b319 ^ c319;
  assign sub319 = a319 ^ b_inv319 ^ c319;
  assign and319 = a319 & b319;
  assign or319  = a319 | b319;
  assign c320 = (a319 & b319) | (a319 & c319) | (b319 & c319);
  wire c_sub320;
  assign c_sub320 = (a319 & b_inv319) | (a319 & c319) | (b_inv319 & c319);
  wire s320, sub320, and320, or320;
  wire b_inv320;
  assign b_inv320 = ~b320;
  assign s320  = a320 ^ b320 ^ c320;
  assign sub320 = a320 ^ b_inv320 ^ c320;
  assign and320 = a320 & b320;
  assign or320  = a320 | b320;
  assign c321 = (a320 & b320) | (a320 & c320) | (b320 & c320);
  wire c_sub321;
  assign c_sub321 = (a320 & b_inv320) | (a320 & c320) | (b_inv320 & c320);
  wire s321, sub321, and321, or321;
  wire b_inv321;
  assign b_inv321 = ~b321;
  assign s321  = a321 ^ b321 ^ c321;
  assign sub321 = a321 ^ b_inv321 ^ c321;
  assign and321 = a321 & b321;
  assign or321  = a321 | b321;
  assign c322 = (a321 & b321) | (a321 & c321) | (b321 & c321);
  wire c_sub322;
  assign c_sub322 = (a321 & b_inv321) | (a321 & c321) | (b_inv321 & c321);
  wire s322, sub322, and322, or322;
  wire b_inv322;
  assign b_inv322 = ~b322;
  assign s322  = a322 ^ b322 ^ c322;
  assign sub322 = a322 ^ b_inv322 ^ c322;
  assign and322 = a322 & b322;
  assign or322  = a322 | b322;
  assign c323 = (a322 & b322) | (a322 & c322) | (b322 & c322);
  wire c_sub323;
  assign c_sub323 = (a322 & b_inv322) | (a322 & c322) | (b_inv322 & c322);
  wire s323, sub323, and323, or323;
  wire b_inv323;
  assign b_inv323 = ~b323;
  assign s323  = a323 ^ b323 ^ c323;
  assign sub323 = a323 ^ b_inv323 ^ c323;
  assign and323 = a323 & b323;
  assign or323  = a323 | b323;
  assign c324 = (a323 & b323) | (a323 & c323) | (b323 & c323);
  wire c_sub324;
  assign c_sub324 = (a323 & b_inv323) | (a323 & c323) | (b_inv323 & c323);
  wire s324, sub324, and324, or324;
  wire b_inv324;
  assign b_inv324 = ~b324;
  assign s324  = a324 ^ b324 ^ c324;
  assign sub324 = a324 ^ b_inv324 ^ c324;
  assign and324 = a324 & b324;
  assign or324  = a324 | b324;
  assign c325 = (a324 & b324) | (a324 & c324) | (b324 & c324);
  wire c_sub325;
  assign c_sub325 = (a324 & b_inv324) | (a324 & c324) | (b_inv324 & c324);
  wire s325, sub325, and325, or325;
  wire b_inv325;
  assign b_inv325 = ~b325;
  assign s325  = a325 ^ b325 ^ c325;
  assign sub325 = a325 ^ b_inv325 ^ c325;
  assign and325 = a325 & b325;
  assign or325  = a325 | b325;
  assign c326 = (a325 & b325) | (a325 & c325) | (b325 & c325);
  wire c_sub326;
  assign c_sub326 = (a325 & b_inv325) | (a325 & c325) | (b_inv325 & c325);
  wire s326, sub326, and326, or326;
  wire b_inv326;
  assign b_inv326 = ~b326;
  assign s326  = a326 ^ b326 ^ c326;
  assign sub326 = a326 ^ b_inv326 ^ c326;
  assign and326 = a326 & b326;
  assign or326  = a326 | b326;
  assign c327 = (a326 & b326) | (a326 & c326) | (b326 & c326);
  wire c_sub327;
  assign c_sub327 = (a326 & b_inv326) | (a326 & c326) | (b_inv326 & c326);
  wire s327, sub327, and327, or327;
  wire b_inv327;
  assign b_inv327 = ~b327;
  assign s327  = a327 ^ b327 ^ c327;
  assign sub327 = a327 ^ b_inv327 ^ c327;
  assign and327 = a327 & b327;
  assign or327  = a327 | b327;
  assign c328 = (a327 & b327) | (a327 & c327) | (b327 & c327);
  wire c_sub328;
  assign c_sub328 = (a327 & b_inv327) | (a327 & c327) | (b_inv327 & c327);
  wire s328, sub328, and328, or328;
  wire b_inv328;
  assign b_inv328 = ~b328;
  assign s328  = a328 ^ b328 ^ c328;
  assign sub328 = a328 ^ b_inv328 ^ c328;
  assign and328 = a328 & b328;
  assign or328  = a328 | b328;
  assign c329 = (a328 & b328) | (a328 & c328) | (b328 & c328);
  wire c_sub329;
  assign c_sub329 = (a328 & b_inv328) | (a328 & c328) | (b_inv328 & c328);
  wire s329, sub329, and329, or329;
  wire b_inv329;
  assign b_inv329 = ~b329;
  assign s329  = a329 ^ b329 ^ c329;
  assign sub329 = a329 ^ b_inv329 ^ c329;
  assign and329 = a329 & b329;
  assign or329  = a329 | b329;
  assign c330 = (a329 & b329) | (a329 & c329) | (b329 & c329);
  wire c_sub330;
  assign c_sub330 = (a329 & b_inv329) | (a329 & c329) | (b_inv329 & c329);
  wire s330, sub330, and330, or330;
  wire b_inv330;
  assign b_inv330 = ~b330;
  assign s330  = a330 ^ b330 ^ c330;
  assign sub330 = a330 ^ b_inv330 ^ c330;
  assign and330 = a330 & b330;
  assign or330  = a330 | b330;
  assign c331 = (a330 & b330) | (a330 & c330) | (b330 & c330);
  wire c_sub331;
  assign c_sub331 = (a330 & b_inv330) | (a330 & c330) | (b_inv330 & c330);
  wire s331, sub331, and331, or331;
  wire b_inv331;
  assign b_inv331 = ~b331;
  assign s331  = a331 ^ b331 ^ c331;
  assign sub331 = a331 ^ b_inv331 ^ c331;
  assign and331 = a331 & b331;
  assign or331  = a331 | b331;
  assign c332 = (a331 & b331) | (a331 & c331) | (b331 & c331);
  wire c_sub332;
  assign c_sub332 = (a331 & b_inv331) | (a331 & c331) | (b_inv331 & c331);
  wire s332, sub332, and332, or332;
  wire b_inv332;
  assign b_inv332 = ~b332;
  assign s332  = a332 ^ b332 ^ c332;
  assign sub332 = a332 ^ b_inv332 ^ c332;
  assign and332 = a332 & b332;
  assign or332  = a332 | b332;
  assign c333 = (a332 & b332) | (a332 & c332) | (b332 & c332);
  wire c_sub333;
  assign c_sub333 = (a332 & b_inv332) | (a332 & c332) | (b_inv332 & c332);
  wire s333, sub333, and333, or333;
  wire b_inv333;
  assign b_inv333 = ~b333;
  assign s333  = a333 ^ b333 ^ c333;
  assign sub333 = a333 ^ b_inv333 ^ c333;
  assign and333 = a333 & b333;
  assign or333  = a333 | b333;
  assign c334 = (a333 & b333) | (a333 & c333) | (b333 & c333);
  wire c_sub334;
  assign c_sub334 = (a333 & b_inv333) | (a333 & c333) | (b_inv333 & c333);
  wire s334, sub334, and334, or334;
  wire b_inv334;
  assign b_inv334 = ~b334;
  assign s334  = a334 ^ b334 ^ c334;
  assign sub334 = a334 ^ b_inv334 ^ c334;
  assign and334 = a334 & b334;
  assign or334  = a334 | b334;
  assign c335 = (a334 & b334) | (a334 & c334) | (b334 & c334);
  wire c_sub335;
  assign c_sub335 = (a334 & b_inv334) | (a334 & c334) | (b_inv334 & c334);
  wire s335, sub335, and335, or335;
  wire b_inv335;
  assign b_inv335 = ~b335;
  assign s335  = a335 ^ b335 ^ c335;
  assign sub335 = a335 ^ b_inv335 ^ c335;
  assign and335 = a335 & b335;
  assign or335  = a335 | b335;
  assign c336 = (a335 & b335) | (a335 & c335) | (b335 & c335);
  wire c_sub336;
  assign c_sub336 = (a335 & b_inv335) | (a335 & c335) | (b_inv335 & c335);
  wire s336, sub336, and336, or336;
  wire b_inv336;
  assign b_inv336 = ~b336;
  assign s336  = a336 ^ b336 ^ c336;
  assign sub336 = a336 ^ b_inv336 ^ c336;
  assign and336 = a336 & b336;
  assign or336  = a336 | b336;
  assign c337 = (a336 & b336) | (a336 & c336) | (b336 & c336);
  wire c_sub337;
  assign c_sub337 = (a336 & b_inv336) | (a336 & c336) | (b_inv336 & c336);
  wire s337, sub337, and337, or337;
  wire b_inv337;
  assign b_inv337 = ~b337;
  assign s337  = a337 ^ b337 ^ c337;
  assign sub337 = a337 ^ b_inv337 ^ c337;
  assign and337 = a337 & b337;
  assign or337  = a337 | b337;
  assign c338 = (a337 & b337) | (a337 & c337) | (b337 & c337);
  wire c_sub338;
  assign c_sub338 = (a337 & b_inv337) | (a337 & c337) | (b_inv337 & c337);
  wire s338, sub338, and338, or338;
  wire b_inv338;
  assign b_inv338 = ~b338;
  assign s338  = a338 ^ b338 ^ c338;
  assign sub338 = a338 ^ b_inv338 ^ c338;
  assign and338 = a338 & b338;
  assign or338  = a338 | b338;
  assign c339 = (a338 & b338) | (a338 & c338) | (b338 & c338);
  wire c_sub339;
  assign c_sub339 = (a338 & b_inv338) | (a338 & c338) | (b_inv338 & c338);
  wire s339, sub339, and339, or339;
  wire b_inv339;
  assign b_inv339 = ~b339;
  assign s339  = a339 ^ b339 ^ c339;
  assign sub339 = a339 ^ b_inv339 ^ c339;
  assign and339 = a339 & b339;
  assign or339  = a339 | b339;
  assign c340 = (a339 & b339) | (a339 & c339) | (b339 & c339);
  wire c_sub340;
  assign c_sub340 = (a339 & b_inv339) | (a339 & c339) | (b_inv339 & c339);
  wire s340, sub340, and340, or340;
  wire b_inv340;
  assign b_inv340 = ~b340;
  assign s340  = a340 ^ b340 ^ c340;
  assign sub340 = a340 ^ b_inv340 ^ c340;
  assign and340 = a340 & b340;
  assign or340  = a340 | b340;
  assign c341 = (a340 & b340) | (a340 & c340) | (b340 & c340);
  wire c_sub341;
  assign c_sub341 = (a340 & b_inv340) | (a340 & c340) | (b_inv340 & c340);
  wire s341, sub341, and341, or341;
  wire b_inv341;
  assign b_inv341 = ~b341;
  assign s341  = a341 ^ b341 ^ c341;
  assign sub341 = a341 ^ b_inv341 ^ c341;
  assign and341 = a341 & b341;
  assign or341  = a341 | b341;
  assign c342 = (a341 & b341) | (a341 & c341) | (b341 & c341);
  wire c_sub342;
  assign c_sub342 = (a341 & b_inv341) | (a341 & c341) | (b_inv341 & c341);
  wire s342, sub342, and342, or342;
  wire b_inv342;
  assign b_inv342 = ~b342;
  assign s342  = a342 ^ b342 ^ c342;
  assign sub342 = a342 ^ b_inv342 ^ c342;
  assign and342 = a342 & b342;
  assign or342  = a342 | b342;
  assign c343 = (a342 & b342) | (a342 & c342) | (b342 & c342);
  wire c_sub343;
  assign c_sub343 = (a342 & b_inv342) | (a342 & c342) | (b_inv342 & c342);
  wire s343, sub343, and343, or343;
  wire b_inv343;
  assign b_inv343 = ~b343;
  assign s343  = a343 ^ b343 ^ c343;
  assign sub343 = a343 ^ b_inv343 ^ c343;
  assign and343 = a343 & b343;
  assign or343  = a343 | b343;
  assign c344 = (a343 & b343) | (a343 & c343) | (b343 & c343);
  wire c_sub344;
  assign c_sub344 = (a343 & b_inv343) | (a343 & c343) | (b_inv343 & c343);
  wire s344, sub344, and344, or344;
  wire b_inv344;
  assign b_inv344 = ~b344;
  assign s344  = a344 ^ b344 ^ c344;
  assign sub344 = a344 ^ b_inv344 ^ c344;
  assign and344 = a344 & b344;
  assign or344  = a344 | b344;
  assign c345 = (a344 & b344) | (a344 & c344) | (b344 & c344);
  wire c_sub345;
  assign c_sub345 = (a344 & b_inv344) | (a344 & c344) | (b_inv344 & c344);
  wire s345, sub345, and345, or345;
  wire b_inv345;
  assign b_inv345 = ~b345;
  assign s345  = a345 ^ b345 ^ c345;
  assign sub345 = a345 ^ b_inv345 ^ c345;
  assign and345 = a345 & b345;
  assign or345  = a345 | b345;
  assign c346 = (a345 & b345) | (a345 & c345) | (b345 & c345);
  wire c_sub346;
  assign c_sub346 = (a345 & b_inv345) | (a345 & c345) | (b_inv345 & c345);
  wire s346, sub346, and346, or346;
  wire b_inv346;
  assign b_inv346 = ~b346;
  assign s346  = a346 ^ b346 ^ c346;
  assign sub346 = a346 ^ b_inv346 ^ c346;
  assign and346 = a346 & b346;
  assign or346  = a346 | b346;
  assign c347 = (a346 & b346) | (a346 & c346) | (b346 & c346);
  wire c_sub347;
  assign c_sub347 = (a346 & b_inv346) | (a346 & c346) | (b_inv346 & c346);
  wire s347, sub347, and347, or347;
  wire b_inv347;
  assign b_inv347 = ~b347;
  assign s347  = a347 ^ b347 ^ c347;
  assign sub347 = a347 ^ b_inv347 ^ c347;
  assign and347 = a347 & b347;
  assign or347  = a347 | b347;
  assign c348 = (a347 & b347) | (a347 & c347) | (b347 & c347);
  wire c_sub348;
  assign c_sub348 = (a347 & b_inv347) | (a347 & c347) | (b_inv347 & c347);
  wire s348, sub348, and348, or348;
  wire b_inv348;
  assign b_inv348 = ~b348;
  assign s348  = a348 ^ b348 ^ c348;
  assign sub348 = a348 ^ b_inv348 ^ c348;
  assign and348 = a348 & b348;
  assign or348  = a348 | b348;
  assign c349 = (a348 & b348) | (a348 & c348) | (b348 & c348);
  wire c_sub349;
  assign c_sub349 = (a348 & b_inv348) | (a348 & c348) | (b_inv348 & c348);
  wire s349, sub349, and349, or349;
  wire b_inv349;
  assign b_inv349 = ~b349;
  assign s349  = a349 ^ b349 ^ c349;
  assign sub349 = a349 ^ b_inv349 ^ c349;
  assign and349 = a349 & b349;
  assign or349  = a349 | b349;
  assign c350 = (a349 & b349) | (a349 & c349) | (b349 & c349);
  wire c_sub350;
  assign c_sub350 = (a349 & b_inv349) | (a349 & c349) | (b_inv349 & c349);
  wire s350, sub350, and350, or350;
  wire b_inv350;
  assign b_inv350 = ~b350;
  assign s350  = a350 ^ b350 ^ c350;
  assign sub350 = a350 ^ b_inv350 ^ c350;
  assign and350 = a350 & b350;
  assign or350  = a350 | b350;
  assign c351 = (a350 & b350) | (a350 & c350) | (b350 & c350);
  wire c_sub351;
  assign c_sub351 = (a350 & b_inv350) | (a350 & c350) | (b_inv350 & c350);
  wire s351, sub351, and351, or351;
  wire b_inv351;
  assign b_inv351 = ~b351;
  assign s351  = a351 ^ b351 ^ c351;
  assign sub351 = a351 ^ b_inv351 ^ c351;
  assign and351 = a351 & b351;
  assign or351  = a351 | b351;
  assign c352 = (a351 & b351) | (a351 & c351) | (b351 & c351);
  wire c_sub352;
  assign c_sub352 = (a351 & b_inv351) | (a351 & c351) | (b_inv351 & c351);
  wire s352, sub352, and352, or352;
  wire b_inv352;
  assign b_inv352 = ~b352;
  assign s352  = a352 ^ b352 ^ c352;
  assign sub352 = a352 ^ b_inv352 ^ c352;
  assign and352 = a352 & b352;
  assign or352  = a352 | b352;
  assign c353 = (a352 & b352) | (a352 & c352) | (b352 & c352);
  wire c_sub353;
  assign c_sub353 = (a352 & b_inv352) | (a352 & c352) | (b_inv352 & c352);
  wire s353, sub353, and353, or353;
  wire b_inv353;
  assign b_inv353 = ~b353;
  assign s353  = a353 ^ b353 ^ c353;
  assign sub353 = a353 ^ b_inv353 ^ c353;
  assign and353 = a353 & b353;
  assign or353  = a353 | b353;
  assign c354 = (a353 & b353) | (a353 & c353) | (b353 & c353);
  wire c_sub354;
  assign c_sub354 = (a353 & b_inv353) | (a353 & c353) | (b_inv353 & c353);
  wire s354, sub354, and354, or354;
  wire b_inv354;
  assign b_inv354 = ~b354;
  assign s354  = a354 ^ b354 ^ c354;
  assign sub354 = a354 ^ b_inv354 ^ c354;
  assign and354 = a354 & b354;
  assign or354  = a354 | b354;
  assign c355 = (a354 & b354) | (a354 & c354) | (b354 & c354);
  wire c_sub355;
  assign c_sub355 = (a354 & b_inv354) | (a354 & c354) | (b_inv354 & c354);
  wire s355, sub355, and355, or355;
  wire b_inv355;
  assign b_inv355 = ~b355;
  assign s355  = a355 ^ b355 ^ c355;
  assign sub355 = a355 ^ b_inv355 ^ c355;
  assign and355 = a355 & b355;
  assign or355  = a355 | b355;
  assign c356 = (a355 & b355) | (a355 & c355) | (b355 & c355);
  wire c_sub356;
  assign c_sub356 = (a355 & b_inv355) | (a355 & c355) | (b_inv355 & c355);
  wire s356, sub356, and356, or356;
  wire b_inv356;
  assign b_inv356 = ~b356;
  assign s356  = a356 ^ b356 ^ c356;
  assign sub356 = a356 ^ b_inv356 ^ c356;
  assign and356 = a356 & b356;
  assign or356  = a356 | b356;
  assign c357 = (a356 & b356) | (a356 & c356) | (b356 & c356);
  wire c_sub357;
  assign c_sub357 = (a356 & b_inv356) | (a356 & c356) | (b_inv356 & c356);
  wire s357, sub357, and357, or357;
  wire b_inv357;
  assign b_inv357 = ~b357;
  assign s357  = a357 ^ b357 ^ c357;
  assign sub357 = a357 ^ b_inv357 ^ c357;
  assign and357 = a357 & b357;
  assign or357  = a357 | b357;
  assign c358 = (a357 & b357) | (a357 & c357) | (b357 & c357);
  wire c_sub358;
  assign c_sub358 = (a357 & b_inv357) | (a357 & c357) | (b_inv357 & c357);
  wire s358, sub358, and358, or358;
  wire b_inv358;
  assign b_inv358 = ~b358;
  assign s358  = a358 ^ b358 ^ c358;
  assign sub358 = a358 ^ b_inv358 ^ c358;
  assign and358 = a358 & b358;
  assign or358  = a358 | b358;
  assign c359 = (a358 & b358) | (a358 & c358) | (b358 & c358);
  wire c_sub359;
  assign c_sub359 = (a358 & b_inv358) | (a358 & c358) | (b_inv358 & c358);
  wire s359, sub359, and359, or359;
  wire b_inv359;
  assign b_inv359 = ~b359;
  assign s359  = a359 ^ b359 ^ c359;
  assign sub359 = a359 ^ b_inv359 ^ c359;
  assign and359 = a359 & b359;
  assign or359  = a359 | b359;
  assign c360 = (a359 & b359) | (a359 & c359) | (b359 & c359);
  wire c_sub360;
  assign c_sub360 = (a359 & b_inv359) | (a359 & c359) | (b_inv359 & c359);
  wire s360, sub360, and360, or360;
  wire b_inv360;
  assign b_inv360 = ~b360;
  assign s360  = a360 ^ b360 ^ c360;
  assign sub360 = a360 ^ b_inv360 ^ c360;
  assign and360 = a360 & b360;
  assign or360  = a360 | b360;
  assign c361 = (a360 & b360) | (a360 & c360) | (b360 & c360);
  wire c_sub361;
  assign c_sub361 = (a360 & b_inv360) | (a360 & c360) | (b_inv360 & c360);
  wire s361, sub361, and361, or361;
  wire b_inv361;
  assign b_inv361 = ~b361;
  assign s361  = a361 ^ b361 ^ c361;
  assign sub361 = a361 ^ b_inv361 ^ c361;
  assign and361 = a361 & b361;
  assign or361  = a361 | b361;
  assign c362 = (a361 & b361) | (a361 & c361) | (b361 & c361);
  wire c_sub362;
  assign c_sub362 = (a361 & b_inv361) | (a361 & c361) | (b_inv361 & c361);
  wire s362, sub362, and362, or362;
  wire b_inv362;
  assign b_inv362 = ~b362;
  assign s362  = a362 ^ b362 ^ c362;
  assign sub362 = a362 ^ b_inv362 ^ c362;
  assign and362 = a362 & b362;
  assign or362  = a362 | b362;
  assign c363 = (a362 & b362) | (a362 & c362) | (b362 & c362);
  wire c_sub363;
  assign c_sub363 = (a362 & b_inv362) | (a362 & c362) | (b_inv362 & c362);
  wire s363, sub363, and363, or363;
  wire b_inv363;
  assign b_inv363 = ~b363;
  assign s363  = a363 ^ b363 ^ c363;
  assign sub363 = a363 ^ b_inv363 ^ c363;
  assign and363 = a363 & b363;
  assign or363  = a363 | b363;
  assign c364 = (a363 & b363) | (a363 & c363) | (b363 & c363);
  wire c_sub364;
  assign c_sub364 = (a363 & b_inv363) | (a363 & c363) | (b_inv363 & c363);
  wire s364, sub364, and364, or364;
  wire b_inv364;
  assign b_inv364 = ~b364;
  assign s364  = a364 ^ b364 ^ c364;
  assign sub364 = a364 ^ b_inv364 ^ c364;
  assign and364 = a364 & b364;
  assign or364  = a364 | b364;
  assign c365 = (a364 & b364) | (a364 & c364) | (b364 & c364);
  wire c_sub365;
  assign c_sub365 = (a364 & b_inv364) | (a364 & c364) | (b_inv364 & c364);
  wire s365, sub365, and365, or365;
  wire b_inv365;
  assign b_inv365 = ~b365;
  assign s365  = a365 ^ b365 ^ c365;
  assign sub365 = a365 ^ b_inv365 ^ c365;
  assign and365 = a365 & b365;
  assign or365  = a365 | b365;
  assign c366 = (a365 & b365) | (a365 & c365) | (b365 & c365);
  wire c_sub366;
  assign c_sub366 = (a365 & b_inv365) | (a365 & c365) | (b_inv365 & c365);
  wire s366, sub366, and366, or366;
  wire b_inv366;
  assign b_inv366 = ~b366;
  assign s366  = a366 ^ b366 ^ c366;
  assign sub366 = a366 ^ b_inv366 ^ c366;
  assign and366 = a366 & b366;
  assign or366  = a366 | b366;
  assign c367 = (a366 & b366) | (a366 & c366) | (b366 & c366);
  wire c_sub367;
  assign c_sub367 = (a366 & b_inv366) | (a366 & c366) | (b_inv366 & c366);
  wire s367, sub367, and367, or367;
  wire b_inv367;
  assign b_inv367 = ~b367;
  assign s367  = a367 ^ b367 ^ c367;
  assign sub367 = a367 ^ b_inv367 ^ c367;
  assign and367 = a367 & b367;
  assign or367  = a367 | b367;
  assign c368 = (a367 & b367) | (a367 & c367) | (b367 & c367);
  wire c_sub368;
  assign c_sub368 = (a367 & b_inv367) | (a367 & c367) | (b_inv367 & c367);
  wire s368, sub368, and368, or368;
  wire b_inv368;
  assign b_inv368 = ~b368;
  assign s368  = a368 ^ b368 ^ c368;
  assign sub368 = a368 ^ b_inv368 ^ c368;
  assign and368 = a368 & b368;
  assign or368  = a368 | b368;
  assign c369 = (a368 & b368) | (a368 & c368) | (b368 & c368);
  wire c_sub369;
  assign c_sub369 = (a368 & b_inv368) | (a368 & c368) | (b_inv368 & c368);
  wire s369, sub369, and369, or369;
  wire b_inv369;
  assign b_inv369 = ~b369;
  assign s369  = a369 ^ b369 ^ c369;
  assign sub369 = a369 ^ b_inv369 ^ c369;
  assign and369 = a369 & b369;
  assign or369  = a369 | b369;
  assign c370 = (a369 & b369) | (a369 & c369) | (b369 & c369);
  wire c_sub370;
  assign c_sub370 = (a369 & b_inv369) | (a369 & c369) | (b_inv369 & c369);
  wire s370, sub370, and370, or370;
  wire b_inv370;
  assign b_inv370 = ~b370;
  assign s370  = a370 ^ b370 ^ c370;
  assign sub370 = a370 ^ b_inv370 ^ c370;
  assign and370 = a370 & b370;
  assign or370  = a370 | b370;
  assign c371 = (a370 & b370) | (a370 & c370) | (b370 & c370);
  wire c_sub371;
  assign c_sub371 = (a370 & b_inv370) | (a370 & c370) | (b_inv370 & c370);
  wire s371, sub371, and371, or371;
  wire b_inv371;
  assign b_inv371 = ~b371;
  assign s371  = a371 ^ b371 ^ c371;
  assign sub371 = a371 ^ b_inv371 ^ c371;
  assign and371 = a371 & b371;
  assign or371  = a371 | b371;
  assign c372 = (a371 & b371) | (a371 & c371) | (b371 & c371);
  wire c_sub372;
  assign c_sub372 = (a371 & b_inv371) | (a371 & c371) | (b_inv371 & c371);
  wire s372, sub372, and372, or372;
  wire b_inv372;
  assign b_inv372 = ~b372;
  assign s372  = a372 ^ b372 ^ c372;
  assign sub372 = a372 ^ b_inv372 ^ c372;
  assign and372 = a372 & b372;
  assign or372  = a372 | b372;
  assign c373 = (a372 & b372) | (a372 & c372) | (b372 & c372);
  wire c_sub373;
  assign c_sub373 = (a372 & b_inv372) | (a372 & c372) | (b_inv372 & c372);
  wire s373, sub373, and373, or373;
  wire b_inv373;
  assign b_inv373 = ~b373;
  assign s373  = a373 ^ b373 ^ c373;
  assign sub373 = a373 ^ b_inv373 ^ c373;
  assign and373 = a373 & b373;
  assign or373  = a373 | b373;
  assign c374 = (a373 & b373) | (a373 & c373) | (b373 & c373);
  wire c_sub374;
  assign c_sub374 = (a373 & b_inv373) | (a373 & c373) | (b_inv373 & c373);
  wire s374, sub374, and374, or374;
  wire b_inv374;
  assign b_inv374 = ~b374;
  assign s374  = a374 ^ b374 ^ c374;
  assign sub374 = a374 ^ b_inv374 ^ c374;
  assign and374 = a374 & b374;
  assign or374  = a374 | b374;
  assign c375 = (a374 & b374) | (a374 & c374) | (b374 & c374);
  wire c_sub375;
  assign c_sub375 = (a374 & b_inv374) | (a374 & c374) | (b_inv374 & c374);
  wire s375, sub375, and375, or375;
  wire b_inv375;
  assign b_inv375 = ~b375;
  assign s375  = a375 ^ b375 ^ c375;
  assign sub375 = a375 ^ b_inv375 ^ c375;
  assign and375 = a375 & b375;
  assign or375  = a375 | b375;
  assign c376 = (a375 & b375) | (a375 & c375) | (b375 & c375);
  wire c_sub376;
  assign c_sub376 = (a375 & b_inv375) | (a375 & c375) | (b_inv375 & c375);
  wire s376, sub376, and376, or376;
  wire b_inv376;
  assign b_inv376 = ~b376;
  assign s376  = a376 ^ b376 ^ c376;
  assign sub376 = a376 ^ b_inv376 ^ c376;
  assign and376 = a376 & b376;
  assign or376  = a376 | b376;
  assign c377 = (a376 & b376) | (a376 & c376) | (b376 & c376);
  wire c_sub377;
  assign c_sub377 = (a376 & b_inv376) | (a376 & c376) | (b_inv376 & c376);
  wire s377, sub377, and377, or377;
  wire b_inv377;
  assign b_inv377 = ~b377;
  assign s377  = a377 ^ b377 ^ c377;
  assign sub377 = a377 ^ b_inv377 ^ c377;
  assign and377 = a377 & b377;
  assign or377  = a377 | b377;
  assign c378 = (a377 & b377) | (a377 & c377) | (b377 & c377);
  wire c_sub378;
  assign c_sub378 = (a377 & b_inv377) | (a377 & c377) | (b_inv377 & c377);
  wire s378, sub378, and378, or378;
  wire b_inv378;
  assign b_inv378 = ~b378;
  assign s378  = a378 ^ b378 ^ c378;
  assign sub378 = a378 ^ b_inv378 ^ c378;
  assign and378 = a378 & b378;
  assign or378  = a378 | b378;
  assign c379 = (a378 & b378) | (a378 & c378) | (b378 & c378);
  wire c_sub379;
  assign c_sub379 = (a378 & b_inv378) | (a378 & c378) | (b_inv378 & c378);
  wire s379, sub379, and379, or379;
  wire b_inv379;
  assign b_inv379 = ~b379;
  assign s379  = a379 ^ b379 ^ c379;
  assign sub379 = a379 ^ b_inv379 ^ c379;
  assign and379 = a379 & b379;
  assign or379  = a379 | b379;
  assign c380 = (a379 & b379) | (a379 & c379) | (b379 & c379);
  wire c_sub380;
  assign c_sub380 = (a379 & b_inv379) | (a379 & c379) | (b_inv379 & c379);
  wire s380, sub380, and380, or380;
  wire b_inv380;
  assign b_inv380 = ~b380;
  assign s380  = a380 ^ b380 ^ c380;
  assign sub380 = a380 ^ b_inv380 ^ c380;
  assign and380 = a380 & b380;
  assign or380  = a380 | b380;
  assign c381 = (a380 & b380) | (a380 & c380) | (b380 & c380);
  wire c_sub381;
  assign c_sub381 = (a380 & b_inv380) | (a380 & c380) | (b_inv380 & c380);
  wire s381, sub381, and381, or381;
  wire b_inv381;
  assign b_inv381 = ~b381;
  assign s381  = a381 ^ b381 ^ c381;
  assign sub381 = a381 ^ b_inv381 ^ c381;
  assign and381 = a381 & b381;
  assign or381  = a381 | b381;
  assign c382 = (a381 & b381) | (a381 & c381) | (b381 & c381);
  wire c_sub382;
  assign c_sub382 = (a381 & b_inv381) | (a381 & c381) | (b_inv381 & c381);
  wire s382, sub382, and382, or382;
  wire b_inv382;
  assign b_inv382 = ~b382;
  assign s382  = a382 ^ b382 ^ c382;
  assign sub382 = a382 ^ b_inv382 ^ c382;
  assign and382 = a382 & b382;
  assign or382  = a382 | b382;
  assign c383 = (a382 & b382) | (a382 & c382) | (b382 & c382);
  wire c_sub383;
  assign c_sub383 = (a382 & b_inv382) | (a382 & c382) | (b_inv382 & c382);
  wire s383, sub383, and383, or383;
  wire b_inv383;
  assign b_inv383 = ~b383;
  assign s383  = a383 ^ b383 ^ c383;
  assign sub383 = a383 ^ b_inv383 ^ c383;
  assign and383 = a383 & b383;
  assign or383  = a383 | b383;
  assign c384 = (a383 & b383) | (a383 & c383) | (b383 & c383);
  wire c_sub384;
  assign c_sub384 = (a383 & b_inv383) | (a383 & c383) | (b_inv383 & c383);
  wire s384, sub384, and384, or384;
  wire b_inv384;
  assign b_inv384 = ~b384;
  assign s384  = a384 ^ b384 ^ c384;
  assign sub384 = a384 ^ b_inv384 ^ c384;
  assign and384 = a384 & b384;
  assign or384  = a384 | b384;
  assign c385 = (a384 & b384) | (a384 & c384) | (b384 & c384);
  wire c_sub385;
  assign c_sub385 = (a384 & b_inv384) | (a384 & c384) | (b_inv384 & c384);
  wire s385, sub385, and385, or385;
  wire b_inv385;
  assign b_inv385 = ~b385;
  assign s385  = a385 ^ b385 ^ c385;
  assign sub385 = a385 ^ b_inv385 ^ c385;
  assign and385 = a385 & b385;
  assign or385  = a385 | b385;
  assign c386 = (a385 & b385) | (a385 & c385) | (b385 & c385);
  wire c_sub386;
  assign c_sub386 = (a385 & b_inv385) | (a385 & c385) | (b_inv385 & c385);
  wire s386, sub386, and386, or386;
  wire b_inv386;
  assign b_inv386 = ~b386;
  assign s386  = a386 ^ b386 ^ c386;
  assign sub386 = a386 ^ b_inv386 ^ c386;
  assign and386 = a386 & b386;
  assign or386  = a386 | b386;
  assign c387 = (a386 & b386) | (a386 & c386) | (b386 & c386);
  wire c_sub387;
  assign c_sub387 = (a386 & b_inv386) | (a386 & c386) | (b_inv386 & c386);
  wire s387, sub387, and387, or387;
  wire b_inv387;
  assign b_inv387 = ~b387;
  assign s387  = a387 ^ b387 ^ c387;
  assign sub387 = a387 ^ b_inv387 ^ c387;
  assign and387 = a387 & b387;
  assign or387  = a387 | b387;
  assign c388 = (a387 & b387) | (a387 & c387) | (b387 & c387);
  wire c_sub388;
  assign c_sub388 = (a387 & b_inv387) | (a387 & c387) | (b_inv387 & c387);
  wire s388, sub388, and388, or388;
  wire b_inv388;
  assign b_inv388 = ~b388;
  assign s388  = a388 ^ b388 ^ c388;
  assign sub388 = a388 ^ b_inv388 ^ c388;
  assign and388 = a388 & b388;
  assign or388  = a388 | b388;
  assign c389 = (a388 & b388) | (a388 & c388) | (b388 & c388);
  wire c_sub389;
  assign c_sub389 = (a388 & b_inv388) | (a388 & c388) | (b_inv388 & c388);
  wire s389, sub389, and389, or389;
  wire b_inv389;
  assign b_inv389 = ~b389;
  assign s389  = a389 ^ b389 ^ c389;
  assign sub389 = a389 ^ b_inv389 ^ c389;
  assign and389 = a389 & b389;
  assign or389  = a389 | b389;
  assign c390 = (a389 & b389) | (a389 & c389) | (b389 & c389);
  wire c_sub390;
  assign c_sub390 = (a389 & b_inv389) | (a389 & c389) | (b_inv389 & c389);
  wire s390, sub390, and390, or390;
  wire b_inv390;
  assign b_inv390 = ~b390;
  assign s390  = a390 ^ b390 ^ c390;
  assign sub390 = a390 ^ b_inv390 ^ c390;
  assign and390 = a390 & b390;
  assign or390  = a390 | b390;
  assign c391 = (a390 & b390) | (a390 & c390) | (b390 & c390);
  wire c_sub391;
  assign c_sub391 = (a390 & b_inv390) | (a390 & c390) | (b_inv390 & c390);
  wire s391, sub391, and391, or391;
  wire b_inv391;
  assign b_inv391 = ~b391;
  assign s391  = a391 ^ b391 ^ c391;
  assign sub391 = a391 ^ b_inv391 ^ c391;
  assign and391 = a391 & b391;
  assign or391  = a391 | b391;
  assign c392 = (a391 & b391) | (a391 & c391) | (b391 & c391);
  wire c_sub392;
  assign c_sub392 = (a391 & b_inv391) | (a391 & c391) | (b_inv391 & c391);
  wire s392, sub392, and392, or392;
  wire b_inv392;
  assign b_inv392 = ~b392;
  assign s392  = a392 ^ b392 ^ c392;
  assign sub392 = a392 ^ b_inv392 ^ c392;
  assign and392 = a392 & b392;
  assign or392  = a392 | b392;
  assign c393 = (a392 & b392) | (a392 & c392) | (b392 & c392);
  wire c_sub393;
  assign c_sub393 = (a392 & b_inv392) | (a392 & c392) | (b_inv392 & c392);
  wire s393, sub393, and393, or393;
  wire b_inv393;
  assign b_inv393 = ~b393;
  assign s393  = a393 ^ b393 ^ c393;
  assign sub393 = a393 ^ b_inv393 ^ c393;
  assign and393 = a393 & b393;
  assign or393  = a393 | b393;
  assign c394 = (a393 & b393) | (a393 & c393) | (b393 & c393);
  wire c_sub394;
  assign c_sub394 = (a393 & b_inv393) | (a393 & c393) | (b_inv393 & c393);
  wire s394, sub394, and394, or394;
  wire b_inv394;
  assign b_inv394 = ~b394;
  assign s394  = a394 ^ b394 ^ c394;
  assign sub394 = a394 ^ b_inv394 ^ c394;
  assign and394 = a394 & b394;
  assign or394  = a394 | b394;
  assign c395 = (a394 & b394) | (a394 & c394) | (b394 & c394);
  wire c_sub395;
  assign c_sub395 = (a394 & b_inv394) | (a394 & c394) | (b_inv394 & c394);
  wire s395, sub395, and395, or395;
  wire b_inv395;
  assign b_inv395 = ~b395;
  assign s395  = a395 ^ b395 ^ c395;
  assign sub395 = a395 ^ b_inv395 ^ c395;
  assign and395 = a395 & b395;
  assign or395  = a395 | b395;
  assign c396 = (a395 & b395) | (a395 & c395) | (b395 & c395);
  wire c_sub396;
  assign c_sub396 = (a395 & b_inv395) | (a395 & c395) | (b_inv395 & c395);
  wire s396, sub396, and396, or396;
  wire b_inv396;
  assign b_inv396 = ~b396;
  assign s396  = a396 ^ b396 ^ c396;
  assign sub396 = a396 ^ b_inv396 ^ c396;
  assign and396 = a396 & b396;
  assign or396  = a396 | b396;
  assign c397 = (a396 & b396) | (a396 & c396) | (b396 & c396);
  wire c_sub397;
  assign c_sub397 = (a396 & b_inv396) | (a396 & c396) | (b_inv396 & c396);
  wire s397, sub397, and397, or397;
  wire b_inv397;
  assign b_inv397 = ~b397;
  assign s397  = a397 ^ b397 ^ c397;
  assign sub397 = a397 ^ b_inv397 ^ c397;
  assign and397 = a397 & b397;
  assign or397  = a397 | b397;
  assign c398 = (a397 & b397) | (a397 & c397) | (b397 & c397);
  wire c_sub398;
  assign c_sub398 = (a397 & b_inv397) | (a397 & c397) | (b_inv397 & c397);
  wire s398, sub398, and398, or398;
  wire b_inv398;
  assign b_inv398 = ~b398;
  assign s398  = a398 ^ b398 ^ c398;
  assign sub398 = a398 ^ b_inv398 ^ c398;
  assign and398 = a398 & b398;
  assign or398  = a398 | b398;
  assign c399 = (a398 & b398) | (a398 & c398) | (b398 & c398);
  wire c_sub399;
  assign c_sub399 = (a398 & b_inv398) | (a398 & c398) | (b_inv398 & c398);
  wire s399, sub399, and399, or399;
  wire b_inv399;
  assign b_inv399 = ~b399;
  assign s399  = a399 ^ b399 ^ c399;
  assign sub399 = a399 ^ b_inv399 ^ c399;
  assign and399 = a399 & b399;
  assign or399  = a399 | b399;
  assign c400 = (a399 & b399) | (a399 & c399) | (b399 & c399);
  wire c_sub400;
  assign c_sub400 = (a399 & b_inv399) | (a399 & c399) | (b_inv399 & c399);
  wire s400, sub400, and400, or400;
  wire b_inv400;
  assign b_inv400 = ~b400;
  assign s400  = a400 ^ b400 ^ c400;
  assign sub400 = a400 ^ b_inv400 ^ c400;
  assign and400 = a400 & b400;
  assign or400  = a400 | b400;
  assign c401 = (a400 & b400) | (a400 & c400) | (b400 & c400);
  wire c_sub401;
  assign c_sub401 = (a400 & b_inv400) | (a400 & c400) | (b_inv400 & c400);
  wire s401, sub401, and401, or401;
  wire b_inv401;
  assign b_inv401 = ~b401;
  assign s401  = a401 ^ b401 ^ c401;
  assign sub401 = a401 ^ b_inv401 ^ c401;
  assign and401 = a401 & b401;
  assign or401  = a401 | b401;
  assign c402 = (a401 & b401) | (a401 & c401) | (b401 & c401);
  wire c_sub402;
  assign c_sub402 = (a401 & b_inv401) | (a401 & c401) | (b_inv401 & c401);
  wire s402, sub402, and402, or402;
  wire b_inv402;
  assign b_inv402 = ~b402;
  assign s402  = a402 ^ b402 ^ c402;
  assign sub402 = a402 ^ b_inv402 ^ c402;
  assign and402 = a402 & b402;
  assign or402  = a402 | b402;
  assign c403 = (a402 & b402) | (a402 & c402) | (b402 & c402);
  wire c_sub403;
  assign c_sub403 = (a402 & b_inv402) | (a402 & c402) | (b_inv402 & c402);
  wire s403, sub403, and403, or403;
  wire b_inv403;
  assign b_inv403 = ~b403;
  assign s403  = a403 ^ b403 ^ c403;
  assign sub403 = a403 ^ b_inv403 ^ c403;
  assign and403 = a403 & b403;
  assign or403  = a403 | b403;
  assign c404 = (a403 & b403) | (a403 & c403) | (b403 & c403);
  wire c_sub404;
  assign c_sub404 = (a403 & b_inv403) | (a403 & c403) | (b_inv403 & c403);
  wire s404, sub404, and404, or404;
  wire b_inv404;
  assign b_inv404 = ~b404;
  assign s404  = a404 ^ b404 ^ c404;
  assign sub404 = a404 ^ b_inv404 ^ c404;
  assign and404 = a404 & b404;
  assign or404  = a404 | b404;
  assign c405 = (a404 & b404) | (a404 & c404) | (b404 & c404);
  wire c_sub405;
  assign c_sub405 = (a404 & b_inv404) | (a404 & c404) | (b_inv404 & c404);
  wire s405, sub405, and405, or405;
  wire b_inv405;
  assign b_inv405 = ~b405;
  assign s405  = a405 ^ b405 ^ c405;
  assign sub405 = a405 ^ b_inv405 ^ c405;
  assign and405 = a405 & b405;
  assign or405  = a405 | b405;
  assign c406 = (a405 & b405) | (a405 & c405) | (b405 & c405);
  wire c_sub406;
  assign c_sub406 = (a405 & b_inv405) | (a405 & c405) | (b_inv405 & c405);
  wire s406, sub406, and406, or406;
  wire b_inv406;
  assign b_inv406 = ~b406;
  assign s406  = a406 ^ b406 ^ c406;
  assign sub406 = a406 ^ b_inv406 ^ c406;
  assign and406 = a406 & b406;
  assign or406  = a406 | b406;
  assign c407 = (a406 & b406) | (a406 & c406) | (b406 & c406);
  wire c_sub407;
  assign c_sub407 = (a406 & b_inv406) | (a406 & c406) | (b_inv406 & c406);
  wire s407, sub407, and407, or407;
  wire b_inv407;
  assign b_inv407 = ~b407;
  assign s407  = a407 ^ b407 ^ c407;
  assign sub407 = a407 ^ b_inv407 ^ c407;
  assign and407 = a407 & b407;
  assign or407  = a407 | b407;
  assign c408 = (a407 & b407) | (a407 & c407) | (b407 & c407);
  wire c_sub408;
  assign c_sub408 = (a407 & b_inv407) | (a407 & c407) | (b_inv407 & c407);
  wire s408, sub408, and408, or408;
  wire b_inv408;
  assign b_inv408 = ~b408;
  assign s408  = a408 ^ b408 ^ c408;
  assign sub408 = a408 ^ b_inv408 ^ c408;
  assign and408 = a408 & b408;
  assign or408  = a408 | b408;
  assign c409 = (a408 & b408) | (a408 & c408) | (b408 & c408);
  wire c_sub409;
  assign c_sub409 = (a408 & b_inv408) | (a408 & c408) | (b_inv408 & c408);
  wire s409, sub409, and409, or409;
  wire b_inv409;
  assign b_inv409 = ~b409;
  assign s409  = a409 ^ b409 ^ c409;
  assign sub409 = a409 ^ b_inv409 ^ c409;
  assign and409 = a409 & b409;
  assign or409  = a409 | b409;
  assign c410 = (a409 & b409) | (a409 & c409) | (b409 & c409);
  wire c_sub410;
  assign c_sub410 = (a409 & b_inv409) | (a409 & c409) | (b_inv409 & c409);
  wire s410, sub410, and410, or410;
  wire b_inv410;
  assign b_inv410 = ~b410;
  assign s410  = a410 ^ b410 ^ c410;
  assign sub410 = a410 ^ b_inv410 ^ c410;
  assign and410 = a410 & b410;
  assign or410  = a410 | b410;
  assign c411 = (a410 & b410) | (a410 & c410) | (b410 & c410);
  wire c_sub411;
  assign c_sub411 = (a410 & b_inv410) | (a410 & c410) | (b_inv410 & c410);
  wire s411, sub411, and411, or411;
  wire b_inv411;
  assign b_inv411 = ~b411;
  assign s411  = a411 ^ b411 ^ c411;
  assign sub411 = a411 ^ b_inv411 ^ c411;
  assign and411 = a411 & b411;
  assign or411  = a411 | b411;
  assign c412 = (a411 & b411) | (a411 & c411) | (b411 & c411);
  wire c_sub412;
  assign c_sub412 = (a411 & b_inv411) | (a411 & c411) | (b_inv411 & c411);
  wire s412, sub412, and412, or412;
  wire b_inv412;
  assign b_inv412 = ~b412;
  assign s412  = a412 ^ b412 ^ c412;
  assign sub412 = a412 ^ b_inv412 ^ c412;
  assign and412 = a412 & b412;
  assign or412  = a412 | b412;
  assign c413 = (a412 & b412) | (a412 & c412) | (b412 & c412);
  wire c_sub413;
  assign c_sub413 = (a412 & b_inv412) | (a412 & c412) | (b_inv412 & c412);
  wire s413, sub413, and413, or413;
  wire b_inv413;
  assign b_inv413 = ~b413;
  assign s413  = a413 ^ b413 ^ c413;
  assign sub413 = a413 ^ b_inv413 ^ c413;
  assign and413 = a413 & b413;
  assign or413  = a413 | b413;
  assign c414 = (a413 & b413) | (a413 & c413) | (b413 & c413);
  wire c_sub414;
  assign c_sub414 = (a413 & b_inv413) | (a413 & c413) | (b_inv413 & c413);
  wire s414, sub414, and414, or414;
  wire b_inv414;
  assign b_inv414 = ~b414;
  assign s414  = a414 ^ b414 ^ c414;
  assign sub414 = a414 ^ b_inv414 ^ c414;
  assign and414 = a414 & b414;
  assign or414  = a414 | b414;
  assign c415 = (a414 & b414) | (a414 & c414) | (b414 & c414);
  wire c_sub415;
  assign c_sub415 = (a414 & b_inv414) | (a414 & c414) | (b_inv414 & c414);
  wire s415, sub415, and415, or415;
  wire b_inv415;
  assign b_inv415 = ~b415;
  assign s415  = a415 ^ b415 ^ c415;
  assign sub415 = a415 ^ b_inv415 ^ c415;
  assign and415 = a415 & b415;
  assign or415  = a415 | b415;
  assign c416 = (a415 & b415) | (a415 & c415) | (b415 & c415);
  wire c_sub416;
  assign c_sub416 = (a415 & b_inv415) | (a415 & c415) | (b_inv415 & c415);
  wire s416, sub416, and416, or416;
  wire b_inv416;
  assign b_inv416 = ~b416;
  assign s416  = a416 ^ b416 ^ c416;
  assign sub416 = a416 ^ b_inv416 ^ c416;
  assign and416 = a416 & b416;
  assign or416  = a416 | b416;
  assign c417 = (a416 & b416) | (a416 & c416) | (b416 & c416);
  wire c_sub417;
  assign c_sub417 = (a416 & b_inv416) | (a416 & c416) | (b_inv416 & c416);
  wire s417, sub417, and417, or417;
  wire b_inv417;
  assign b_inv417 = ~b417;
  assign s417  = a417 ^ b417 ^ c417;
  assign sub417 = a417 ^ b_inv417 ^ c417;
  assign and417 = a417 & b417;
  assign or417  = a417 | b417;
  assign c418 = (a417 & b417) | (a417 & c417) | (b417 & c417);
  wire c_sub418;
  assign c_sub418 = (a417 & b_inv417) | (a417 & c417) | (b_inv417 & c417);
  wire s418, sub418, and418, or418;
  wire b_inv418;
  assign b_inv418 = ~b418;
  assign s418  = a418 ^ b418 ^ c418;
  assign sub418 = a418 ^ b_inv418 ^ c418;
  assign and418 = a418 & b418;
  assign or418  = a418 | b418;
  assign c419 = (a418 & b418) | (a418 & c418) | (b418 & c418);
  wire c_sub419;
  assign c_sub419 = (a418 & b_inv418) | (a418 & c418) | (b_inv418 & c418);
  wire s419, sub419, and419, or419;
  wire b_inv419;
  assign b_inv419 = ~b419;
  assign s419  = a419 ^ b419 ^ c419;
  assign sub419 = a419 ^ b_inv419 ^ c419;
  assign and419 = a419 & b419;
  assign or419  = a419 | b419;
  assign c420 = (a419 & b419) | (a419 & c419) | (b419 & c419);
  wire c_sub420;
  assign c_sub420 = (a419 & b_inv419) | (a419 & c419) | (b_inv419 & c419);
  wire s420, sub420, and420, or420;
  wire b_inv420;
  assign b_inv420 = ~b420;
  assign s420  = a420 ^ b420 ^ c420;
  assign sub420 = a420 ^ b_inv420 ^ c420;
  assign and420 = a420 & b420;
  assign or420  = a420 | b420;
  assign c421 = (a420 & b420) | (a420 & c420) | (b420 & c420);
  wire c_sub421;
  assign c_sub421 = (a420 & b_inv420) | (a420 & c420) | (b_inv420 & c420);
  wire s421, sub421, and421, or421;
  wire b_inv421;
  assign b_inv421 = ~b421;
  assign s421  = a421 ^ b421 ^ c421;
  assign sub421 = a421 ^ b_inv421 ^ c421;
  assign and421 = a421 & b421;
  assign or421  = a421 | b421;
  assign c422 = (a421 & b421) | (a421 & c421) | (b421 & c421);
  wire c_sub422;
  assign c_sub422 = (a421 & b_inv421) | (a421 & c421) | (b_inv421 & c421);
  wire s422, sub422, and422, or422;
  wire b_inv422;
  assign b_inv422 = ~b422;
  assign s422  = a422 ^ b422 ^ c422;
  assign sub422 = a422 ^ b_inv422 ^ c422;
  assign and422 = a422 & b422;
  assign or422  = a422 | b422;
  assign c423 = (a422 & b422) | (a422 & c422) | (b422 & c422);
  wire c_sub423;
  assign c_sub423 = (a422 & b_inv422) | (a422 & c422) | (b_inv422 & c422);
  wire s423, sub423, and423, or423;
  wire b_inv423;
  assign b_inv423 = ~b423;
  assign s423  = a423 ^ b423 ^ c423;
  assign sub423 = a423 ^ b_inv423 ^ c423;
  assign and423 = a423 & b423;
  assign or423  = a423 | b423;
  assign c424 = (a423 & b423) | (a423 & c423) | (b423 & c423);
  wire c_sub424;
  assign c_sub424 = (a423 & b_inv423) | (a423 & c423) | (b_inv423 & c423);
  wire s424, sub424, and424, or424;
  wire b_inv424;
  assign b_inv424 = ~b424;
  assign s424  = a424 ^ b424 ^ c424;
  assign sub424 = a424 ^ b_inv424 ^ c424;
  assign and424 = a424 & b424;
  assign or424  = a424 | b424;
  assign c425 = (a424 & b424) | (a424 & c424) | (b424 & c424);
  wire c_sub425;
  assign c_sub425 = (a424 & b_inv424) | (a424 & c424) | (b_inv424 & c424);
  wire s425, sub425, and425, or425;
  wire b_inv425;
  assign b_inv425 = ~b425;
  assign s425  = a425 ^ b425 ^ c425;
  assign sub425 = a425 ^ b_inv425 ^ c425;
  assign and425 = a425 & b425;
  assign or425  = a425 | b425;
  assign c426 = (a425 & b425) | (a425 & c425) | (b425 & c425);
  wire c_sub426;
  assign c_sub426 = (a425 & b_inv425) | (a425 & c425) | (b_inv425 & c425);
  wire s426, sub426, and426, or426;
  wire b_inv426;
  assign b_inv426 = ~b426;
  assign s426  = a426 ^ b426 ^ c426;
  assign sub426 = a426 ^ b_inv426 ^ c426;
  assign and426 = a426 & b426;
  assign or426  = a426 | b426;
  assign c427 = (a426 & b426) | (a426 & c426) | (b426 & c426);
  wire c_sub427;
  assign c_sub427 = (a426 & b_inv426) | (a426 & c426) | (b_inv426 & c426);
  wire s427, sub427, and427, or427;
  wire b_inv427;
  assign b_inv427 = ~b427;
  assign s427  = a427 ^ b427 ^ c427;
  assign sub427 = a427 ^ b_inv427 ^ c427;
  assign and427 = a427 & b427;
  assign or427  = a427 | b427;
  assign c428 = (a427 & b427) | (a427 & c427) | (b427 & c427);
  wire c_sub428;
  assign c_sub428 = (a427 & b_inv427) | (a427 & c427) | (b_inv427 & c427);
  wire s428, sub428, and428, or428;
  wire b_inv428;
  assign b_inv428 = ~b428;
  assign s428  = a428 ^ b428 ^ c428;
  assign sub428 = a428 ^ b_inv428 ^ c428;
  assign and428 = a428 & b428;
  assign or428  = a428 | b428;
  assign c429 = (a428 & b428) | (a428 & c428) | (b428 & c428);
  wire c_sub429;
  assign c_sub429 = (a428 & b_inv428) | (a428 & c428) | (b_inv428 & c428);
  wire s429, sub429, and429, or429;
  wire b_inv429;
  assign b_inv429 = ~b429;
  assign s429  = a429 ^ b429 ^ c429;
  assign sub429 = a429 ^ b_inv429 ^ c429;
  assign and429 = a429 & b429;
  assign or429  = a429 | b429;
  assign c430 = (a429 & b429) | (a429 & c429) | (b429 & c429);
  wire c_sub430;
  assign c_sub430 = (a429 & b_inv429) | (a429 & c429) | (b_inv429 & c429);
  wire s430, sub430, and430, or430;
  wire b_inv430;
  assign b_inv430 = ~b430;
  assign s430  = a430 ^ b430 ^ c430;
  assign sub430 = a430 ^ b_inv430 ^ c430;
  assign and430 = a430 & b430;
  assign or430  = a430 | b430;
  assign c431 = (a430 & b430) | (a430 & c430) | (b430 & c430);
  wire c_sub431;
  assign c_sub431 = (a430 & b_inv430) | (a430 & c430) | (b_inv430 & c430);
  wire s431, sub431, and431, or431;
  wire b_inv431;
  assign b_inv431 = ~b431;
  assign s431  = a431 ^ b431 ^ c431;
  assign sub431 = a431 ^ b_inv431 ^ c431;
  assign and431 = a431 & b431;
  assign or431  = a431 | b431;
  assign c432 = (a431 & b431) | (a431 & c431) | (b431 & c431);
  wire c_sub432;
  assign c_sub432 = (a431 & b_inv431) | (a431 & c431) | (b_inv431 & c431);
  wire s432, sub432, and432, or432;
  wire b_inv432;
  assign b_inv432 = ~b432;
  assign s432  = a432 ^ b432 ^ c432;
  assign sub432 = a432 ^ b_inv432 ^ c432;
  assign and432 = a432 & b432;
  assign or432  = a432 | b432;
  assign c433 = (a432 & b432) | (a432 & c432) | (b432 & c432);
  wire c_sub433;
  assign c_sub433 = (a432 & b_inv432) | (a432 & c432) | (b_inv432 & c432);
  wire s433, sub433, and433, or433;
  wire b_inv433;
  assign b_inv433 = ~b433;
  assign s433  = a433 ^ b433 ^ c433;
  assign sub433 = a433 ^ b_inv433 ^ c433;
  assign and433 = a433 & b433;
  assign or433  = a433 | b433;
  assign c434 = (a433 & b433) | (a433 & c433) | (b433 & c433);
  wire c_sub434;
  assign c_sub434 = (a433 & b_inv433) | (a433 & c433) | (b_inv433 & c433);
  wire s434, sub434, and434, or434;
  wire b_inv434;
  assign b_inv434 = ~b434;
  assign s434  = a434 ^ b434 ^ c434;
  assign sub434 = a434 ^ b_inv434 ^ c434;
  assign and434 = a434 & b434;
  assign or434  = a434 | b434;
  assign c435 = (a434 & b434) | (a434 & c434) | (b434 & c434);
  wire c_sub435;
  assign c_sub435 = (a434 & b_inv434) | (a434 & c434) | (b_inv434 & c434);
  wire s435, sub435, and435, or435;
  wire b_inv435;
  assign b_inv435 = ~b435;
  assign s435  = a435 ^ b435 ^ c435;
  assign sub435 = a435 ^ b_inv435 ^ c435;
  assign and435 = a435 & b435;
  assign or435  = a435 | b435;
  assign c436 = (a435 & b435) | (a435 & c435) | (b435 & c435);
  wire c_sub436;
  assign c_sub436 = (a435 & b_inv435) | (a435 & c435) | (b_inv435 & c435);
  wire s436, sub436, and436, or436;
  wire b_inv436;
  assign b_inv436 = ~b436;
  assign s436  = a436 ^ b436 ^ c436;
  assign sub436 = a436 ^ b_inv436 ^ c436;
  assign and436 = a436 & b436;
  assign or436  = a436 | b436;
  assign c437 = (a436 & b436) | (a436 & c436) | (b436 & c436);
  wire c_sub437;
  assign c_sub437 = (a436 & b_inv436) | (a436 & c436) | (b_inv436 & c436);
  wire s437, sub437, and437, or437;
  wire b_inv437;
  assign b_inv437 = ~b437;
  assign s437  = a437 ^ b437 ^ c437;
  assign sub437 = a437 ^ b_inv437 ^ c437;
  assign and437 = a437 & b437;
  assign or437  = a437 | b437;
  assign c438 = (a437 & b437) | (a437 & c437) | (b437 & c437);
  wire c_sub438;
  assign c_sub438 = (a437 & b_inv437) | (a437 & c437) | (b_inv437 & c437);
  wire s438, sub438, and438, or438;
  wire b_inv438;
  assign b_inv438 = ~b438;
  assign s438  = a438 ^ b438 ^ c438;
  assign sub438 = a438 ^ b_inv438 ^ c438;
  assign and438 = a438 & b438;
  assign or438  = a438 | b438;
  assign c439 = (a438 & b438) | (a438 & c438) | (b438 & c438);
  wire c_sub439;
  assign c_sub439 = (a438 & b_inv438) | (a438 & c438) | (b_inv438 & c438);
  wire s439, sub439, and439, or439;
  wire b_inv439;
  assign b_inv439 = ~b439;
  assign s439  = a439 ^ b439 ^ c439;
  assign sub439 = a439 ^ b_inv439 ^ c439;
  assign and439 = a439 & b439;
  assign or439  = a439 | b439;
  assign c440 = (a439 & b439) | (a439 & c439) | (b439 & c439);
  wire c_sub440;
  assign c_sub440 = (a439 & b_inv439) | (a439 & c439) | (b_inv439 & c439);
  wire s440, sub440, and440, or440;
  wire b_inv440;
  assign b_inv440 = ~b440;
  assign s440  = a440 ^ b440 ^ c440;
  assign sub440 = a440 ^ b_inv440 ^ c440;
  assign and440 = a440 & b440;
  assign or440  = a440 | b440;
  assign c441 = (a440 & b440) | (a440 & c440) | (b440 & c440);
  wire c_sub441;
  assign c_sub441 = (a440 & b_inv440) | (a440 & c440) | (b_inv440 & c440);
  wire s441, sub441, and441, or441;
  wire b_inv441;
  assign b_inv441 = ~b441;
  assign s441  = a441 ^ b441 ^ c441;
  assign sub441 = a441 ^ b_inv441 ^ c441;
  assign and441 = a441 & b441;
  assign or441  = a441 | b441;
  assign c442 = (a441 & b441) | (a441 & c441) | (b441 & c441);
  wire c_sub442;
  assign c_sub442 = (a441 & b_inv441) | (a441 & c441) | (b_inv441 & c441);
  wire s442, sub442, and442, or442;
  wire b_inv442;
  assign b_inv442 = ~b442;
  assign s442  = a442 ^ b442 ^ c442;
  assign sub442 = a442 ^ b_inv442 ^ c442;
  assign and442 = a442 & b442;
  assign or442  = a442 | b442;
  assign c443 = (a442 & b442) | (a442 & c442) | (b442 & c442);
  wire c_sub443;
  assign c_sub443 = (a442 & b_inv442) | (a442 & c442) | (b_inv442 & c442);
  wire s443, sub443, and443, or443;
  wire b_inv443;
  assign b_inv443 = ~b443;
  assign s443  = a443 ^ b443 ^ c443;
  assign sub443 = a443 ^ b_inv443 ^ c443;
  assign and443 = a443 & b443;
  assign or443  = a443 | b443;
  assign c444 = (a443 & b443) | (a443 & c443) | (b443 & c443);
  wire c_sub444;
  assign c_sub444 = (a443 & b_inv443) | (a443 & c443) | (b_inv443 & c443);
  wire s444, sub444, and444, or444;
  wire b_inv444;
  assign b_inv444 = ~b444;
  assign s444  = a444 ^ b444 ^ c444;
  assign sub444 = a444 ^ b_inv444 ^ c444;
  assign and444 = a444 & b444;
  assign or444  = a444 | b444;
  assign c445 = (a444 & b444) | (a444 & c444) | (b444 & c444);
  wire c_sub445;
  assign c_sub445 = (a444 & b_inv444) | (a444 & c444) | (b_inv444 & c444);
  wire s445, sub445, and445, or445;
  wire b_inv445;
  assign b_inv445 = ~b445;
  assign s445  = a445 ^ b445 ^ c445;
  assign sub445 = a445 ^ b_inv445 ^ c445;
  assign and445 = a445 & b445;
  assign or445  = a445 | b445;
  assign c446 = (a445 & b445) | (a445 & c445) | (b445 & c445);
  wire c_sub446;
  assign c_sub446 = (a445 & b_inv445) | (a445 & c445) | (b_inv445 & c445);
  wire s446, sub446, and446, or446;
  wire b_inv446;
  assign b_inv446 = ~b446;
  assign s446  = a446 ^ b446 ^ c446;
  assign sub446 = a446 ^ b_inv446 ^ c446;
  assign and446 = a446 & b446;
  assign or446  = a446 | b446;
  assign c447 = (a446 & b446) | (a446 & c446) | (b446 & c446);
  wire c_sub447;
  assign c_sub447 = (a446 & b_inv446) | (a446 & c446) | (b_inv446 & c446);
  wire s447, sub447, and447, or447;
  wire b_inv447;
  assign b_inv447 = ~b447;
  assign s447  = a447 ^ b447 ^ c447;
  assign sub447 = a447 ^ b_inv447 ^ c447;
  assign and447 = a447 & b447;
  assign or447  = a447 | b447;
  assign c448 = (a447 & b447) | (a447 & c447) | (b447 & c447);
  wire c_sub448;
  assign c_sub448 = (a447 & b_inv447) | (a447 & c447) | (b_inv447 & c447);
  wire s448, sub448, and448, or448;
  wire b_inv448;
  assign b_inv448 = ~b448;
  assign s448  = a448 ^ b448 ^ c448;
  assign sub448 = a448 ^ b_inv448 ^ c448;
  assign and448 = a448 & b448;
  assign or448  = a448 | b448;
  assign c449 = (a448 & b448) | (a448 & c448) | (b448 & c448);
  wire c_sub449;
  assign c_sub449 = (a448 & b_inv448) | (a448 & c448) | (b_inv448 & c448);
  wire s449, sub449, and449, or449;
  wire b_inv449;
  assign b_inv449 = ~b449;
  assign s449  = a449 ^ b449 ^ c449;
  assign sub449 = a449 ^ b_inv449 ^ c449;
  assign and449 = a449 & b449;
  assign or449  = a449 | b449;
  assign c450 = (a449 & b449) | (a449 & c449) | (b449 & c449);
  wire c_sub450;
  assign c_sub450 = (a449 & b_inv449) | (a449 & c449) | (b_inv449 & c449);
  wire s450, sub450, and450, or450;
  wire b_inv450;
  assign b_inv450 = ~b450;
  assign s450  = a450 ^ b450 ^ c450;
  assign sub450 = a450 ^ b_inv450 ^ c450;
  assign and450 = a450 & b450;
  assign or450  = a450 | b450;
  assign c451 = (a450 & b450) | (a450 & c450) | (b450 & c450);
  wire c_sub451;
  assign c_sub451 = (a450 & b_inv450) | (a450 & c450) | (b_inv450 & c450);
  wire s451, sub451, and451, or451;
  wire b_inv451;
  assign b_inv451 = ~b451;
  assign s451  = a451 ^ b451 ^ c451;
  assign sub451 = a451 ^ b_inv451 ^ c451;
  assign and451 = a451 & b451;
  assign or451  = a451 | b451;
  assign c452 = (a451 & b451) | (a451 & c451) | (b451 & c451);
  wire c_sub452;
  assign c_sub452 = (a451 & b_inv451) | (a451 & c451) | (b_inv451 & c451);
  wire s452, sub452, and452, or452;
  wire b_inv452;
  assign b_inv452 = ~b452;
  assign s452  = a452 ^ b452 ^ c452;
  assign sub452 = a452 ^ b_inv452 ^ c452;
  assign and452 = a452 & b452;
  assign or452  = a452 | b452;
  assign c453 = (a452 & b452) | (a452 & c452) | (b452 & c452);
  wire c_sub453;
  assign c_sub453 = (a452 & b_inv452) | (a452 & c452) | (b_inv452 & c452);
  wire s453, sub453, and453, or453;
  wire b_inv453;
  assign b_inv453 = ~b453;
  assign s453  = a453 ^ b453 ^ c453;
  assign sub453 = a453 ^ b_inv453 ^ c453;
  assign and453 = a453 & b453;
  assign or453  = a453 | b453;
  assign c454 = (a453 & b453) | (a453 & c453) | (b453 & c453);
  wire c_sub454;
  assign c_sub454 = (a453 & b_inv453) | (a453 & c453) | (b_inv453 & c453);
  wire s454, sub454, and454, or454;
  wire b_inv454;
  assign b_inv454 = ~b454;
  assign s454  = a454 ^ b454 ^ c454;
  assign sub454 = a454 ^ b_inv454 ^ c454;
  assign and454 = a454 & b454;
  assign or454  = a454 | b454;
  assign c455 = (a454 & b454) | (a454 & c454) | (b454 & c454);
  wire c_sub455;
  assign c_sub455 = (a454 & b_inv454) | (a454 & c454) | (b_inv454 & c454);
  wire s455, sub455, and455, or455;
  wire b_inv455;
  assign b_inv455 = ~b455;
  assign s455  = a455 ^ b455 ^ c455;
  assign sub455 = a455 ^ b_inv455 ^ c455;
  assign and455 = a455 & b455;
  assign or455  = a455 | b455;
  assign c456 = (a455 & b455) | (a455 & c455) | (b455 & c455);
  wire c_sub456;
  assign c_sub456 = (a455 & b_inv455) | (a455 & c455) | (b_inv455 & c455);
  wire s456, sub456, and456, or456;
  wire b_inv456;
  assign b_inv456 = ~b456;
  assign s456  = a456 ^ b456 ^ c456;
  assign sub456 = a456 ^ b_inv456 ^ c456;
  assign and456 = a456 & b456;
  assign or456  = a456 | b456;
  assign c457 = (a456 & b456) | (a456 & c456) | (b456 & c456);
  wire c_sub457;
  assign c_sub457 = (a456 & b_inv456) | (a456 & c456) | (b_inv456 & c456);
  wire s457, sub457, and457, or457;
  wire b_inv457;
  assign b_inv457 = ~b457;
  assign s457  = a457 ^ b457 ^ c457;
  assign sub457 = a457 ^ b_inv457 ^ c457;
  assign and457 = a457 & b457;
  assign or457  = a457 | b457;
  assign c458 = (a457 & b457) | (a457 & c457) | (b457 & c457);
  wire c_sub458;
  assign c_sub458 = (a457 & b_inv457) | (a457 & c457) | (b_inv457 & c457);
  wire s458, sub458, and458, or458;
  wire b_inv458;
  assign b_inv458 = ~b458;
  assign s458  = a458 ^ b458 ^ c458;
  assign sub458 = a458 ^ b_inv458 ^ c458;
  assign and458 = a458 & b458;
  assign or458  = a458 | b458;
  assign c459 = (a458 & b458) | (a458 & c458) | (b458 & c458);
  wire c_sub459;
  assign c_sub459 = (a458 & b_inv458) | (a458 & c458) | (b_inv458 & c458);
  wire s459, sub459, and459, or459;
  wire b_inv459;
  assign b_inv459 = ~b459;
  assign s459  = a459 ^ b459 ^ c459;
  assign sub459 = a459 ^ b_inv459 ^ c459;
  assign and459 = a459 & b459;
  assign or459  = a459 | b459;
  assign c460 = (a459 & b459) | (a459 & c459) | (b459 & c459);
  wire c_sub460;
  assign c_sub460 = (a459 & b_inv459) | (a459 & c459) | (b_inv459 & c459);
  wire s460, sub460, and460, or460;
  wire b_inv460;
  assign b_inv460 = ~b460;
  assign s460  = a460 ^ b460 ^ c460;
  assign sub460 = a460 ^ b_inv460 ^ c460;
  assign and460 = a460 & b460;
  assign or460  = a460 | b460;
  assign c461 = (a460 & b460) | (a460 & c460) | (b460 & c460);
  wire c_sub461;
  assign c_sub461 = (a460 & b_inv460) | (a460 & c460) | (b_inv460 & c460);
  wire s461, sub461, and461, or461;
  wire b_inv461;
  assign b_inv461 = ~b461;
  assign s461  = a461 ^ b461 ^ c461;
  assign sub461 = a461 ^ b_inv461 ^ c461;
  assign and461 = a461 & b461;
  assign or461  = a461 | b461;
  assign c462 = (a461 & b461) | (a461 & c461) | (b461 & c461);
  wire c_sub462;
  assign c_sub462 = (a461 & b_inv461) | (a461 & c461) | (b_inv461 & c461);
  wire s462, sub462, and462, or462;
  wire b_inv462;
  assign b_inv462 = ~b462;
  assign s462  = a462 ^ b462 ^ c462;
  assign sub462 = a462 ^ b_inv462 ^ c462;
  assign and462 = a462 & b462;
  assign or462  = a462 | b462;
  assign c463 = (a462 & b462) | (a462 & c462) | (b462 & c462);
  wire c_sub463;
  assign c_sub463 = (a462 & b_inv462) | (a462 & c462) | (b_inv462 & c462);
  wire s463, sub463, and463, or463;
  wire b_inv463;
  assign b_inv463 = ~b463;
  assign s463  = a463 ^ b463 ^ c463;
  assign sub463 = a463 ^ b_inv463 ^ c463;
  assign and463 = a463 & b463;
  assign or463  = a463 | b463;
  assign c464 = (a463 & b463) | (a463 & c463) | (b463 & c463);
  wire c_sub464;
  assign c_sub464 = (a463 & b_inv463) | (a463 & c463) | (b_inv463 & c463);
  wire s464, sub464, and464, or464;
  wire b_inv464;
  assign b_inv464 = ~b464;
  assign s464  = a464 ^ b464 ^ c464;
  assign sub464 = a464 ^ b_inv464 ^ c464;
  assign and464 = a464 & b464;
  assign or464  = a464 | b464;
  assign c465 = (a464 & b464) | (a464 & c464) | (b464 & c464);
  wire c_sub465;
  assign c_sub465 = (a464 & b_inv464) | (a464 & c464) | (b_inv464 & c464);
  wire s465, sub465, and465, or465;
  wire b_inv465;
  assign b_inv465 = ~b465;
  assign s465  = a465 ^ b465 ^ c465;
  assign sub465 = a465 ^ b_inv465 ^ c465;
  assign and465 = a465 & b465;
  assign or465  = a465 | b465;
  assign c466 = (a465 & b465) | (a465 & c465) | (b465 & c465);
  wire c_sub466;
  assign c_sub466 = (a465 & b_inv465) | (a465 & c465) | (b_inv465 & c465);
  wire s466, sub466, and466, or466;
  wire b_inv466;
  assign b_inv466 = ~b466;
  assign s466  = a466 ^ b466 ^ c466;
  assign sub466 = a466 ^ b_inv466 ^ c466;
  assign and466 = a466 & b466;
  assign or466  = a466 | b466;
  assign c467 = (a466 & b466) | (a466 & c466) | (b466 & c466);
  wire c_sub467;
  assign c_sub467 = (a466 & b_inv466) | (a466 & c466) | (b_inv466 & c466);
  wire s467, sub467, and467, or467;
  wire b_inv467;
  assign b_inv467 = ~b467;
  assign s467  = a467 ^ b467 ^ c467;
  assign sub467 = a467 ^ b_inv467 ^ c467;
  assign and467 = a467 & b467;
  assign or467  = a467 | b467;
  assign c468 = (a467 & b467) | (a467 & c467) | (b467 & c467);
  wire c_sub468;
  assign c_sub468 = (a467 & b_inv467) | (a467 & c467) | (b_inv467 & c467);
  wire s468, sub468, and468, or468;
  wire b_inv468;
  assign b_inv468 = ~b468;
  assign s468  = a468 ^ b468 ^ c468;
  assign sub468 = a468 ^ b_inv468 ^ c468;
  assign and468 = a468 & b468;
  assign or468  = a468 | b468;
  assign c469 = (a468 & b468) | (a468 & c468) | (b468 & c468);
  wire c_sub469;
  assign c_sub469 = (a468 & b_inv468) | (a468 & c468) | (b_inv468 & c468);
  wire s469, sub469, and469, or469;
  wire b_inv469;
  assign b_inv469 = ~b469;
  assign s469  = a469 ^ b469 ^ c469;
  assign sub469 = a469 ^ b_inv469 ^ c469;
  assign and469 = a469 & b469;
  assign or469  = a469 | b469;
  assign c470 = (a469 & b469) | (a469 & c469) | (b469 & c469);
  wire c_sub470;
  assign c_sub470 = (a469 & b_inv469) | (a469 & c469) | (b_inv469 & c469);
  wire s470, sub470, and470, or470;
  wire b_inv470;
  assign b_inv470 = ~b470;
  assign s470  = a470 ^ b470 ^ c470;
  assign sub470 = a470 ^ b_inv470 ^ c470;
  assign and470 = a470 & b470;
  assign or470  = a470 | b470;
  assign c471 = (a470 & b470) | (a470 & c470) | (b470 & c470);
  wire c_sub471;
  assign c_sub471 = (a470 & b_inv470) | (a470 & c470) | (b_inv470 & c470);
  wire s471, sub471, and471, or471;
  wire b_inv471;
  assign b_inv471 = ~b471;
  assign s471  = a471 ^ b471 ^ c471;
  assign sub471 = a471 ^ b_inv471 ^ c471;
  assign and471 = a471 & b471;
  assign or471  = a471 | b471;
  assign c472 = (a471 & b471) | (a471 & c471) | (b471 & c471);
  wire c_sub472;
  assign c_sub472 = (a471 & b_inv471) | (a471 & c471) | (b_inv471 & c471);
  wire s472, sub472, and472, or472;
  wire b_inv472;
  assign b_inv472 = ~b472;
  assign s472  = a472 ^ b472 ^ c472;
  assign sub472 = a472 ^ b_inv472 ^ c472;
  assign and472 = a472 & b472;
  assign or472  = a472 | b472;
  assign c473 = (a472 & b472) | (a472 & c472) | (b472 & c472);
  wire c_sub473;
  assign c_sub473 = (a472 & b_inv472) | (a472 & c472) | (b_inv472 & c472);
  wire s473, sub473, and473, or473;
  wire b_inv473;
  assign b_inv473 = ~b473;
  assign s473  = a473 ^ b473 ^ c473;
  assign sub473 = a473 ^ b_inv473 ^ c473;
  assign and473 = a473 & b473;
  assign or473  = a473 | b473;
  assign c474 = (a473 & b473) | (a473 & c473) | (b473 & c473);
  wire c_sub474;
  assign c_sub474 = (a473 & b_inv473) | (a473 & c473) | (b_inv473 & c473);
  wire s474, sub474, and474, or474;
  wire b_inv474;
  assign b_inv474 = ~b474;
  assign s474  = a474 ^ b474 ^ c474;
  assign sub474 = a474 ^ b_inv474 ^ c474;
  assign and474 = a474 & b474;
  assign or474  = a474 | b474;
  assign c475 = (a474 & b474) | (a474 & c474) | (b474 & c474);
  wire c_sub475;
  assign c_sub475 = (a474 & b_inv474) | (a474 & c474) | (b_inv474 & c474);
  wire s475, sub475, and475, or475;
  wire b_inv475;
  assign b_inv475 = ~b475;
  assign s475  = a475 ^ b475 ^ c475;
  assign sub475 = a475 ^ b_inv475 ^ c475;
  assign and475 = a475 & b475;
  assign or475  = a475 | b475;
  assign c476 = (a475 & b475) | (a475 & c475) | (b475 & c475);
  wire c_sub476;
  assign c_sub476 = (a475 & b_inv475) | (a475 & c475) | (b_inv475 & c475);
  wire s476, sub476, and476, or476;
  wire b_inv476;
  assign b_inv476 = ~b476;
  assign s476  = a476 ^ b476 ^ c476;
  assign sub476 = a476 ^ b_inv476 ^ c476;
  assign and476 = a476 & b476;
  assign or476  = a476 | b476;
  assign c477 = (a476 & b476) | (a476 & c476) | (b476 & c476);
  wire c_sub477;
  assign c_sub477 = (a476 & b_inv476) | (a476 & c476) | (b_inv476 & c476);
  wire s477, sub477, and477, or477;
  wire b_inv477;
  assign b_inv477 = ~b477;
  assign s477  = a477 ^ b477 ^ c477;
  assign sub477 = a477 ^ b_inv477 ^ c477;
  assign and477 = a477 & b477;
  assign or477  = a477 | b477;
  assign c478 = (a477 & b477) | (a477 & c477) | (b477 & c477);
  wire c_sub478;
  assign c_sub478 = (a477 & b_inv477) | (a477 & c477) | (b_inv477 & c477);
  wire s478, sub478, and478, or478;
  wire b_inv478;
  assign b_inv478 = ~b478;
  assign s478  = a478 ^ b478 ^ c478;
  assign sub478 = a478 ^ b_inv478 ^ c478;
  assign and478 = a478 & b478;
  assign or478  = a478 | b478;
  assign c479 = (a478 & b478) | (a478 & c478) | (b478 & c478);
  wire c_sub479;
  assign c_sub479 = (a478 & b_inv478) | (a478 & c478) | (b_inv478 & c478);
  wire s479, sub479, and479, or479;
  wire b_inv479;
  assign b_inv479 = ~b479;
  assign s479  = a479 ^ b479 ^ c479;
  assign sub479 = a479 ^ b_inv479 ^ c479;
  assign and479 = a479 & b479;
  assign or479  = a479 | b479;
  assign c480 = (a479 & b479) | (a479 & c479) | (b479 & c479);
  wire c_sub480;
  assign c_sub480 = (a479 & b_inv479) | (a479 & c479) | (b_inv479 & c479);
  wire s480, sub480, and480, or480;
  wire b_inv480;
  assign b_inv480 = ~b480;
  assign s480  = a480 ^ b480 ^ c480;
  assign sub480 = a480 ^ b_inv480 ^ c480;
  assign and480 = a480 & b480;
  assign or480  = a480 | b480;
  assign c481 = (a480 & b480) | (a480 & c480) | (b480 & c480);
  wire c_sub481;
  assign c_sub481 = (a480 & b_inv480) | (a480 & c480) | (b_inv480 & c480);
  wire s481, sub481, and481, or481;
  wire b_inv481;
  assign b_inv481 = ~b481;
  assign s481  = a481 ^ b481 ^ c481;
  assign sub481 = a481 ^ b_inv481 ^ c481;
  assign and481 = a481 & b481;
  assign or481  = a481 | b481;
  assign c482 = (a481 & b481) | (a481 & c481) | (b481 & c481);
  wire c_sub482;
  assign c_sub482 = (a481 & b_inv481) | (a481 & c481) | (b_inv481 & c481);
  wire s482, sub482, and482, or482;
  wire b_inv482;
  assign b_inv482 = ~b482;
  assign s482  = a482 ^ b482 ^ c482;
  assign sub482 = a482 ^ b_inv482 ^ c482;
  assign and482 = a482 & b482;
  assign or482  = a482 | b482;
  assign c483 = (a482 & b482) | (a482 & c482) | (b482 & c482);
  wire c_sub483;
  assign c_sub483 = (a482 & b_inv482) | (a482 & c482) | (b_inv482 & c482);
  wire s483, sub483, and483, or483;
  wire b_inv483;
  assign b_inv483 = ~b483;
  assign s483  = a483 ^ b483 ^ c483;
  assign sub483 = a483 ^ b_inv483 ^ c483;
  assign and483 = a483 & b483;
  assign or483  = a483 | b483;
  assign c484 = (a483 & b483) | (a483 & c483) | (b483 & c483);
  wire c_sub484;
  assign c_sub484 = (a483 & b_inv483) | (a483 & c483) | (b_inv483 & c483);
  wire s484, sub484, and484, or484;
  wire b_inv484;
  assign b_inv484 = ~b484;
  assign s484  = a484 ^ b484 ^ c484;
  assign sub484 = a484 ^ b_inv484 ^ c484;
  assign and484 = a484 & b484;
  assign or484  = a484 | b484;
  assign c485 = (a484 & b484) | (a484 & c484) | (b484 & c484);
  wire c_sub485;
  assign c_sub485 = (a484 & b_inv484) | (a484 & c484) | (b_inv484 & c484);
  wire s485, sub485, and485, or485;
  wire b_inv485;
  assign b_inv485 = ~b485;
  assign s485  = a485 ^ b485 ^ c485;
  assign sub485 = a485 ^ b_inv485 ^ c485;
  assign and485 = a485 & b485;
  assign or485  = a485 | b485;
  assign c486 = (a485 & b485) | (a485 & c485) | (b485 & c485);
  wire c_sub486;
  assign c_sub486 = (a485 & b_inv485) | (a485 & c485) | (b_inv485 & c485);
  wire s486, sub486, and486, or486;
  wire b_inv486;
  assign b_inv486 = ~b486;
  assign s486  = a486 ^ b486 ^ c486;
  assign sub486 = a486 ^ b_inv486 ^ c486;
  assign and486 = a486 & b486;
  assign or486  = a486 | b486;
  assign c487 = (a486 & b486) | (a486 & c486) | (b486 & c486);
  wire c_sub487;
  assign c_sub487 = (a486 & b_inv486) | (a486 & c486) | (b_inv486 & c486);
  wire s487, sub487, and487, or487;
  wire b_inv487;
  assign b_inv487 = ~b487;
  assign s487  = a487 ^ b487 ^ c487;
  assign sub487 = a487 ^ b_inv487 ^ c487;
  assign and487 = a487 & b487;
  assign or487  = a487 | b487;
  assign c488 = (a487 & b487) | (a487 & c487) | (b487 & c487);
  wire c_sub488;
  assign c_sub488 = (a487 & b_inv487) | (a487 & c487) | (b_inv487 & c487);
  wire s488, sub488, and488, or488;
  wire b_inv488;
  assign b_inv488 = ~b488;
  assign s488  = a488 ^ b488 ^ c488;
  assign sub488 = a488 ^ b_inv488 ^ c488;
  assign and488 = a488 & b488;
  assign or488  = a488 | b488;
  assign c489 = (a488 & b488) | (a488 & c488) | (b488 & c488);
  wire c_sub489;
  assign c_sub489 = (a488 & b_inv488) | (a488 & c488) | (b_inv488 & c488);
  wire s489, sub489, and489, or489;
  wire b_inv489;
  assign b_inv489 = ~b489;
  assign s489  = a489 ^ b489 ^ c489;
  assign sub489 = a489 ^ b_inv489 ^ c489;
  assign and489 = a489 & b489;
  assign or489  = a489 | b489;
  assign c490 = (a489 & b489) | (a489 & c489) | (b489 & c489);
  wire c_sub490;
  assign c_sub490 = (a489 & b_inv489) | (a489 & c489) | (b_inv489 & c489);
  wire s490, sub490, and490, or490;
  wire b_inv490;
  assign b_inv490 = ~b490;
  assign s490  = a490 ^ b490 ^ c490;
  assign sub490 = a490 ^ b_inv490 ^ c490;
  assign and490 = a490 & b490;
  assign or490  = a490 | b490;
  assign c491 = (a490 & b490) | (a490 & c490) | (b490 & c490);
  wire c_sub491;
  assign c_sub491 = (a490 & b_inv490) | (a490 & c490) | (b_inv490 & c490);
  wire s491, sub491, and491, or491;
  wire b_inv491;
  assign b_inv491 = ~b491;
  assign s491  = a491 ^ b491 ^ c491;
  assign sub491 = a491 ^ b_inv491 ^ c491;
  assign and491 = a491 & b491;
  assign or491  = a491 | b491;
  assign c492 = (a491 & b491) | (a491 & c491) | (b491 & c491);
  wire c_sub492;
  assign c_sub492 = (a491 & b_inv491) | (a491 & c491) | (b_inv491 & c491);
  wire s492, sub492, and492, or492;
  wire b_inv492;
  assign b_inv492 = ~b492;
  assign s492  = a492 ^ b492 ^ c492;
  assign sub492 = a492 ^ b_inv492 ^ c492;
  assign and492 = a492 & b492;
  assign or492  = a492 | b492;
  assign c493 = (a492 & b492) | (a492 & c492) | (b492 & c492);
  wire c_sub493;
  assign c_sub493 = (a492 & b_inv492) | (a492 & c492) | (b_inv492 & c492);
  wire s493, sub493, and493, or493;
  wire b_inv493;
  assign b_inv493 = ~b493;
  assign s493  = a493 ^ b493 ^ c493;
  assign sub493 = a493 ^ b_inv493 ^ c493;
  assign and493 = a493 & b493;
  assign or493  = a493 | b493;
  assign c494 = (a493 & b493) | (a493 & c493) | (b493 & c493);
  wire c_sub494;
  assign c_sub494 = (a493 & b_inv493) | (a493 & c493) | (b_inv493 & c493);
  wire s494, sub494, and494, or494;
  wire b_inv494;
  assign b_inv494 = ~b494;
  assign s494  = a494 ^ b494 ^ c494;
  assign sub494 = a494 ^ b_inv494 ^ c494;
  assign and494 = a494 & b494;
  assign or494  = a494 | b494;
  assign c495 = (a494 & b494) | (a494 & c494) | (b494 & c494);
  wire c_sub495;
  assign c_sub495 = (a494 & b_inv494) | (a494 & c494) | (b_inv494 & c494);
  wire s495, sub495, and495, or495;
  wire b_inv495;
  assign b_inv495 = ~b495;
  assign s495  = a495 ^ b495 ^ c495;
  assign sub495 = a495 ^ b_inv495 ^ c495;
  assign and495 = a495 & b495;
  assign or495  = a495 | b495;
  assign c496 = (a495 & b495) | (a495 & c495) | (b495 & c495);
  wire c_sub496;
  assign c_sub496 = (a495 & b_inv495) | (a495 & c495) | (b_inv495 & c495);
  wire s496, sub496, and496, or496;
  wire b_inv496;
  assign b_inv496 = ~b496;
  assign s496  = a496 ^ b496 ^ c496;
  assign sub496 = a496 ^ b_inv496 ^ c496;
  assign and496 = a496 & b496;
  assign or496  = a496 | b496;
  assign c497 = (a496 & b496) | (a496 & c496) | (b496 & c496);
  wire c_sub497;
  assign c_sub497 = (a496 & b_inv496) | (a496 & c496) | (b_inv496 & c496);
  wire s497, sub497, and497, or497;
  wire b_inv497;
  assign b_inv497 = ~b497;
  assign s497  = a497 ^ b497 ^ c497;
  assign sub497 = a497 ^ b_inv497 ^ c497;
  assign and497 = a497 & b497;
  assign or497  = a497 | b497;
  assign c498 = (a497 & b497) | (a497 & c497) | (b497 & c497);
  wire c_sub498;
  assign c_sub498 = (a497 & b_inv497) | (a497 & c497) | (b_inv497 & c497);
  wire s498, sub498, and498, or498;
  wire b_inv498;
  assign b_inv498 = ~b498;
  assign s498  = a498 ^ b498 ^ c498;
  assign sub498 = a498 ^ b_inv498 ^ c498;
  assign and498 = a498 & b498;
  assign or498  = a498 | b498;
  assign c499 = (a498 & b498) | (a498 & c498) | (b498 & c498);
  wire c_sub499;
  assign c_sub499 = (a498 & b_inv498) | (a498 & c498) | (b_inv498 & c498);
  wire s499, sub499, and499, or499;
  wire b_inv499;
  assign b_inv499 = ~b499;
  assign s499  = a499 ^ b499 ^ c499;
  assign sub499 = a499 ^ b_inv499 ^ c499;
  assign and499 = a499 & b499;
  assign or499  = a499 | b499;
  assign c500 = (a499 & b499) | (a499 & c499) | (b499 & c499);
  wire c_sub500;
  assign c_sub500 = (a499 & b_inv499) | (a499 & c499) | (b_inv499 & c499);
  wire s500, sub500, and500, or500;
  wire b_inv500;
  assign b_inv500 = ~b500;
  assign s500  = a500 ^ b500 ^ c500;
  assign sub500 = a500 ^ b_inv500 ^ c500;
  assign and500 = a500 & b500;
  assign or500  = a500 | b500;
  assign c501 = (a500 & b500) | (a500 & c500) | (b500 & c500);
  wire c_sub501;
  assign c_sub501 = (a500 & b_inv500) | (a500 & c500) | (b_inv500 & c500);
  wire s501, sub501, and501, or501;
  wire b_inv501;
  assign b_inv501 = ~b501;
  assign s501  = a501 ^ b501 ^ c501;
  assign sub501 = a501 ^ b_inv501 ^ c501;
  assign and501 = a501 & b501;
  assign or501  = a501 | b501;
  assign c502 = (a501 & b501) | (a501 & c501) | (b501 & c501);
  wire c_sub502;
  assign c_sub502 = (a501 & b_inv501) | (a501 & c501) | (b_inv501 & c501);
  wire s502, sub502, and502, or502;
  wire b_inv502;
  assign b_inv502 = ~b502;
  assign s502  = a502 ^ b502 ^ c502;
  assign sub502 = a502 ^ b_inv502 ^ c502;
  assign and502 = a502 & b502;
  assign or502  = a502 | b502;
  assign c503 = (a502 & b502) | (a502 & c502) | (b502 & c502);
  wire c_sub503;
  assign c_sub503 = (a502 & b_inv502) | (a502 & c502) | (b_inv502 & c502);
  wire s503, sub503, and503, or503;
  wire b_inv503;
  assign b_inv503 = ~b503;
  assign s503  = a503 ^ b503 ^ c503;
  assign sub503 = a503 ^ b_inv503 ^ c503;
  assign and503 = a503 & b503;
  assign or503  = a503 | b503;
  assign c504 = (a503 & b503) | (a503 & c503) | (b503 & c503);
  wire c_sub504;
  assign c_sub504 = (a503 & b_inv503) | (a503 & c503) | (b_inv503 & c503);
  wire s504, sub504, and504, or504;
  wire b_inv504;
  assign b_inv504 = ~b504;
  assign s504  = a504 ^ b504 ^ c504;
  assign sub504 = a504 ^ b_inv504 ^ c504;
  assign and504 = a504 & b504;
  assign or504  = a504 | b504;
  assign c505 = (a504 & b504) | (a504 & c504) | (b504 & c504);
  wire c_sub505;
  assign c_sub505 = (a504 & b_inv504) | (a504 & c504) | (b_inv504 & c504);
  wire s505, sub505, and505, or505;
  wire b_inv505;
  assign b_inv505 = ~b505;
  assign s505  = a505 ^ b505 ^ c505;
  assign sub505 = a505 ^ b_inv505 ^ c505;
  assign and505 = a505 & b505;
  assign or505  = a505 | b505;
  assign c506 = (a505 & b505) | (a505 & c505) | (b505 & c505);
  wire c_sub506;
  assign c_sub506 = (a505 & b_inv505) | (a505 & c505) | (b_inv505 & c505);
  wire s506, sub506, and506, or506;
  wire b_inv506;
  assign b_inv506 = ~b506;
  assign s506  = a506 ^ b506 ^ c506;
  assign sub506 = a506 ^ b_inv506 ^ c506;
  assign and506 = a506 & b506;
  assign or506  = a506 | b506;
  assign c507 = (a506 & b506) | (a506 & c506) | (b506 & c506);
  wire c_sub507;
  assign c_sub507 = (a506 & b_inv506) | (a506 & c506) | (b_inv506 & c506);
  wire s507, sub507, and507, or507;
  wire b_inv507;
  assign b_inv507 = ~b507;
  assign s507  = a507 ^ b507 ^ c507;
  assign sub507 = a507 ^ b_inv507 ^ c507;
  assign and507 = a507 & b507;
  assign or507  = a507 | b507;
  assign c508 = (a507 & b507) | (a507 & c507) | (b507 & c507);
  wire c_sub508;
  assign c_sub508 = (a507 & b_inv507) | (a507 & c507) | (b_inv507 & c507);
  wire s508, sub508, and508, or508;
  wire b_inv508;
  assign b_inv508 = ~b508;
  assign s508  = a508 ^ b508 ^ c508;
  assign sub508 = a508 ^ b_inv508 ^ c508;
  assign and508 = a508 & b508;
  assign or508  = a508 | b508;
  assign c509 = (a508 & b508) | (a508 & c508) | (b508 & c508);
  wire c_sub509;
  assign c_sub509 = (a508 & b_inv508) | (a508 & c508) | (b_inv508 & c508);
  wire s509, sub509, and509, or509;
  wire b_inv509;
  assign b_inv509 = ~b509;
  assign s509  = a509 ^ b509 ^ c509;
  assign sub509 = a509 ^ b_inv509 ^ c509;
  assign and509 = a509 & b509;
  assign or509  = a509 | b509;
  assign c510 = (a509 & b509) | (a509 & c509) | (b509 & c509);
  wire c_sub510;
  assign c_sub510 = (a509 & b_inv509) | (a509 & c509) | (b_inv509 & c509);
  wire s510, sub510, and510, or510;
  wire b_inv510;
  assign b_inv510 = ~b510;
  assign s510  = a510 ^ b510 ^ c510;
  assign sub510 = a510 ^ b_inv510 ^ c510;
  assign and510 = a510 & b510;
  assign or510  = a510 | b510;
  assign c511 = (a510 & b510) | (a510 & c510) | (b510 & c510);
  wire c_sub511;
  assign c_sub511 = (a510 & b_inv510) | (a510 & c510) | (b_inv510 & c510);
  wire s511, sub511, and511, or511;
  wire b_inv511;
  assign b_inv511 = ~b511;
  assign s511  = a511 ^ b511 ^ c511;
  assign sub511 = a511 ^ b_inv511 ^ c511;
  assign and511 = a511 & b511;
  assign or511  = a511 | b511;
  assign c512 = (a511 & b511) | (a511 & c511) | (b511 & c511);
  wire c_sub512;
  assign c_sub512 = (a511 & b_inv511) | (a511 & c511) | (b_inv511 & c511);
  wire s512, sub512, and512, or512;
  wire b_inv512;
  assign b_inv512 = ~b512;
  assign s512  = a512 ^ b512 ^ c512;
  assign sub512 = a512 ^ b_inv512 ^ c512;
  assign and512 = a512 & b512;
  assign or512  = a512 | b512;
  assign c513 = (a512 & b512) | (a512 & c512) | (b512 & c512);
  wire c_sub513;
  assign c_sub513 = (a512 & b_inv512) | (a512 & c512) | (b_inv512 & c512);
  wire s513, sub513, and513, or513;
  wire b_inv513;
  assign b_inv513 = ~b513;
  assign s513  = a513 ^ b513 ^ c513;
  assign sub513 = a513 ^ b_inv513 ^ c513;
  assign and513 = a513 & b513;
  assign or513  = a513 | b513;
  assign c514 = (a513 & b513) | (a513 & c513) | (b513 & c513);
  wire c_sub514;
  assign c_sub514 = (a513 & b_inv513) | (a513 & c513) | (b_inv513 & c513);
  wire s514, sub514, and514, or514;
  wire b_inv514;
  assign b_inv514 = ~b514;
  assign s514  = a514 ^ b514 ^ c514;
  assign sub514 = a514 ^ b_inv514 ^ c514;
  assign and514 = a514 & b514;
  assign or514  = a514 | b514;
  assign c515 = (a514 & b514) | (a514 & c514) | (b514 & c514);
  wire c_sub515;
  assign c_sub515 = (a514 & b_inv514) | (a514 & c514) | (b_inv514 & c514);
  wire s515, sub515, and515, or515;
  wire b_inv515;
  assign b_inv515 = ~b515;
  assign s515  = a515 ^ b515 ^ c515;
  assign sub515 = a515 ^ b_inv515 ^ c515;
  assign and515 = a515 & b515;
  assign or515  = a515 | b515;
  assign c516 = (a515 & b515) | (a515 & c515) | (b515 & c515);
  wire c_sub516;
  assign c_sub516 = (a515 & b_inv515) | (a515 & c515) | (b_inv515 & c515);
  wire s516, sub516, and516, or516;
  wire b_inv516;
  assign b_inv516 = ~b516;
  assign s516  = a516 ^ b516 ^ c516;
  assign sub516 = a516 ^ b_inv516 ^ c516;
  assign and516 = a516 & b516;
  assign or516  = a516 | b516;
  assign c517 = (a516 & b516) | (a516 & c516) | (b516 & c516);
  wire c_sub517;
  assign c_sub517 = (a516 & b_inv516) | (a516 & c516) | (b_inv516 & c516);
  wire s517, sub517, and517, or517;
  wire b_inv517;
  assign b_inv517 = ~b517;
  assign s517  = a517 ^ b517 ^ c517;
  assign sub517 = a517 ^ b_inv517 ^ c517;
  assign and517 = a517 & b517;
  assign or517  = a517 | b517;
  assign c518 = (a517 & b517) | (a517 & c517) | (b517 & c517);
  wire c_sub518;
  assign c_sub518 = (a517 & b_inv517) | (a517 & c517) | (b_inv517 & c517);
  wire s518, sub518, and518, or518;
  wire b_inv518;
  assign b_inv518 = ~b518;
  assign s518  = a518 ^ b518 ^ c518;
  assign sub518 = a518 ^ b_inv518 ^ c518;
  assign and518 = a518 & b518;
  assign or518  = a518 | b518;
  assign c519 = (a518 & b518) | (a518 & c518) | (b518 & c518);
  wire c_sub519;
  assign c_sub519 = (a518 & b_inv518) | (a518 & c518) | (b_inv518 & c518);
  wire s519, sub519, and519, or519;
  wire b_inv519;
  assign b_inv519 = ~b519;
  assign s519  = a519 ^ b519 ^ c519;
  assign sub519 = a519 ^ b_inv519 ^ c519;
  assign and519 = a519 & b519;
  assign or519  = a519 | b519;
  assign c520 = (a519 & b519) | (a519 & c519) | (b519 & c519);
  wire c_sub520;
  assign c_sub520 = (a519 & b_inv519) | (a519 & c519) | (b_inv519 & c519);
  wire s520, sub520, and520, or520;
  wire b_inv520;
  assign b_inv520 = ~b520;
  assign s520  = a520 ^ b520 ^ c520;
  assign sub520 = a520 ^ b_inv520 ^ c520;
  assign and520 = a520 & b520;
  assign or520  = a520 | b520;
  assign c521 = (a520 & b520) | (a520 & c520) | (b520 & c520);
  wire c_sub521;
  assign c_sub521 = (a520 & b_inv520) | (a520 & c520) | (b_inv520 & c520);
  wire s521, sub521, and521, or521;
  wire b_inv521;
  assign b_inv521 = ~b521;
  assign s521  = a521 ^ b521 ^ c521;
  assign sub521 = a521 ^ b_inv521 ^ c521;
  assign and521 = a521 & b521;
  assign or521  = a521 | b521;
  assign c522 = (a521 & b521) | (a521 & c521) | (b521 & c521);
  wire c_sub522;
  assign c_sub522 = (a521 & b_inv521) | (a521 & c521) | (b_inv521 & c521);
  wire s522, sub522, and522, or522;
  wire b_inv522;
  assign b_inv522 = ~b522;
  assign s522  = a522 ^ b522 ^ c522;
  assign sub522 = a522 ^ b_inv522 ^ c522;
  assign and522 = a522 & b522;
  assign or522  = a522 | b522;
  assign c523 = (a522 & b522) | (a522 & c522) | (b522 & c522);
  wire c_sub523;
  assign c_sub523 = (a522 & b_inv522) | (a522 & c522) | (b_inv522 & c522);
  wire s523, sub523, and523, or523;
  wire b_inv523;
  assign b_inv523 = ~b523;
  assign s523  = a523 ^ b523 ^ c523;
  assign sub523 = a523 ^ b_inv523 ^ c523;
  assign and523 = a523 & b523;
  assign or523  = a523 | b523;
  assign c524 = (a523 & b523) | (a523 & c523) | (b523 & c523);
  wire c_sub524;
  assign c_sub524 = (a523 & b_inv523) | (a523 & c523) | (b_inv523 & c523);
  wire s524, sub524, and524, or524;
  wire b_inv524;
  assign b_inv524 = ~b524;
  assign s524  = a524 ^ b524 ^ c524;
  assign sub524 = a524 ^ b_inv524 ^ c524;
  assign and524 = a524 & b524;
  assign or524  = a524 | b524;
  assign c525 = (a524 & b524) | (a524 & c524) | (b524 & c524);
  wire c_sub525;
  assign c_sub525 = (a524 & b_inv524) | (a524 & c524) | (b_inv524 & c524);
  wire s525, sub525, and525, or525;
  wire b_inv525;
  assign b_inv525 = ~b525;
  assign s525  = a525 ^ b525 ^ c525;
  assign sub525 = a525 ^ b_inv525 ^ c525;
  assign and525 = a525 & b525;
  assign or525  = a525 | b525;
  assign c526 = (a525 & b525) | (a525 & c525) | (b525 & c525);
  wire c_sub526;
  assign c_sub526 = (a525 & b_inv525) | (a525 & c525) | (b_inv525 & c525);
  wire s526, sub526, and526, or526;
  wire b_inv526;
  assign b_inv526 = ~b526;
  assign s526  = a526 ^ b526 ^ c526;
  assign sub526 = a526 ^ b_inv526 ^ c526;
  assign and526 = a526 & b526;
  assign or526  = a526 | b526;
  assign c527 = (a526 & b526) | (a526 & c526) | (b526 & c526);
  wire c_sub527;
  assign c_sub527 = (a526 & b_inv526) | (a526 & c526) | (b_inv526 & c526);
  wire s527, sub527, and527, or527;
  wire b_inv527;
  assign b_inv527 = ~b527;
  assign s527  = a527 ^ b527 ^ c527;
  assign sub527 = a527 ^ b_inv527 ^ c527;
  assign and527 = a527 & b527;
  assign or527  = a527 | b527;
  assign c528 = (a527 & b527) | (a527 & c527) | (b527 & c527);
  wire c_sub528;
  assign c_sub528 = (a527 & b_inv527) | (a527 & c527) | (b_inv527 & c527);
  wire s528, sub528, and528, or528;
  wire b_inv528;
  assign b_inv528 = ~b528;
  assign s528  = a528 ^ b528 ^ c528;
  assign sub528 = a528 ^ b_inv528 ^ c528;
  assign and528 = a528 & b528;
  assign or528  = a528 | b528;
  assign c529 = (a528 & b528) | (a528 & c528) | (b528 & c528);
  wire c_sub529;
  assign c_sub529 = (a528 & b_inv528) | (a528 & c528) | (b_inv528 & c528);
  wire s529, sub529, and529, or529;
  wire b_inv529;
  assign b_inv529 = ~b529;
  assign s529  = a529 ^ b529 ^ c529;
  assign sub529 = a529 ^ b_inv529 ^ c529;
  assign and529 = a529 & b529;
  assign or529  = a529 | b529;
  assign c530 = (a529 & b529) | (a529 & c529) | (b529 & c529);
  wire c_sub530;
  assign c_sub530 = (a529 & b_inv529) | (a529 & c529) | (b_inv529 & c529);
  wire s530, sub530, and530, or530;
  wire b_inv530;
  assign b_inv530 = ~b530;
  assign s530  = a530 ^ b530 ^ c530;
  assign sub530 = a530 ^ b_inv530 ^ c530;
  assign and530 = a530 & b530;
  assign or530  = a530 | b530;
  assign c531 = (a530 & b530) | (a530 & c530) | (b530 & c530);
  wire c_sub531;
  assign c_sub531 = (a530 & b_inv530) | (a530 & c530) | (b_inv530 & c530);
  wire s531, sub531, and531, or531;
  wire b_inv531;
  assign b_inv531 = ~b531;
  assign s531  = a531 ^ b531 ^ c531;
  assign sub531 = a531 ^ b_inv531 ^ c531;
  assign and531 = a531 & b531;
  assign or531  = a531 | b531;
  assign c532 = (a531 & b531) | (a531 & c531) | (b531 & c531);
  wire c_sub532;
  assign c_sub532 = (a531 & b_inv531) | (a531 & c531) | (b_inv531 & c531);
  wire s532, sub532, and532, or532;
  wire b_inv532;
  assign b_inv532 = ~b532;
  assign s532  = a532 ^ b532 ^ c532;
  assign sub532 = a532 ^ b_inv532 ^ c532;
  assign and532 = a532 & b532;
  assign or532  = a532 | b532;
  assign c533 = (a532 & b532) | (a532 & c532) | (b532 & c532);
  wire c_sub533;
  assign c_sub533 = (a532 & b_inv532) | (a532 & c532) | (b_inv532 & c532);
  wire s533, sub533, and533, or533;
  wire b_inv533;
  assign b_inv533 = ~b533;
  assign s533  = a533 ^ b533 ^ c533;
  assign sub533 = a533 ^ b_inv533 ^ c533;
  assign and533 = a533 & b533;
  assign or533  = a533 | b533;
  assign c534 = (a533 & b533) | (a533 & c533) | (b533 & c533);
  wire c_sub534;
  assign c_sub534 = (a533 & b_inv533) | (a533 & c533) | (b_inv533 & c533);
  wire s534, sub534, and534, or534;
  wire b_inv534;
  assign b_inv534 = ~b534;
  assign s534  = a534 ^ b534 ^ c534;
  assign sub534 = a534 ^ b_inv534 ^ c534;
  assign and534 = a534 & b534;
  assign or534  = a534 | b534;
  assign c535 = (a534 & b534) | (a534 & c534) | (b534 & c534);
  wire c_sub535;
  assign c_sub535 = (a534 & b_inv534) | (a534 & c534) | (b_inv534 & c534);
  wire s535, sub535, and535, or535;
  wire b_inv535;
  assign b_inv535 = ~b535;
  assign s535  = a535 ^ b535 ^ c535;
  assign sub535 = a535 ^ b_inv535 ^ c535;
  assign and535 = a535 & b535;
  assign or535  = a535 | b535;
  assign c536 = (a535 & b535) | (a535 & c535) | (b535 & c535);
  wire c_sub536;
  assign c_sub536 = (a535 & b_inv535) | (a535 & c535) | (b_inv535 & c535);
  wire s536, sub536, and536, or536;
  wire b_inv536;
  assign b_inv536 = ~b536;
  assign s536  = a536 ^ b536 ^ c536;
  assign sub536 = a536 ^ b_inv536 ^ c536;
  assign and536 = a536 & b536;
  assign or536  = a536 | b536;
  assign c537 = (a536 & b536) | (a536 & c536) | (b536 & c536);
  wire c_sub537;
  assign c_sub537 = (a536 & b_inv536) | (a536 & c536) | (b_inv536 & c536);
  wire s537, sub537, and537, or537;
  wire b_inv537;
  assign b_inv537 = ~b537;
  assign s537  = a537 ^ b537 ^ c537;
  assign sub537 = a537 ^ b_inv537 ^ c537;
  assign and537 = a537 & b537;
  assign or537  = a537 | b537;
  assign c538 = (a537 & b537) | (a537 & c537) | (b537 & c537);
  wire c_sub538;
  assign c_sub538 = (a537 & b_inv537) | (a537 & c537) | (b_inv537 & c537);
  wire s538, sub538, and538, or538;
  wire b_inv538;
  assign b_inv538 = ~b538;
  assign s538  = a538 ^ b538 ^ c538;
  assign sub538 = a538 ^ b_inv538 ^ c538;
  assign and538 = a538 & b538;
  assign or538  = a538 | b538;
  assign c539 = (a538 & b538) | (a538 & c538) | (b538 & c538);
  wire c_sub539;
  assign c_sub539 = (a538 & b_inv538) | (a538 & c538) | (b_inv538 & c538);
  wire s539, sub539, and539, or539;
  wire b_inv539;
  assign b_inv539 = ~b539;
  assign s539  = a539 ^ b539 ^ c539;
  assign sub539 = a539 ^ b_inv539 ^ c539;
  assign and539 = a539 & b539;
  assign or539  = a539 | b539;
  assign c540 = (a539 & b539) | (a539 & c539) | (b539 & c539);
  wire c_sub540;
  assign c_sub540 = (a539 & b_inv539) | (a539 & c539) | (b_inv539 & c539);
  wire s540, sub540, and540, or540;
  wire b_inv540;
  assign b_inv540 = ~b540;
  assign s540  = a540 ^ b540 ^ c540;
  assign sub540 = a540 ^ b_inv540 ^ c540;
  assign and540 = a540 & b540;
  assign or540  = a540 | b540;
  assign c541 = (a540 & b540) | (a540 & c540) | (b540 & c540);
  wire c_sub541;
  assign c_sub541 = (a540 & b_inv540) | (a540 & c540) | (b_inv540 & c540);
  wire s541, sub541, and541, or541;
  wire b_inv541;
  assign b_inv541 = ~b541;
  assign s541  = a541 ^ b541 ^ c541;
  assign sub541 = a541 ^ b_inv541 ^ c541;
  assign and541 = a541 & b541;
  assign or541  = a541 | b541;
  assign c542 = (a541 & b541) | (a541 & c541) | (b541 & c541);
  wire c_sub542;
  assign c_sub542 = (a541 & b_inv541) | (a541 & c541) | (b_inv541 & c541);
  wire s542, sub542, and542, or542;
  wire b_inv542;
  assign b_inv542 = ~b542;
  assign s542  = a542 ^ b542 ^ c542;
  assign sub542 = a542 ^ b_inv542 ^ c542;
  assign and542 = a542 & b542;
  assign or542  = a542 | b542;
  assign c543 = (a542 & b542) | (a542 & c542) | (b542 & c542);
  wire c_sub543;
  assign c_sub543 = (a542 & b_inv542) | (a542 & c542) | (b_inv542 & c542);
  wire s543, sub543, and543, or543;
  wire b_inv543;
  assign b_inv543 = ~b543;
  assign s543  = a543 ^ b543 ^ c543;
  assign sub543 = a543 ^ b_inv543 ^ c543;
  assign and543 = a543 & b543;
  assign or543  = a543 | b543;
  assign c544 = (a543 & b543) | (a543 & c543) | (b543 & c543);
  wire c_sub544;
  assign c_sub544 = (a543 & b_inv543) | (a543 & c543) | (b_inv543 & c543);
  wire s544, sub544, and544, or544;
  wire b_inv544;
  assign b_inv544 = ~b544;
  assign s544  = a544 ^ b544 ^ c544;
  assign sub544 = a544 ^ b_inv544 ^ c544;
  assign and544 = a544 & b544;
  assign or544  = a544 | b544;
  assign c545 = (a544 & b544) | (a544 & c544) | (b544 & c544);
  wire c_sub545;
  assign c_sub545 = (a544 & b_inv544) | (a544 & c544) | (b_inv544 & c544);
  wire s545, sub545, and545, or545;
  wire b_inv545;
  assign b_inv545 = ~b545;
  assign s545  = a545 ^ b545 ^ c545;
  assign sub545 = a545 ^ b_inv545 ^ c545;
  assign and545 = a545 & b545;
  assign or545  = a545 | b545;
  assign c546 = (a545 & b545) | (a545 & c545) | (b545 & c545);
  wire c_sub546;
  assign c_sub546 = (a545 & b_inv545) | (a545 & c545) | (b_inv545 & c545);
  wire s546, sub546, and546, or546;
  wire b_inv546;
  assign b_inv546 = ~b546;
  assign s546  = a546 ^ b546 ^ c546;
  assign sub546 = a546 ^ b_inv546 ^ c546;
  assign and546 = a546 & b546;
  assign or546  = a546 | b546;
  assign c547 = (a546 & b546) | (a546 & c546) | (b546 & c546);
  wire c_sub547;
  assign c_sub547 = (a546 & b_inv546) | (a546 & c546) | (b_inv546 & c546);
  wire s547, sub547, and547, or547;
  wire b_inv547;
  assign b_inv547 = ~b547;
  assign s547  = a547 ^ b547 ^ c547;
  assign sub547 = a547 ^ b_inv547 ^ c547;
  assign and547 = a547 & b547;
  assign or547  = a547 | b547;
  assign c548 = (a547 & b547) | (a547 & c547) | (b547 & c547);
  wire c_sub548;
  assign c_sub548 = (a547 & b_inv547) | (a547 & c547) | (b_inv547 & c547);
  wire s548, sub548, and548, or548;
  wire b_inv548;
  assign b_inv548 = ~b548;
  assign s548  = a548 ^ b548 ^ c548;
  assign sub548 = a548 ^ b_inv548 ^ c548;
  assign and548 = a548 & b548;
  assign or548  = a548 | b548;
  assign c549 = (a548 & b548) | (a548 & c548) | (b548 & c548);
  wire c_sub549;
  assign c_sub549 = (a548 & b_inv548) | (a548 & c548) | (b_inv548 & c548);
  wire s549, sub549, and549, or549;
  wire b_inv549;
  assign b_inv549 = ~b549;
  assign s549  = a549 ^ b549 ^ c549;
  assign sub549 = a549 ^ b_inv549 ^ c549;
  assign and549 = a549 & b549;
  assign or549  = a549 | b549;
  assign c550 = (a549 & b549) | (a549 & c549) | (b549 & c549);
  wire c_sub550;
  assign c_sub550 = (a549 & b_inv549) | (a549 & c549) | (b_inv549 & c549);
  wire s550, sub550, and550, or550;
  wire b_inv550;
  assign b_inv550 = ~b550;
  assign s550  = a550 ^ b550 ^ c550;
  assign sub550 = a550 ^ b_inv550 ^ c550;
  assign and550 = a550 & b550;
  assign or550  = a550 | b550;
  assign c551 = (a550 & b550) | (a550 & c550) | (b550 & c550);
  wire c_sub551;
  assign c_sub551 = (a550 & b_inv550) | (a550 & c550) | (b_inv550 & c550);
  wire s551, sub551, and551, or551;
  wire b_inv551;
  assign b_inv551 = ~b551;
  assign s551  = a551 ^ b551 ^ c551;
  assign sub551 = a551 ^ b_inv551 ^ c551;
  assign and551 = a551 & b551;
  assign or551  = a551 | b551;
  assign c552 = (a551 & b551) | (a551 & c551) | (b551 & c551);
  wire c_sub552;
  assign c_sub552 = (a551 & b_inv551) | (a551 & c551) | (b_inv551 & c551);
  wire s552, sub552, and552, or552;
  wire b_inv552;
  assign b_inv552 = ~b552;
  assign s552  = a552 ^ b552 ^ c552;
  assign sub552 = a552 ^ b_inv552 ^ c552;
  assign and552 = a552 & b552;
  assign or552  = a552 | b552;
  assign c553 = (a552 & b552) | (a552 & c552) | (b552 & c552);
  wire c_sub553;
  assign c_sub553 = (a552 & b_inv552) | (a552 & c552) | (b_inv552 & c552);
  wire s553, sub553, and553, or553;
  wire b_inv553;
  assign b_inv553 = ~b553;
  assign s553  = a553 ^ b553 ^ c553;
  assign sub553 = a553 ^ b_inv553 ^ c553;
  assign and553 = a553 & b553;
  assign or553  = a553 | b553;
  assign c554 = (a553 & b553) | (a553 & c553) | (b553 & c553);
  wire c_sub554;
  assign c_sub554 = (a553 & b_inv553) | (a553 & c553) | (b_inv553 & c553);
  wire s554, sub554, and554, or554;
  wire b_inv554;
  assign b_inv554 = ~b554;
  assign s554  = a554 ^ b554 ^ c554;
  assign sub554 = a554 ^ b_inv554 ^ c554;
  assign and554 = a554 & b554;
  assign or554  = a554 | b554;
  assign c555 = (a554 & b554) | (a554 & c554) | (b554 & c554);
  wire c_sub555;
  assign c_sub555 = (a554 & b_inv554) | (a554 & c554) | (b_inv554 & c554);
  wire s555, sub555, and555, or555;
  wire b_inv555;
  assign b_inv555 = ~b555;
  assign s555  = a555 ^ b555 ^ c555;
  assign sub555 = a555 ^ b_inv555 ^ c555;
  assign and555 = a555 & b555;
  assign or555  = a555 | b555;
  assign c556 = (a555 & b555) | (a555 & c555) | (b555 & c555);
  wire c_sub556;
  assign c_sub556 = (a555 & b_inv555) | (a555 & c555) | (b_inv555 & c555);
  wire s556, sub556, and556, or556;
  wire b_inv556;
  assign b_inv556 = ~b556;
  assign s556  = a556 ^ b556 ^ c556;
  assign sub556 = a556 ^ b_inv556 ^ c556;
  assign and556 = a556 & b556;
  assign or556  = a556 | b556;
  assign c557 = (a556 & b556) | (a556 & c556) | (b556 & c556);
  wire c_sub557;
  assign c_sub557 = (a556 & b_inv556) | (a556 & c556) | (b_inv556 & c556);
  wire s557, sub557, and557, or557;
  wire b_inv557;
  assign b_inv557 = ~b557;
  assign s557  = a557 ^ b557 ^ c557;
  assign sub557 = a557 ^ b_inv557 ^ c557;
  assign and557 = a557 & b557;
  assign or557  = a557 | b557;
  assign c558 = (a557 & b557) | (a557 & c557) | (b557 & c557);
  wire c_sub558;
  assign c_sub558 = (a557 & b_inv557) | (a557 & c557) | (b_inv557 & c557);
  wire s558, sub558, and558, or558;
  wire b_inv558;
  assign b_inv558 = ~b558;
  assign s558  = a558 ^ b558 ^ c558;
  assign sub558 = a558 ^ b_inv558 ^ c558;
  assign and558 = a558 & b558;
  assign or558  = a558 | b558;
  assign c559 = (a558 & b558) | (a558 & c558) | (b558 & c558);
  wire c_sub559;
  assign c_sub559 = (a558 & b_inv558) | (a558 & c558) | (b_inv558 & c558);
  wire s559, sub559, and559, or559;
  wire b_inv559;
  assign b_inv559 = ~b559;
  assign s559  = a559 ^ b559 ^ c559;
  assign sub559 = a559 ^ b_inv559 ^ c559;
  assign and559 = a559 & b559;
  assign or559  = a559 | b559;
  assign c560 = (a559 & b559) | (a559 & c559) | (b559 & c559);
  wire c_sub560;
  assign c_sub560 = (a559 & b_inv559) | (a559 & c559) | (b_inv559 & c559);
  wire s560, sub560, and560, or560;
  wire b_inv560;
  assign b_inv560 = ~b560;
  assign s560  = a560 ^ b560 ^ c560;
  assign sub560 = a560 ^ b_inv560 ^ c560;
  assign and560 = a560 & b560;
  assign or560  = a560 | b560;
  assign c561 = (a560 & b560) | (a560 & c560) | (b560 & c560);
  wire c_sub561;
  assign c_sub561 = (a560 & b_inv560) | (a560 & c560) | (b_inv560 & c560);
  wire s561, sub561, and561, or561;
  wire b_inv561;
  assign b_inv561 = ~b561;
  assign s561  = a561 ^ b561 ^ c561;
  assign sub561 = a561 ^ b_inv561 ^ c561;
  assign and561 = a561 & b561;
  assign or561  = a561 | b561;
  assign c562 = (a561 & b561) | (a561 & c561) | (b561 & c561);
  wire c_sub562;
  assign c_sub562 = (a561 & b_inv561) | (a561 & c561) | (b_inv561 & c561);
  wire s562, sub562, and562, or562;
  wire b_inv562;
  assign b_inv562 = ~b562;
  assign s562  = a562 ^ b562 ^ c562;
  assign sub562 = a562 ^ b_inv562 ^ c562;
  assign and562 = a562 & b562;
  assign or562  = a562 | b562;
  assign c563 = (a562 & b562) | (a562 & c562) | (b562 & c562);
  wire c_sub563;
  assign c_sub563 = (a562 & b_inv562) | (a562 & c562) | (b_inv562 & c562);
  wire s563, sub563, and563, or563;
  wire b_inv563;
  assign b_inv563 = ~b563;
  assign s563  = a563 ^ b563 ^ c563;
  assign sub563 = a563 ^ b_inv563 ^ c563;
  assign and563 = a563 & b563;
  assign or563  = a563 | b563;
  assign c564 = (a563 & b563) | (a563 & c563) | (b563 & c563);
  wire c_sub564;
  assign c_sub564 = (a563 & b_inv563) | (a563 & c563) | (b_inv563 & c563);
  wire s564, sub564, and564, or564;
  wire b_inv564;
  assign b_inv564 = ~b564;
  assign s564  = a564 ^ b564 ^ c564;
  assign sub564 = a564 ^ b_inv564 ^ c564;
  assign and564 = a564 & b564;
  assign or564  = a564 | b564;
  assign c565 = (a564 & b564) | (a564 & c564) | (b564 & c564);
  wire c_sub565;
  assign c_sub565 = (a564 & b_inv564) | (a564 & c564) | (b_inv564 & c564);
  wire s565, sub565, and565, or565;
  wire b_inv565;
  assign b_inv565 = ~b565;
  assign s565  = a565 ^ b565 ^ c565;
  assign sub565 = a565 ^ b_inv565 ^ c565;
  assign and565 = a565 & b565;
  assign or565  = a565 | b565;
  assign c566 = (a565 & b565) | (a565 & c565) | (b565 & c565);
  wire c_sub566;
  assign c_sub566 = (a565 & b_inv565) | (a565 & c565) | (b_inv565 & c565);
  wire s566, sub566, and566, or566;
  wire b_inv566;
  assign b_inv566 = ~b566;
  assign s566  = a566 ^ b566 ^ c566;
  assign sub566 = a566 ^ b_inv566 ^ c566;
  assign and566 = a566 & b566;
  assign or566  = a566 | b566;
  assign c567 = (a566 & b566) | (a566 & c566) | (b566 & c566);
  wire c_sub567;
  assign c_sub567 = (a566 & b_inv566) | (a566 & c566) | (b_inv566 & c566);
  wire s567, sub567, and567, or567;
  wire b_inv567;
  assign b_inv567 = ~b567;
  assign s567  = a567 ^ b567 ^ c567;
  assign sub567 = a567 ^ b_inv567 ^ c567;
  assign and567 = a567 & b567;
  assign or567  = a567 | b567;
  assign c568 = (a567 & b567) | (a567 & c567) | (b567 & c567);
  wire c_sub568;
  assign c_sub568 = (a567 & b_inv567) | (a567 & c567) | (b_inv567 & c567);
  wire s568, sub568, and568, or568;
  wire b_inv568;
  assign b_inv568 = ~b568;
  assign s568  = a568 ^ b568 ^ c568;
  assign sub568 = a568 ^ b_inv568 ^ c568;
  assign and568 = a568 & b568;
  assign or568  = a568 | b568;
  assign c569 = (a568 & b568) | (a568 & c568) | (b568 & c568);
  wire c_sub569;
  assign c_sub569 = (a568 & b_inv568) | (a568 & c568) | (b_inv568 & c568);
  wire s569, sub569, and569, or569;
  wire b_inv569;
  assign b_inv569 = ~b569;
  assign s569  = a569 ^ b569 ^ c569;
  assign sub569 = a569 ^ b_inv569 ^ c569;
  assign and569 = a569 & b569;
  assign or569  = a569 | b569;
  assign c570 = (a569 & b569) | (a569 & c569) | (b569 & c569);
  wire c_sub570;
  assign c_sub570 = (a569 & b_inv569) | (a569 & c569) | (b_inv569 & c569);
  wire s570, sub570, and570, or570;
  wire b_inv570;
  assign b_inv570 = ~b570;
  assign s570  = a570 ^ b570 ^ c570;
  assign sub570 = a570 ^ b_inv570 ^ c570;
  assign and570 = a570 & b570;
  assign or570  = a570 | b570;
  assign c571 = (a570 & b570) | (a570 & c570) | (b570 & c570);
  wire c_sub571;
  assign c_sub571 = (a570 & b_inv570) | (a570 & c570) | (b_inv570 & c570);
  wire s571, sub571, and571, or571;
  wire b_inv571;
  assign b_inv571 = ~b571;
  assign s571  = a571 ^ b571 ^ c571;
  assign sub571 = a571 ^ b_inv571 ^ c571;
  assign and571 = a571 & b571;
  assign or571  = a571 | b571;
  assign c572 = (a571 & b571) | (a571 & c571) | (b571 & c571);
  wire c_sub572;
  assign c_sub572 = (a571 & b_inv571) | (a571 & c571) | (b_inv571 & c571);
  wire s572, sub572, and572, or572;
  wire b_inv572;
  assign b_inv572 = ~b572;
  assign s572  = a572 ^ b572 ^ c572;
  assign sub572 = a572 ^ b_inv572 ^ c572;
  assign and572 = a572 & b572;
  assign or572  = a572 | b572;
  assign c573 = (a572 & b572) | (a572 & c572) | (b572 & c572);
  wire c_sub573;
  assign c_sub573 = (a572 & b_inv572) | (a572 & c572) | (b_inv572 & c572);
  wire s573, sub573, and573, or573;
  wire b_inv573;
  assign b_inv573 = ~b573;
  assign s573  = a573 ^ b573 ^ c573;
  assign sub573 = a573 ^ b_inv573 ^ c573;
  assign and573 = a573 & b573;
  assign or573  = a573 | b573;
  assign c574 = (a573 & b573) | (a573 & c573) | (b573 & c573);
  wire c_sub574;
  assign c_sub574 = (a573 & b_inv573) | (a573 & c573) | (b_inv573 & c573);
  wire s574, sub574, and574, or574;
  wire b_inv574;
  assign b_inv574 = ~b574;
  assign s574  = a574 ^ b574 ^ c574;
  assign sub574 = a574 ^ b_inv574 ^ c574;
  assign and574 = a574 & b574;
  assign or574  = a574 | b574;
  assign c575 = (a574 & b574) | (a574 & c574) | (b574 & c574);
  wire c_sub575;
  assign c_sub575 = (a574 & b_inv574) | (a574 & c574) | (b_inv574 & c574);
  wire s575, sub575, and575, or575;
  wire b_inv575;
  assign b_inv575 = ~b575;
  assign s575  = a575 ^ b575 ^ c575;
  assign sub575 = a575 ^ b_inv575 ^ c575;
  assign and575 = a575 & b575;
  assign or575  = a575 | b575;
  assign c576 = (a575 & b575) | (a575 & c575) | (b575 & c575);
  wire c_sub576;
  assign c_sub576 = (a575 & b_inv575) | (a575 & c575) | (b_inv575 & c575);
  wire s576, sub576, and576, or576;
  wire b_inv576;
  assign b_inv576 = ~b576;
  assign s576  = a576 ^ b576 ^ c576;
  assign sub576 = a576 ^ b_inv576 ^ c576;
  assign and576 = a576 & b576;
  assign or576  = a576 | b576;
  assign c577 = (a576 & b576) | (a576 & c576) | (b576 & c576);
  wire c_sub577;
  assign c_sub577 = (a576 & b_inv576) | (a576 & c576) | (b_inv576 & c576);
  wire s577, sub577, and577, or577;
  wire b_inv577;
  assign b_inv577 = ~b577;
  assign s577  = a577 ^ b577 ^ c577;
  assign sub577 = a577 ^ b_inv577 ^ c577;
  assign and577 = a577 & b577;
  assign or577  = a577 | b577;
  assign c578 = (a577 & b577) | (a577 & c577) | (b577 & c577);
  wire c_sub578;
  assign c_sub578 = (a577 & b_inv577) | (a577 & c577) | (b_inv577 & c577);
  wire s578, sub578, and578, or578;
  wire b_inv578;
  assign b_inv578 = ~b578;
  assign s578  = a578 ^ b578 ^ c578;
  assign sub578 = a578 ^ b_inv578 ^ c578;
  assign and578 = a578 & b578;
  assign or578  = a578 | b578;
  assign c579 = (a578 & b578) | (a578 & c578) | (b578 & c578);
  wire c_sub579;
  assign c_sub579 = (a578 & b_inv578) | (a578 & c578) | (b_inv578 & c578);
  wire s579, sub579, and579, or579;
  wire b_inv579;
  assign b_inv579 = ~b579;
  assign s579  = a579 ^ b579 ^ c579;
  assign sub579 = a579 ^ b_inv579 ^ c579;
  assign and579 = a579 & b579;
  assign or579  = a579 | b579;
  assign c580 = (a579 & b579) | (a579 & c579) | (b579 & c579);
  wire c_sub580;
  assign c_sub580 = (a579 & b_inv579) | (a579 & c579) | (b_inv579 & c579);
  wire s580, sub580, and580, or580;
  wire b_inv580;
  assign b_inv580 = ~b580;
  assign s580  = a580 ^ b580 ^ c580;
  assign sub580 = a580 ^ b_inv580 ^ c580;
  assign and580 = a580 & b580;
  assign or580  = a580 | b580;
  assign c581 = (a580 & b580) | (a580 & c580) | (b580 & c580);
  wire c_sub581;
  assign c_sub581 = (a580 & b_inv580) | (a580 & c580) | (b_inv580 & c580);
  wire s581, sub581, and581, or581;
  wire b_inv581;
  assign b_inv581 = ~b581;
  assign s581  = a581 ^ b581 ^ c581;
  assign sub581 = a581 ^ b_inv581 ^ c581;
  assign and581 = a581 & b581;
  assign or581  = a581 | b581;
  assign c582 = (a581 & b581) | (a581 & c581) | (b581 & c581);
  wire c_sub582;
  assign c_sub582 = (a581 & b_inv581) | (a581 & c581) | (b_inv581 & c581);
  wire s582, sub582, and582, or582;
  wire b_inv582;
  assign b_inv582 = ~b582;
  assign s582  = a582 ^ b582 ^ c582;
  assign sub582 = a582 ^ b_inv582 ^ c582;
  assign and582 = a582 & b582;
  assign or582  = a582 | b582;
  assign c583 = (a582 & b582) | (a582 & c582) | (b582 & c582);
  wire c_sub583;
  assign c_sub583 = (a582 & b_inv582) | (a582 & c582) | (b_inv582 & c582);
  wire s583, sub583, and583, or583;
  wire b_inv583;
  assign b_inv583 = ~b583;
  assign s583  = a583 ^ b583 ^ c583;
  assign sub583 = a583 ^ b_inv583 ^ c583;
  assign and583 = a583 & b583;
  assign or583  = a583 | b583;
  assign c584 = (a583 & b583) | (a583 & c583) | (b583 & c583);
  wire c_sub584;
  assign c_sub584 = (a583 & b_inv583) | (a583 & c583) | (b_inv583 & c583);
  wire s584, sub584, and584, or584;
  wire b_inv584;
  assign b_inv584 = ~b584;
  assign s584  = a584 ^ b584 ^ c584;
  assign sub584 = a584 ^ b_inv584 ^ c584;
  assign and584 = a584 & b584;
  assign or584  = a584 | b584;
  assign c585 = (a584 & b584) | (a584 & c584) | (b584 & c584);
  wire c_sub585;
  assign c_sub585 = (a584 & b_inv584) | (a584 & c584) | (b_inv584 & c584);
  wire s585, sub585, and585, or585;
  wire b_inv585;
  assign b_inv585 = ~b585;
  assign s585  = a585 ^ b585 ^ c585;
  assign sub585 = a585 ^ b_inv585 ^ c585;
  assign and585 = a585 & b585;
  assign or585  = a585 | b585;
  assign c586 = (a585 & b585) | (a585 & c585) | (b585 & c585);
  wire c_sub586;
  assign c_sub586 = (a585 & b_inv585) | (a585 & c585) | (b_inv585 & c585);
  wire s586, sub586, and586, or586;
  wire b_inv586;
  assign b_inv586 = ~b586;
  assign s586  = a586 ^ b586 ^ c586;
  assign sub586 = a586 ^ b_inv586 ^ c586;
  assign and586 = a586 & b586;
  assign or586  = a586 | b586;
  assign c587 = (a586 & b586) | (a586 & c586) | (b586 & c586);
  wire c_sub587;
  assign c_sub587 = (a586 & b_inv586) | (a586 & c586) | (b_inv586 & c586);
  wire s587, sub587, and587, or587;
  wire b_inv587;
  assign b_inv587 = ~b587;
  assign s587  = a587 ^ b587 ^ c587;
  assign sub587 = a587 ^ b_inv587 ^ c587;
  assign and587 = a587 & b587;
  assign or587  = a587 | b587;
  assign c588 = (a587 & b587) | (a587 & c587) | (b587 & c587);
  wire c_sub588;
  assign c_sub588 = (a587 & b_inv587) | (a587 & c587) | (b_inv587 & c587);
  wire s588, sub588, and588, or588;
  wire b_inv588;
  assign b_inv588 = ~b588;
  assign s588  = a588 ^ b588 ^ c588;
  assign sub588 = a588 ^ b_inv588 ^ c588;
  assign and588 = a588 & b588;
  assign or588  = a588 | b588;
  assign c589 = (a588 & b588) | (a588 & c588) | (b588 & c588);
  wire c_sub589;
  assign c_sub589 = (a588 & b_inv588) | (a588 & c588) | (b_inv588 & c588);
  wire s589, sub589, and589, or589;
  wire b_inv589;
  assign b_inv589 = ~b589;
  assign s589  = a589 ^ b589 ^ c589;
  assign sub589 = a589 ^ b_inv589 ^ c589;
  assign and589 = a589 & b589;
  assign or589  = a589 | b589;
  assign c590 = (a589 & b589) | (a589 & c589) | (b589 & c589);
  wire c_sub590;
  assign c_sub590 = (a589 & b_inv589) | (a589 & c589) | (b_inv589 & c589);
  wire s590, sub590, and590, or590;
  wire b_inv590;
  assign b_inv590 = ~b590;
  assign s590  = a590 ^ b590 ^ c590;
  assign sub590 = a590 ^ b_inv590 ^ c590;
  assign and590 = a590 & b590;
  assign or590  = a590 | b590;
  assign c591 = (a590 & b590) | (a590 & c590) | (b590 & c590);
  wire c_sub591;
  assign c_sub591 = (a590 & b_inv590) | (a590 & c590) | (b_inv590 & c590);
  wire s591, sub591, and591, or591;
  wire b_inv591;
  assign b_inv591 = ~b591;
  assign s591  = a591 ^ b591 ^ c591;
  assign sub591 = a591 ^ b_inv591 ^ c591;
  assign and591 = a591 & b591;
  assign or591  = a591 | b591;
  assign c592 = (a591 & b591) | (a591 & c591) | (b591 & c591);
  wire c_sub592;
  assign c_sub592 = (a591 & b_inv591) | (a591 & c591) | (b_inv591 & c591);
  wire s592, sub592, and592, or592;
  wire b_inv592;
  assign b_inv592 = ~b592;
  assign s592  = a592 ^ b592 ^ c592;
  assign sub592 = a592 ^ b_inv592 ^ c592;
  assign and592 = a592 & b592;
  assign or592  = a592 | b592;
  assign c593 = (a592 & b592) | (a592 & c592) | (b592 & c592);
  wire c_sub593;
  assign c_sub593 = (a592 & b_inv592) | (a592 & c592) | (b_inv592 & c592);
  wire s593, sub593, and593, or593;
  wire b_inv593;
  assign b_inv593 = ~b593;
  assign s593  = a593 ^ b593 ^ c593;
  assign sub593 = a593 ^ b_inv593 ^ c593;
  assign and593 = a593 & b593;
  assign or593  = a593 | b593;
  assign c594 = (a593 & b593) | (a593 & c593) | (b593 & c593);
  wire c_sub594;
  assign c_sub594 = (a593 & b_inv593) | (a593 & c593) | (b_inv593 & c593);
  wire s594, sub594, and594, or594;
  wire b_inv594;
  assign b_inv594 = ~b594;
  assign s594  = a594 ^ b594 ^ c594;
  assign sub594 = a594 ^ b_inv594 ^ c594;
  assign and594 = a594 & b594;
  assign or594  = a594 | b594;
  assign c595 = (a594 & b594) | (a594 & c594) | (b594 & c594);
  wire c_sub595;
  assign c_sub595 = (a594 & b_inv594) | (a594 & c594) | (b_inv594 & c594);
  wire s595, sub595, and595, or595;
  wire b_inv595;
  assign b_inv595 = ~b595;
  assign s595  = a595 ^ b595 ^ c595;
  assign sub595 = a595 ^ b_inv595 ^ c595;
  assign and595 = a595 & b595;
  assign or595  = a595 | b595;
  assign c596 = (a595 & b595) | (a595 & c595) | (b595 & c595);
  wire c_sub596;
  assign c_sub596 = (a595 & b_inv595) | (a595 & c595) | (b_inv595 & c595);
  wire s596, sub596, and596, or596;
  wire b_inv596;
  assign b_inv596 = ~b596;
  assign s596  = a596 ^ b596 ^ c596;
  assign sub596 = a596 ^ b_inv596 ^ c596;
  assign and596 = a596 & b596;
  assign or596  = a596 | b596;
  assign c597 = (a596 & b596) | (a596 & c596) | (b596 & c596);
  wire c_sub597;
  assign c_sub597 = (a596 & b_inv596) | (a596 & c596) | (b_inv596 & c596);
  wire s597, sub597, and597, or597;
  wire b_inv597;
  assign b_inv597 = ~b597;
  assign s597  = a597 ^ b597 ^ c597;
  assign sub597 = a597 ^ b_inv597 ^ c597;
  assign and597 = a597 & b597;
  assign or597  = a597 | b597;
  assign c598 = (a597 & b597) | (a597 & c597) | (b597 & c597);
  wire c_sub598;
  assign c_sub598 = (a597 & b_inv597) | (a597 & c597) | (b_inv597 & c597);
  wire s598, sub598, and598, or598;
  wire b_inv598;
  assign b_inv598 = ~b598;
  assign s598  = a598 ^ b598 ^ c598;
  assign sub598 = a598 ^ b_inv598 ^ c598;
  assign and598 = a598 & b598;
  assign or598  = a598 | b598;
  assign c599 = (a598 & b598) | (a598 & c598) | (b598 & c598);
  wire c_sub599;
  assign c_sub599 = (a598 & b_inv598) | (a598 & c598) | (b_inv598 & c598);
  wire s599, sub599, and599, or599;
  wire b_inv599;
  assign b_inv599 = ~b599;
  assign s599  = a599 ^ b599 ^ c599;
  assign sub599 = a599 ^ b_inv599 ^ c599;
  assign and599 = a599 & b599;
  assign or599  = a599 | b599;
  assign c600 = (a599 & b599) | (a599 & c599) | (b599 & c599);
  wire c_sub600;
  assign c_sub600 = (a599 & b_inv599) | (a599 & c599) | (b_inv599 & c599);
  wire s600, sub600, and600, or600;
  wire b_inv600;
  assign b_inv600 = ~b600;
  assign s600  = a600 ^ b600 ^ c600;
  assign sub600 = a600 ^ b_inv600 ^ c600;
  assign and600 = a600 & b600;
  assign or600  = a600 | b600;
  assign c601 = (a600 & b600) | (a600 & c600) | (b600 & c600);
  wire c_sub601;
  assign c_sub601 = (a600 & b_inv600) | (a600 & c600) | (b_inv600 & c600);
  wire s601, sub601, and601, or601;
  wire b_inv601;
  assign b_inv601 = ~b601;
  assign s601  = a601 ^ b601 ^ c601;
  assign sub601 = a601 ^ b_inv601 ^ c601;
  assign and601 = a601 & b601;
  assign or601  = a601 | b601;
  assign c602 = (a601 & b601) | (a601 & c601) | (b601 & c601);
  wire c_sub602;
  assign c_sub602 = (a601 & b_inv601) | (a601 & c601) | (b_inv601 & c601);
  wire s602, sub602, and602, or602;
  wire b_inv602;
  assign b_inv602 = ~b602;
  assign s602  = a602 ^ b602 ^ c602;
  assign sub602 = a602 ^ b_inv602 ^ c602;
  assign and602 = a602 & b602;
  assign or602  = a602 | b602;
  assign c603 = (a602 & b602) | (a602 & c602) | (b602 & c602);
  wire c_sub603;
  assign c_sub603 = (a602 & b_inv602) | (a602 & c602) | (b_inv602 & c602);
  wire s603, sub603, and603, or603;
  wire b_inv603;
  assign b_inv603 = ~b603;
  assign s603  = a603 ^ b603 ^ c603;
  assign sub603 = a603 ^ b_inv603 ^ c603;
  assign and603 = a603 & b603;
  assign or603  = a603 | b603;
  assign c604 = (a603 & b603) | (a603 & c603) | (b603 & c603);
  wire c_sub604;
  assign c_sub604 = (a603 & b_inv603) | (a603 & c603) | (b_inv603 & c603);
  wire s604, sub604, and604, or604;
  wire b_inv604;
  assign b_inv604 = ~b604;
  assign s604  = a604 ^ b604 ^ c604;
  assign sub604 = a604 ^ b_inv604 ^ c604;
  assign and604 = a604 & b604;
  assign or604  = a604 | b604;
  assign c605 = (a604 & b604) | (a604 & c604) | (b604 & c604);
  wire c_sub605;
  assign c_sub605 = (a604 & b_inv604) | (a604 & c604) | (b_inv604 & c604);
  wire s605, sub605, and605, or605;
  wire b_inv605;
  assign b_inv605 = ~b605;
  assign s605  = a605 ^ b605 ^ c605;
  assign sub605 = a605 ^ b_inv605 ^ c605;
  assign and605 = a605 & b605;
  assign or605  = a605 | b605;
  assign c606 = (a605 & b605) | (a605 & c605) | (b605 & c605);
  wire c_sub606;
  assign c_sub606 = (a605 & b_inv605) | (a605 & c605) | (b_inv605 & c605);
  wire s606, sub606, and606, or606;
  wire b_inv606;
  assign b_inv606 = ~b606;
  assign s606  = a606 ^ b606 ^ c606;
  assign sub606 = a606 ^ b_inv606 ^ c606;
  assign and606 = a606 & b606;
  assign or606  = a606 | b606;
  assign c607 = (a606 & b606) | (a606 & c606) | (b606 & c606);
  wire c_sub607;
  assign c_sub607 = (a606 & b_inv606) | (a606 & c606) | (b_inv606 & c606);
  wire s607, sub607, and607, or607;
  wire b_inv607;
  assign b_inv607 = ~b607;
  assign s607  = a607 ^ b607 ^ c607;
  assign sub607 = a607 ^ b_inv607 ^ c607;
  assign and607 = a607 & b607;
  assign or607  = a607 | b607;
  assign c608 = (a607 & b607) | (a607 & c607) | (b607 & c607);
  wire c_sub608;
  assign c_sub608 = (a607 & b_inv607) | (a607 & c607) | (b_inv607 & c607);
  wire s608, sub608, and608, or608;
  wire b_inv608;
  assign b_inv608 = ~b608;
  assign s608  = a608 ^ b608 ^ c608;
  assign sub608 = a608 ^ b_inv608 ^ c608;
  assign and608 = a608 & b608;
  assign or608  = a608 | b608;
  assign c609 = (a608 & b608) | (a608 & c608) | (b608 & c608);
  wire c_sub609;
  assign c_sub609 = (a608 & b_inv608) | (a608 & c608) | (b_inv608 & c608);
  wire s609, sub609, and609, or609;
  wire b_inv609;
  assign b_inv609 = ~b609;
  assign s609  = a609 ^ b609 ^ c609;
  assign sub609 = a609 ^ b_inv609 ^ c609;
  assign and609 = a609 & b609;
  assign or609  = a609 | b609;
  assign c610 = (a609 & b609) | (a609 & c609) | (b609 & c609);
  wire c_sub610;
  assign c_sub610 = (a609 & b_inv609) | (a609 & c609) | (b_inv609 & c609);
  wire s610, sub610, and610, or610;
  wire b_inv610;
  assign b_inv610 = ~b610;
  assign s610  = a610 ^ b610 ^ c610;
  assign sub610 = a610 ^ b_inv610 ^ c610;
  assign and610 = a610 & b610;
  assign or610  = a610 | b610;
  assign c611 = (a610 & b610) | (a610 & c610) | (b610 & c610);
  wire c_sub611;
  assign c_sub611 = (a610 & b_inv610) | (a610 & c610) | (b_inv610 & c610);
  wire s611, sub611, and611, or611;
  wire b_inv611;
  assign b_inv611 = ~b611;
  assign s611  = a611 ^ b611 ^ c611;
  assign sub611 = a611 ^ b_inv611 ^ c611;
  assign and611 = a611 & b611;
  assign or611  = a611 | b611;
  assign c612 = (a611 & b611) | (a611 & c611) | (b611 & c611);
  wire c_sub612;
  assign c_sub612 = (a611 & b_inv611) | (a611 & c611) | (b_inv611 & c611);
  wire s612, sub612, and612, or612;
  wire b_inv612;
  assign b_inv612 = ~b612;
  assign s612  = a612 ^ b612 ^ c612;
  assign sub612 = a612 ^ b_inv612 ^ c612;
  assign and612 = a612 & b612;
  assign or612  = a612 | b612;
  assign c613 = (a612 & b612) | (a612 & c612) | (b612 & c612);
  wire c_sub613;
  assign c_sub613 = (a612 & b_inv612) | (a612 & c612) | (b_inv612 & c612);
  wire s613, sub613, and613, or613;
  wire b_inv613;
  assign b_inv613 = ~b613;
  assign s613  = a613 ^ b613 ^ c613;
  assign sub613 = a613 ^ b_inv613 ^ c613;
  assign and613 = a613 & b613;
  assign or613  = a613 | b613;
  assign c614 = (a613 & b613) | (a613 & c613) | (b613 & c613);
  wire c_sub614;
  assign c_sub614 = (a613 & b_inv613) | (a613 & c613) | (b_inv613 & c613);
  wire s614, sub614, and614, or614;
  wire b_inv614;
  assign b_inv614 = ~b614;
  assign s614  = a614 ^ b614 ^ c614;
  assign sub614 = a614 ^ b_inv614 ^ c614;
  assign and614 = a614 & b614;
  assign or614  = a614 | b614;
  assign c615 = (a614 & b614) | (a614 & c614) | (b614 & c614);
  wire c_sub615;
  assign c_sub615 = (a614 & b_inv614) | (a614 & c614) | (b_inv614 & c614);
  wire s615, sub615, and615, or615;
  wire b_inv615;
  assign b_inv615 = ~b615;
  assign s615  = a615 ^ b615 ^ c615;
  assign sub615 = a615 ^ b_inv615 ^ c615;
  assign and615 = a615 & b615;
  assign or615  = a615 | b615;
  assign c616 = (a615 & b615) | (a615 & c615) | (b615 & c615);
  wire c_sub616;
  assign c_sub616 = (a615 & b_inv615) | (a615 & c615) | (b_inv615 & c615);
  wire s616, sub616, and616, or616;
  wire b_inv616;
  assign b_inv616 = ~b616;
  assign s616  = a616 ^ b616 ^ c616;
  assign sub616 = a616 ^ b_inv616 ^ c616;
  assign and616 = a616 & b616;
  assign or616  = a616 | b616;
  assign c617 = (a616 & b616) | (a616 & c616) | (b616 & c616);
  wire c_sub617;
  assign c_sub617 = (a616 & b_inv616) | (a616 & c616) | (b_inv616 & c616);
  wire s617, sub617, and617, or617;
  wire b_inv617;
  assign b_inv617 = ~b617;
  assign s617  = a617 ^ b617 ^ c617;
  assign sub617 = a617 ^ b_inv617 ^ c617;
  assign and617 = a617 & b617;
  assign or617  = a617 | b617;
  assign c618 = (a617 & b617) | (a617 & c617) | (b617 & c617);
  wire c_sub618;
  assign c_sub618 = (a617 & b_inv617) | (a617 & c617) | (b_inv617 & c617);
  wire s618, sub618, and618, or618;
  wire b_inv618;
  assign b_inv618 = ~b618;
  assign s618  = a618 ^ b618 ^ c618;
  assign sub618 = a618 ^ b_inv618 ^ c618;
  assign and618 = a618 & b618;
  assign or618  = a618 | b618;
  assign c619 = (a618 & b618) | (a618 & c618) | (b618 & c618);
  wire c_sub619;
  assign c_sub619 = (a618 & b_inv618) | (a618 & c618) | (b_inv618 & c618);
  wire s619, sub619, and619, or619;
  wire b_inv619;
  assign b_inv619 = ~b619;
  assign s619  = a619 ^ b619 ^ c619;
  assign sub619 = a619 ^ b_inv619 ^ c619;
  assign and619 = a619 & b619;
  assign or619  = a619 | b619;
  assign c620 = (a619 & b619) | (a619 & c619) | (b619 & c619);
  wire c_sub620;
  assign c_sub620 = (a619 & b_inv619) | (a619 & c619) | (b_inv619 & c619);
  wire s620, sub620, and620, or620;
  wire b_inv620;
  assign b_inv620 = ~b620;
  assign s620  = a620 ^ b620 ^ c620;
  assign sub620 = a620 ^ b_inv620 ^ c620;
  assign and620 = a620 & b620;
  assign or620  = a620 | b620;
  assign c621 = (a620 & b620) | (a620 & c620) | (b620 & c620);
  wire c_sub621;
  assign c_sub621 = (a620 & b_inv620) | (a620 & c620) | (b_inv620 & c620);
  wire s621, sub621, and621, or621;
  wire b_inv621;
  assign b_inv621 = ~b621;
  assign s621  = a621 ^ b621 ^ c621;
  assign sub621 = a621 ^ b_inv621 ^ c621;
  assign and621 = a621 & b621;
  assign or621  = a621 | b621;
  assign c622 = (a621 & b621) | (a621 & c621) | (b621 & c621);
  wire c_sub622;
  assign c_sub622 = (a621 & b_inv621) | (a621 & c621) | (b_inv621 & c621);
  wire s622, sub622, and622, or622;
  wire b_inv622;
  assign b_inv622 = ~b622;
  assign s622  = a622 ^ b622 ^ c622;
  assign sub622 = a622 ^ b_inv622 ^ c622;
  assign and622 = a622 & b622;
  assign or622  = a622 | b622;
  assign c623 = (a622 & b622) | (a622 & c622) | (b622 & c622);
  wire c_sub623;
  assign c_sub623 = (a622 & b_inv622) | (a622 & c622) | (b_inv622 & c622);
  wire s623, sub623, and623, or623;
  wire b_inv623;
  assign b_inv623 = ~b623;
  assign s623  = a623 ^ b623 ^ c623;
  assign sub623 = a623 ^ b_inv623 ^ c623;
  assign and623 = a623 & b623;
  assign or623  = a623 | b623;
  assign c624 = (a623 & b623) | (a623 & c623) | (b623 & c623);
  wire c_sub624;
  assign c_sub624 = (a623 & b_inv623) | (a623 & c623) | (b_inv623 & c623);
  wire s624, sub624, and624, or624;
  wire b_inv624;
  assign b_inv624 = ~b624;
  assign s624  = a624 ^ b624 ^ c624;
  assign sub624 = a624 ^ b_inv624 ^ c624;
  assign and624 = a624 & b624;
  assign or624  = a624 | b624;
  assign c625 = (a624 & b624) | (a624 & c624) | (b624 & c624);
  wire c_sub625;
  assign c_sub625 = (a624 & b_inv624) | (a624 & c624) | (b_inv624 & c624);
  wire s625, sub625, and625, or625;
  wire b_inv625;
  assign b_inv625 = ~b625;
  assign s625  = a625 ^ b625 ^ c625;
  assign sub625 = a625 ^ b_inv625 ^ c625;
  assign and625 = a625 & b625;
  assign or625  = a625 | b625;
  assign c626 = (a625 & b625) | (a625 & c625) | (b625 & c625);
  wire c_sub626;
  assign c_sub626 = (a625 & b_inv625) | (a625 & c625) | (b_inv625 & c625);
  wire s626, sub626, and626, or626;
  wire b_inv626;
  assign b_inv626 = ~b626;
  assign s626  = a626 ^ b626 ^ c626;
  assign sub626 = a626 ^ b_inv626 ^ c626;
  assign and626 = a626 & b626;
  assign or626  = a626 | b626;
  assign c627 = (a626 & b626) | (a626 & c626) | (b626 & c626);
  wire c_sub627;
  assign c_sub627 = (a626 & b_inv626) | (a626 & c626) | (b_inv626 & c626);
  wire s627, sub627, and627, or627;
  wire b_inv627;
  assign b_inv627 = ~b627;
  assign s627  = a627 ^ b627 ^ c627;
  assign sub627 = a627 ^ b_inv627 ^ c627;
  assign and627 = a627 & b627;
  assign or627  = a627 | b627;
  assign c628 = (a627 & b627) | (a627 & c627) | (b627 & c627);
  wire c_sub628;
  assign c_sub628 = (a627 & b_inv627) | (a627 & c627) | (b_inv627 & c627);
  wire s628, sub628, and628, or628;
  wire b_inv628;
  assign b_inv628 = ~b628;
  assign s628  = a628 ^ b628 ^ c628;
  assign sub628 = a628 ^ b_inv628 ^ c628;
  assign and628 = a628 & b628;
  assign or628  = a628 | b628;
  assign c629 = (a628 & b628) | (a628 & c628) | (b628 & c628);
  wire c_sub629;
  assign c_sub629 = (a628 & b_inv628) | (a628 & c628) | (b_inv628 & c628);
  wire s629, sub629, and629, or629;
  wire b_inv629;
  assign b_inv629 = ~b629;
  assign s629  = a629 ^ b629 ^ c629;
  assign sub629 = a629 ^ b_inv629 ^ c629;
  assign and629 = a629 & b629;
  assign or629  = a629 | b629;
  assign c630 = (a629 & b629) | (a629 & c629) | (b629 & c629);
  wire c_sub630;
  assign c_sub630 = (a629 & b_inv629) | (a629 & c629) | (b_inv629 & c629);
  wire s630, sub630, and630, or630;
  wire b_inv630;
  assign b_inv630 = ~b630;
  assign s630  = a630 ^ b630 ^ c630;
  assign sub630 = a630 ^ b_inv630 ^ c630;
  assign and630 = a630 & b630;
  assign or630  = a630 | b630;
  assign c631 = (a630 & b630) | (a630 & c630) | (b630 & c630);
  wire c_sub631;
  assign c_sub631 = (a630 & b_inv630) | (a630 & c630) | (b_inv630 & c630);
  wire s631, sub631, and631, or631;
  wire b_inv631;
  assign b_inv631 = ~b631;
  assign s631  = a631 ^ b631 ^ c631;
  assign sub631 = a631 ^ b_inv631 ^ c631;
  assign and631 = a631 & b631;
  assign or631  = a631 | b631;
  assign c632 = (a631 & b631) | (a631 & c631) | (b631 & c631);
  wire c_sub632;
  assign c_sub632 = (a631 & b_inv631) | (a631 & c631) | (b_inv631 & c631);
  wire s632, sub632, and632, or632;
  wire b_inv632;
  assign b_inv632 = ~b632;
  assign s632  = a632 ^ b632 ^ c632;
  assign sub632 = a632 ^ b_inv632 ^ c632;
  assign and632 = a632 & b632;
  assign or632  = a632 | b632;
  assign c633 = (a632 & b632) | (a632 & c632) | (b632 & c632);
  wire c_sub633;
  assign c_sub633 = (a632 & b_inv632) | (a632 & c632) | (b_inv632 & c632);
  wire s633, sub633, and633, or633;
  wire b_inv633;
  assign b_inv633 = ~b633;
  assign s633  = a633 ^ b633 ^ c633;
  assign sub633 = a633 ^ b_inv633 ^ c633;
  assign and633 = a633 & b633;
  assign or633  = a633 | b633;
  assign c634 = (a633 & b633) | (a633 & c633) | (b633 & c633);
  wire c_sub634;
  assign c_sub634 = (a633 & b_inv633) | (a633 & c633) | (b_inv633 & c633);
  wire s634, sub634, and634, or634;
  wire b_inv634;
  assign b_inv634 = ~b634;
  assign s634  = a634 ^ b634 ^ c634;
  assign sub634 = a634 ^ b_inv634 ^ c634;
  assign and634 = a634 & b634;
  assign or634  = a634 | b634;
  assign c635 = (a634 & b634) | (a634 & c634) | (b634 & c634);
  wire c_sub635;
  assign c_sub635 = (a634 & b_inv634) | (a634 & c634) | (b_inv634 & c634);
  wire s635, sub635, and635, or635;
  wire b_inv635;
  assign b_inv635 = ~b635;
  assign s635  = a635 ^ b635 ^ c635;
  assign sub635 = a635 ^ b_inv635 ^ c635;
  assign and635 = a635 & b635;
  assign or635  = a635 | b635;
  assign c636 = (a635 & b635) | (a635 & c635) | (b635 & c635);
  wire c_sub636;
  assign c_sub636 = (a635 & b_inv635) | (a635 & c635) | (b_inv635 & c635);
  wire s636, sub636, and636, or636;
  wire b_inv636;
  assign b_inv636 = ~b636;
  assign s636  = a636 ^ b636 ^ c636;
  assign sub636 = a636 ^ b_inv636 ^ c636;
  assign and636 = a636 & b636;
  assign or636  = a636 | b636;
  assign c637 = (a636 & b636) | (a636 & c636) | (b636 & c636);
  wire c_sub637;
  assign c_sub637 = (a636 & b_inv636) | (a636 & c636) | (b_inv636 & c636);
  wire s637, sub637, and637, or637;
  wire b_inv637;
  assign b_inv637 = ~b637;
  assign s637  = a637 ^ b637 ^ c637;
  assign sub637 = a637 ^ b_inv637 ^ c637;
  assign and637 = a637 & b637;
  assign or637  = a637 | b637;
  assign c638 = (a637 & b637) | (a637 & c637) | (b637 & c637);
  wire c_sub638;
  assign c_sub638 = (a637 & b_inv637) | (a637 & c637) | (b_inv637 & c637);
  wire s638, sub638, and638, or638;
  wire b_inv638;
  assign b_inv638 = ~b638;
  assign s638  = a638 ^ b638 ^ c638;
  assign sub638 = a638 ^ b_inv638 ^ c638;
  assign and638 = a638 & b638;
  assign or638  = a638 | b638;
  assign c639 = (a638 & b638) | (a638 & c638) | (b638 & c638);
  wire c_sub639;
  assign c_sub639 = (a638 & b_inv638) | (a638 & c638) | (b_inv638 & c638);
  wire s639, sub639, and639, or639;
  wire b_inv639;
  assign b_inv639 = ~b639;
  assign s639  = a639 ^ b639 ^ c639;
  assign sub639 = a639 ^ b_inv639 ^ c639;
  assign and639 = a639 & b639;
  assign or639  = a639 | b639;
  assign c640 = (a639 & b639) | (a639 & c639) | (b639 & c639);
  wire c_sub640;
  assign c_sub640 = (a639 & b_inv639) | (a639 & c639) | (b_inv639 & c639);
  wire s640, sub640, and640, or640;
  wire b_inv640;
  assign b_inv640 = ~b640;
  assign s640  = a640 ^ b640 ^ c640;
  assign sub640 = a640 ^ b_inv640 ^ c640;
  assign and640 = a640 & b640;
  assign or640  = a640 | b640;
  assign c641 = (a640 & b640) | (a640 & c640) | (b640 & c640);
  wire c_sub641;
  assign c_sub641 = (a640 & b_inv640) | (a640 & c640) | (b_inv640 & c640);
  wire s641, sub641, and641, or641;
  wire b_inv641;
  assign b_inv641 = ~b641;
  assign s641  = a641 ^ b641 ^ c641;
  assign sub641 = a641 ^ b_inv641 ^ c641;
  assign and641 = a641 & b641;
  assign or641  = a641 | b641;
  assign c642 = (a641 & b641) | (a641 & c641) | (b641 & c641);
  wire c_sub642;
  assign c_sub642 = (a641 & b_inv641) | (a641 & c641) | (b_inv641 & c641);
  wire s642, sub642, and642, or642;
  wire b_inv642;
  assign b_inv642 = ~b642;
  assign s642  = a642 ^ b642 ^ c642;
  assign sub642 = a642 ^ b_inv642 ^ c642;
  assign and642 = a642 & b642;
  assign or642  = a642 | b642;
  assign c643 = (a642 & b642) | (a642 & c642) | (b642 & c642);
  wire c_sub643;
  assign c_sub643 = (a642 & b_inv642) | (a642 & c642) | (b_inv642 & c642);
  wire s643, sub643, and643, or643;
  wire b_inv643;
  assign b_inv643 = ~b643;
  assign s643  = a643 ^ b643 ^ c643;
  assign sub643 = a643 ^ b_inv643 ^ c643;
  assign and643 = a643 & b643;
  assign or643  = a643 | b643;
  assign c644 = (a643 & b643) | (a643 & c643) | (b643 & c643);
  wire c_sub644;
  assign c_sub644 = (a643 & b_inv643) | (a643 & c643) | (b_inv643 & c643);
  wire s644, sub644, and644, or644;
  wire b_inv644;
  assign b_inv644 = ~b644;
  assign s644  = a644 ^ b644 ^ c644;
  assign sub644 = a644 ^ b_inv644 ^ c644;
  assign and644 = a644 & b644;
  assign or644  = a644 | b644;
  assign c645 = (a644 & b644) | (a644 & c644) | (b644 & c644);
  wire c_sub645;
  assign c_sub645 = (a644 & b_inv644) | (a644 & c644) | (b_inv644 & c644);
  wire s645, sub645, and645, or645;
  wire b_inv645;
  assign b_inv645 = ~b645;
  assign s645  = a645 ^ b645 ^ c645;
  assign sub645 = a645 ^ b_inv645 ^ c645;
  assign and645 = a645 & b645;
  assign or645  = a645 | b645;
  assign c646 = (a645 & b645) | (a645 & c645) | (b645 & c645);
  wire c_sub646;
  assign c_sub646 = (a645 & b_inv645) | (a645 & c645) | (b_inv645 & c645);
  wire s646, sub646, and646, or646;
  wire b_inv646;
  assign b_inv646 = ~b646;
  assign s646  = a646 ^ b646 ^ c646;
  assign sub646 = a646 ^ b_inv646 ^ c646;
  assign and646 = a646 & b646;
  assign or646  = a646 | b646;
  assign c647 = (a646 & b646) | (a646 & c646) | (b646 & c646);
  wire c_sub647;
  assign c_sub647 = (a646 & b_inv646) | (a646 & c646) | (b_inv646 & c646);
  wire s647, sub647, and647, or647;
  wire b_inv647;
  assign b_inv647 = ~b647;
  assign s647  = a647 ^ b647 ^ c647;
  assign sub647 = a647 ^ b_inv647 ^ c647;
  assign and647 = a647 & b647;
  assign or647  = a647 | b647;
  assign c648 = (a647 & b647) | (a647 & c647) | (b647 & c647);
  wire c_sub648;
  assign c_sub648 = (a647 & b_inv647) | (a647 & c647) | (b_inv647 & c647);
  wire s648, sub648, and648, or648;
  wire b_inv648;
  assign b_inv648 = ~b648;
  assign s648  = a648 ^ b648 ^ c648;
  assign sub648 = a648 ^ b_inv648 ^ c648;
  assign and648 = a648 & b648;
  assign or648  = a648 | b648;
  assign c649 = (a648 & b648) | (a648 & c648) | (b648 & c648);
  wire c_sub649;
  assign c_sub649 = (a648 & b_inv648) | (a648 & c648) | (b_inv648 & c648);
  wire s649, sub649, and649, or649;
  wire b_inv649;
  assign b_inv649 = ~b649;
  assign s649  = a649 ^ b649 ^ c649;
  assign sub649 = a649 ^ b_inv649 ^ c649;
  assign and649 = a649 & b649;
  assign or649  = a649 | b649;
  assign c650 = (a649 & b649) | (a649 & c649) | (b649 & c649);
  wire c_sub650;
  assign c_sub650 = (a649 & b_inv649) | (a649 & c649) | (b_inv649 & c649);
  wire s650, sub650, and650, or650;
  wire b_inv650;
  assign b_inv650 = ~b650;
  assign s650  = a650 ^ b650 ^ c650;
  assign sub650 = a650 ^ b_inv650 ^ c650;
  assign and650 = a650 & b650;
  assign or650  = a650 | b650;
  assign c651 = (a650 & b650) | (a650 & c650) | (b650 & c650);
  wire c_sub651;
  assign c_sub651 = (a650 & b_inv650) | (a650 & c650) | (b_inv650 & c650);
  wire s651, sub651, and651, or651;
  wire b_inv651;
  assign b_inv651 = ~b651;
  assign s651  = a651 ^ b651 ^ c651;
  assign sub651 = a651 ^ b_inv651 ^ c651;
  assign and651 = a651 & b651;
  assign or651  = a651 | b651;
  assign c652 = (a651 & b651) | (a651 & c651) | (b651 & c651);
  wire c_sub652;
  assign c_sub652 = (a651 & b_inv651) | (a651 & c651) | (b_inv651 & c651);
  wire s652, sub652, and652, or652;
  wire b_inv652;
  assign b_inv652 = ~b652;
  assign s652  = a652 ^ b652 ^ c652;
  assign sub652 = a652 ^ b_inv652 ^ c652;
  assign and652 = a652 & b652;
  assign or652  = a652 | b652;
  assign c653 = (a652 & b652) | (a652 & c652) | (b652 & c652);
  wire c_sub653;
  assign c_sub653 = (a652 & b_inv652) | (a652 & c652) | (b_inv652 & c652);
  wire s653, sub653, and653, or653;
  wire b_inv653;
  assign b_inv653 = ~b653;
  assign s653  = a653 ^ b653 ^ c653;
  assign sub653 = a653 ^ b_inv653 ^ c653;
  assign and653 = a653 & b653;
  assign or653  = a653 | b653;
  assign c654 = (a653 & b653) | (a653 & c653) | (b653 & c653);
  wire c_sub654;
  assign c_sub654 = (a653 & b_inv653) | (a653 & c653) | (b_inv653 & c653);
  wire s654, sub654, and654, or654;
  wire b_inv654;
  assign b_inv654 = ~b654;
  assign s654  = a654 ^ b654 ^ c654;
  assign sub654 = a654 ^ b_inv654 ^ c654;
  assign and654 = a654 & b654;
  assign or654  = a654 | b654;
  assign c655 = (a654 & b654) | (a654 & c654) | (b654 & c654);
  wire c_sub655;
  assign c_sub655 = (a654 & b_inv654) | (a654 & c654) | (b_inv654 & c654);
  wire s655, sub655, and655, or655;
  wire b_inv655;
  assign b_inv655 = ~b655;
  assign s655  = a655 ^ b655 ^ c655;
  assign sub655 = a655 ^ b_inv655 ^ c655;
  assign and655 = a655 & b655;
  assign or655  = a655 | b655;
  assign c656 = (a655 & b655) | (a655 & c655) | (b655 & c655);
  wire c_sub656;
  assign c_sub656 = (a655 & b_inv655) | (a655 & c655) | (b_inv655 & c655);
  wire s656, sub656, and656, or656;
  wire b_inv656;
  assign b_inv656 = ~b656;
  assign s656  = a656 ^ b656 ^ c656;
  assign sub656 = a656 ^ b_inv656 ^ c656;
  assign and656 = a656 & b656;
  assign or656  = a656 | b656;
  assign c657 = (a656 & b656) | (a656 & c656) | (b656 & c656);
  wire c_sub657;
  assign c_sub657 = (a656 & b_inv656) | (a656 & c656) | (b_inv656 & c656);
  wire s657, sub657, and657, or657;
  wire b_inv657;
  assign b_inv657 = ~b657;
  assign s657  = a657 ^ b657 ^ c657;
  assign sub657 = a657 ^ b_inv657 ^ c657;
  assign and657 = a657 & b657;
  assign or657  = a657 | b657;
  assign c658 = (a657 & b657) | (a657 & c657) | (b657 & c657);
  wire c_sub658;
  assign c_sub658 = (a657 & b_inv657) | (a657 & c657) | (b_inv657 & c657);
  wire s658, sub658, and658, or658;
  wire b_inv658;
  assign b_inv658 = ~b658;
  assign s658  = a658 ^ b658 ^ c658;
  assign sub658 = a658 ^ b_inv658 ^ c658;
  assign and658 = a658 & b658;
  assign or658  = a658 | b658;
  assign c659 = (a658 & b658) | (a658 & c658) | (b658 & c658);
  wire c_sub659;
  assign c_sub659 = (a658 & b_inv658) | (a658 & c658) | (b_inv658 & c658);
  wire s659, sub659, and659, or659;
  wire b_inv659;
  assign b_inv659 = ~b659;
  assign s659  = a659 ^ b659 ^ c659;
  assign sub659 = a659 ^ b_inv659 ^ c659;
  assign and659 = a659 & b659;
  assign or659  = a659 | b659;
  assign c660 = (a659 & b659) | (a659 & c659) | (b659 & c659);
  wire c_sub660;
  assign c_sub660 = (a659 & b_inv659) | (a659 & c659) | (b_inv659 & c659);
  wire s660, sub660, and660, or660;
  wire b_inv660;
  assign b_inv660 = ~b660;
  assign s660  = a660 ^ b660 ^ c660;
  assign sub660 = a660 ^ b_inv660 ^ c660;
  assign and660 = a660 & b660;
  assign or660  = a660 | b660;
  assign c661 = (a660 & b660) | (a660 & c660) | (b660 & c660);
  wire c_sub661;
  assign c_sub661 = (a660 & b_inv660) | (a660 & c660) | (b_inv660 & c660);
  wire s661, sub661, and661, or661;
  wire b_inv661;
  assign b_inv661 = ~b661;
  assign s661  = a661 ^ b661 ^ c661;
  assign sub661 = a661 ^ b_inv661 ^ c661;
  assign and661 = a661 & b661;
  assign or661  = a661 | b661;
  assign c662 = (a661 & b661) | (a661 & c661) | (b661 & c661);
  wire c_sub662;
  assign c_sub662 = (a661 & b_inv661) | (a661 & c661) | (b_inv661 & c661);
  wire s662, sub662, and662, or662;
  wire b_inv662;
  assign b_inv662 = ~b662;
  assign s662  = a662 ^ b662 ^ c662;
  assign sub662 = a662 ^ b_inv662 ^ c662;
  assign and662 = a662 & b662;
  assign or662  = a662 | b662;
  assign c663 = (a662 & b662) | (a662 & c662) | (b662 & c662);
  wire c_sub663;
  assign c_sub663 = (a662 & b_inv662) | (a662 & c662) | (b_inv662 & c662);
  wire s663, sub663, and663, or663;
  wire b_inv663;
  assign b_inv663 = ~b663;
  assign s663  = a663 ^ b663 ^ c663;
  assign sub663 = a663 ^ b_inv663 ^ c663;
  assign and663 = a663 & b663;
  assign or663  = a663 | b663;
  assign c664 = (a663 & b663) | (a663 & c663) | (b663 & c663);
  wire c_sub664;
  assign c_sub664 = (a663 & b_inv663) | (a663 & c663) | (b_inv663 & c663);
  wire s664, sub664, and664, or664;
  wire b_inv664;
  assign b_inv664 = ~b664;
  assign s664  = a664 ^ b664 ^ c664;
  assign sub664 = a664 ^ b_inv664 ^ c664;
  assign and664 = a664 & b664;
  assign or664  = a664 | b664;
  assign c665 = (a664 & b664) | (a664 & c664) | (b664 & c664);
  wire c_sub665;
  assign c_sub665 = (a664 & b_inv664) | (a664 & c664) | (b_inv664 & c664);
  wire s665, sub665, and665, or665;
  wire b_inv665;
  assign b_inv665 = ~b665;
  assign s665  = a665 ^ b665 ^ c665;
  assign sub665 = a665 ^ b_inv665 ^ c665;
  assign and665 = a665 & b665;
  assign or665  = a665 | b665;
  assign c666 = (a665 & b665) | (a665 & c665) | (b665 & c665);
  wire c_sub666;
  assign c_sub666 = (a665 & b_inv665) | (a665 & c665) | (b_inv665 & c665);
  wire s666, sub666, and666, or666;
  wire b_inv666;
  assign b_inv666 = ~b666;
  assign s666  = a666 ^ b666 ^ c666;
  assign sub666 = a666 ^ b_inv666 ^ c666;
  assign and666 = a666 & b666;
  assign or666  = a666 | b666;
  assign c667 = (a666 & b666) | (a666 & c666) | (b666 & c666);
  wire c_sub667;
  assign c_sub667 = (a666 & b_inv666) | (a666 & c666) | (b_inv666 & c666);
  wire s667, sub667, and667, or667;
  wire b_inv667;
  assign b_inv667 = ~b667;
  assign s667  = a667 ^ b667 ^ c667;
  assign sub667 = a667 ^ b_inv667 ^ c667;
  assign and667 = a667 & b667;
  assign or667  = a667 | b667;
  assign c668 = (a667 & b667) | (a667 & c667) | (b667 & c667);
  wire c_sub668;
  assign c_sub668 = (a667 & b_inv667) | (a667 & c667) | (b_inv667 & c667);
  wire s668, sub668, and668, or668;
  wire b_inv668;
  assign b_inv668 = ~b668;
  assign s668  = a668 ^ b668 ^ c668;
  assign sub668 = a668 ^ b_inv668 ^ c668;
  assign and668 = a668 & b668;
  assign or668  = a668 | b668;
  assign c669 = (a668 & b668) | (a668 & c668) | (b668 & c668);
  wire c_sub669;
  assign c_sub669 = (a668 & b_inv668) | (a668 & c668) | (b_inv668 & c668);
  wire s669, sub669, and669, or669;
  wire b_inv669;
  assign b_inv669 = ~b669;
  assign s669  = a669 ^ b669 ^ c669;
  assign sub669 = a669 ^ b_inv669 ^ c669;
  assign and669 = a669 & b669;
  assign or669  = a669 | b669;
  assign c670 = (a669 & b669) | (a669 & c669) | (b669 & c669);
  wire c_sub670;
  assign c_sub670 = (a669 & b_inv669) | (a669 & c669) | (b_inv669 & c669);
  wire s670, sub670, and670, or670;
  wire b_inv670;
  assign b_inv670 = ~b670;
  assign s670  = a670 ^ b670 ^ c670;
  assign sub670 = a670 ^ b_inv670 ^ c670;
  assign and670 = a670 & b670;
  assign or670  = a670 | b670;
  assign c671 = (a670 & b670) | (a670 & c670) | (b670 & c670);
  wire c_sub671;
  assign c_sub671 = (a670 & b_inv670) | (a670 & c670) | (b_inv670 & c670);
  wire s671, sub671, and671, or671;
  wire b_inv671;
  assign b_inv671 = ~b671;
  assign s671  = a671 ^ b671 ^ c671;
  assign sub671 = a671 ^ b_inv671 ^ c671;
  assign and671 = a671 & b671;
  assign or671  = a671 | b671;
  assign c672 = (a671 & b671) | (a671 & c671) | (b671 & c671);
  wire c_sub672;
  assign c_sub672 = (a671 & b_inv671) | (a671 & c671) | (b_inv671 & c671);
  wire s672, sub672, and672, or672;
  wire b_inv672;
  assign b_inv672 = ~b672;
  assign s672  = a672 ^ b672 ^ c672;
  assign sub672 = a672 ^ b_inv672 ^ c672;
  assign and672 = a672 & b672;
  assign or672  = a672 | b672;
  assign c673 = (a672 & b672) | (a672 & c672) | (b672 & c672);
  wire c_sub673;
  assign c_sub673 = (a672 & b_inv672) | (a672 & c672) | (b_inv672 & c672);
  wire s673, sub673, and673, or673;
  wire b_inv673;
  assign b_inv673 = ~b673;
  assign s673  = a673 ^ b673 ^ c673;
  assign sub673 = a673 ^ b_inv673 ^ c673;
  assign and673 = a673 & b673;
  assign or673  = a673 | b673;
  assign c674 = (a673 & b673) | (a673 & c673) | (b673 & c673);
  wire c_sub674;
  assign c_sub674 = (a673 & b_inv673) | (a673 & c673) | (b_inv673 & c673);
  wire s674, sub674, and674, or674;
  wire b_inv674;
  assign b_inv674 = ~b674;
  assign s674  = a674 ^ b674 ^ c674;
  assign sub674 = a674 ^ b_inv674 ^ c674;
  assign and674 = a674 & b674;
  assign or674  = a674 | b674;
  assign c675 = (a674 & b674) | (a674 & c674) | (b674 & c674);
  wire c_sub675;
  assign c_sub675 = (a674 & b_inv674) | (a674 & c674) | (b_inv674 & c674);
  wire s675, sub675, and675, or675;
  wire b_inv675;
  assign b_inv675 = ~b675;
  assign s675  = a675 ^ b675 ^ c675;
  assign sub675 = a675 ^ b_inv675 ^ c675;
  assign and675 = a675 & b675;
  assign or675  = a675 | b675;
  assign c676 = (a675 & b675) | (a675 & c675) | (b675 & c675);
  wire c_sub676;
  assign c_sub676 = (a675 & b_inv675) | (a675 & c675) | (b_inv675 & c675);
  wire s676, sub676, and676, or676;
  wire b_inv676;
  assign b_inv676 = ~b676;
  assign s676  = a676 ^ b676 ^ c676;
  assign sub676 = a676 ^ b_inv676 ^ c676;
  assign and676 = a676 & b676;
  assign or676  = a676 | b676;
  assign c677 = (a676 & b676) | (a676 & c676) | (b676 & c676);
  wire c_sub677;
  assign c_sub677 = (a676 & b_inv676) | (a676 & c676) | (b_inv676 & c676);
  wire s677, sub677, and677, or677;
  wire b_inv677;
  assign b_inv677 = ~b677;
  assign s677  = a677 ^ b677 ^ c677;
  assign sub677 = a677 ^ b_inv677 ^ c677;
  assign and677 = a677 & b677;
  assign or677  = a677 | b677;
  assign c678 = (a677 & b677) | (a677 & c677) | (b677 & c677);
  wire c_sub678;
  assign c_sub678 = (a677 & b_inv677) | (a677 & c677) | (b_inv677 & c677);
  wire s678, sub678, and678, or678;
  wire b_inv678;
  assign b_inv678 = ~b678;
  assign s678  = a678 ^ b678 ^ c678;
  assign sub678 = a678 ^ b_inv678 ^ c678;
  assign and678 = a678 & b678;
  assign or678  = a678 | b678;
  assign c679 = (a678 & b678) | (a678 & c678) | (b678 & c678);
  wire c_sub679;
  assign c_sub679 = (a678 & b_inv678) | (a678 & c678) | (b_inv678 & c678);
  wire s679, sub679, and679, or679;
  wire b_inv679;
  assign b_inv679 = ~b679;
  assign s679  = a679 ^ b679 ^ c679;
  assign sub679 = a679 ^ b_inv679 ^ c679;
  assign and679 = a679 & b679;
  assign or679  = a679 | b679;
  assign c680 = (a679 & b679) | (a679 & c679) | (b679 & c679);
  wire c_sub680;
  assign c_sub680 = (a679 & b_inv679) | (a679 & c679) | (b_inv679 & c679);
  wire s680, sub680, and680, or680;
  wire b_inv680;
  assign b_inv680 = ~b680;
  assign s680  = a680 ^ b680 ^ c680;
  assign sub680 = a680 ^ b_inv680 ^ c680;
  assign and680 = a680 & b680;
  assign or680  = a680 | b680;
  assign c681 = (a680 & b680) | (a680 & c680) | (b680 & c680);
  wire c_sub681;
  assign c_sub681 = (a680 & b_inv680) | (a680 & c680) | (b_inv680 & c680);
  wire s681, sub681, and681, or681;
  wire b_inv681;
  assign b_inv681 = ~b681;
  assign s681  = a681 ^ b681 ^ c681;
  assign sub681 = a681 ^ b_inv681 ^ c681;
  assign and681 = a681 & b681;
  assign or681  = a681 | b681;
  assign c682 = (a681 & b681) | (a681 & c681) | (b681 & c681);
  wire c_sub682;
  assign c_sub682 = (a681 & b_inv681) | (a681 & c681) | (b_inv681 & c681);
  wire s682, sub682, and682, or682;
  wire b_inv682;
  assign b_inv682 = ~b682;
  assign s682  = a682 ^ b682 ^ c682;
  assign sub682 = a682 ^ b_inv682 ^ c682;
  assign and682 = a682 & b682;
  assign or682  = a682 | b682;
  assign c683 = (a682 & b682) | (a682 & c682) | (b682 & c682);
  wire c_sub683;
  assign c_sub683 = (a682 & b_inv682) | (a682 & c682) | (b_inv682 & c682);
  wire s683, sub683, and683, or683;
  wire b_inv683;
  assign b_inv683 = ~b683;
  assign s683  = a683 ^ b683 ^ c683;
  assign sub683 = a683 ^ b_inv683 ^ c683;
  assign and683 = a683 & b683;
  assign or683  = a683 | b683;
  assign c684 = (a683 & b683) | (a683 & c683) | (b683 & c683);
  wire c_sub684;
  assign c_sub684 = (a683 & b_inv683) | (a683 & c683) | (b_inv683 & c683);
  wire s684, sub684, and684, or684;
  wire b_inv684;
  assign b_inv684 = ~b684;
  assign s684  = a684 ^ b684 ^ c684;
  assign sub684 = a684 ^ b_inv684 ^ c684;
  assign and684 = a684 & b684;
  assign or684  = a684 | b684;
  assign c685 = (a684 & b684) | (a684 & c684) | (b684 & c684);
  wire c_sub685;
  assign c_sub685 = (a684 & b_inv684) | (a684 & c684) | (b_inv684 & c684);
  wire s685, sub685, and685, or685;
  wire b_inv685;
  assign b_inv685 = ~b685;
  assign s685  = a685 ^ b685 ^ c685;
  assign sub685 = a685 ^ b_inv685 ^ c685;
  assign and685 = a685 & b685;
  assign or685  = a685 | b685;
  assign c686 = (a685 & b685) | (a685 & c685) | (b685 & c685);
  wire c_sub686;
  assign c_sub686 = (a685 & b_inv685) | (a685 & c685) | (b_inv685 & c685);
  wire s686, sub686, and686, or686;
  wire b_inv686;
  assign b_inv686 = ~b686;
  assign s686  = a686 ^ b686 ^ c686;
  assign sub686 = a686 ^ b_inv686 ^ c686;
  assign and686 = a686 & b686;
  assign or686  = a686 | b686;
  assign c687 = (a686 & b686) | (a686 & c686) | (b686 & c686);
  wire c_sub687;
  assign c_sub687 = (a686 & b_inv686) | (a686 & c686) | (b_inv686 & c686);
  wire s687, sub687, and687, or687;
  wire b_inv687;
  assign b_inv687 = ~b687;
  assign s687  = a687 ^ b687 ^ c687;
  assign sub687 = a687 ^ b_inv687 ^ c687;
  assign and687 = a687 & b687;
  assign or687  = a687 | b687;
  assign c688 = (a687 & b687) | (a687 & c687) | (b687 & c687);
  wire c_sub688;
  assign c_sub688 = (a687 & b_inv687) | (a687 & c687) | (b_inv687 & c687);
  wire s688, sub688, and688, or688;
  wire b_inv688;
  assign b_inv688 = ~b688;
  assign s688  = a688 ^ b688 ^ c688;
  assign sub688 = a688 ^ b_inv688 ^ c688;
  assign and688 = a688 & b688;
  assign or688  = a688 | b688;
  assign c689 = (a688 & b688) | (a688 & c688) | (b688 & c688);
  wire c_sub689;
  assign c_sub689 = (a688 & b_inv688) | (a688 & c688) | (b_inv688 & c688);
  wire s689, sub689, and689, or689;
  wire b_inv689;
  assign b_inv689 = ~b689;
  assign s689  = a689 ^ b689 ^ c689;
  assign sub689 = a689 ^ b_inv689 ^ c689;
  assign and689 = a689 & b689;
  assign or689  = a689 | b689;
  assign c690 = (a689 & b689) | (a689 & c689) | (b689 & c689);
  wire c_sub690;
  assign c_sub690 = (a689 & b_inv689) | (a689 & c689) | (b_inv689 & c689);
  wire s690, sub690, and690, or690;
  wire b_inv690;
  assign b_inv690 = ~b690;
  assign s690  = a690 ^ b690 ^ c690;
  assign sub690 = a690 ^ b_inv690 ^ c690;
  assign and690 = a690 & b690;
  assign or690  = a690 | b690;
  assign c691 = (a690 & b690) | (a690 & c690) | (b690 & c690);
  wire c_sub691;
  assign c_sub691 = (a690 & b_inv690) | (a690 & c690) | (b_inv690 & c690);
  wire s691, sub691, and691, or691;
  wire b_inv691;
  assign b_inv691 = ~b691;
  assign s691  = a691 ^ b691 ^ c691;
  assign sub691 = a691 ^ b_inv691 ^ c691;
  assign and691 = a691 & b691;
  assign or691  = a691 | b691;
  assign c692 = (a691 & b691) | (a691 & c691) | (b691 & c691);
  wire c_sub692;
  assign c_sub692 = (a691 & b_inv691) | (a691 & c691) | (b_inv691 & c691);
  wire s692, sub692, and692, or692;
  wire b_inv692;
  assign b_inv692 = ~b692;
  assign s692  = a692 ^ b692 ^ c692;
  assign sub692 = a692 ^ b_inv692 ^ c692;
  assign and692 = a692 & b692;
  assign or692  = a692 | b692;
  assign c693 = (a692 & b692) | (a692 & c692) | (b692 & c692);
  wire c_sub693;
  assign c_sub693 = (a692 & b_inv692) | (a692 & c692) | (b_inv692 & c692);
  wire s693, sub693, and693, or693;
  wire b_inv693;
  assign b_inv693 = ~b693;
  assign s693  = a693 ^ b693 ^ c693;
  assign sub693 = a693 ^ b_inv693 ^ c693;
  assign and693 = a693 & b693;
  assign or693  = a693 | b693;
  assign c694 = (a693 & b693) | (a693 & c693) | (b693 & c693);
  wire c_sub694;
  assign c_sub694 = (a693 & b_inv693) | (a693 & c693) | (b_inv693 & c693);
  wire s694, sub694, and694, or694;
  wire b_inv694;
  assign b_inv694 = ~b694;
  assign s694  = a694 ^ b694 ^ c694;
  assign sub694 = a694 ^ b_inv694 ^ c694;
  assign and694 = a694 & b694;
  assign or694  = a694 | b694;
  assign c695 = (a694 & b694) | (a694 & c694) | (b694 & c694);
  wire c_sub695;
  assign c_sub695 = (a694 & b_inv694) | (a694 & c694) | (b_inv694 & c694);
  wire s695, sub695, and695, or695;
  wire b_inv695;
  assign b_inv695 = ~b695;
  assign s695  = a695 ^ b695 ^ c695;
  assign sub695 = a695 ^ b_inv695 ^ c695;
  assign and695 = a695 & b695;
  assign or695  = a695 | b695;
  assign c696 = (a695 & b695) | (a695 & c695) | (b695 & c695);
  wire c_sub696;
  assign c_sub696 = (a695 & b_inv695) | (a695 & c695) | (b_inv695 & c695);
  wire s696, sub696, and696, or696;
  wire b_inv696;
  assign b_inv696 = ~b696;
  assign s696  = a696 ^ b696 ^ c696;
  assign sub696 = a696 ^ b_inv696 ^ c696;
  assign and696 = a696 & b696;
  assign or696  = a696 | b696;
  assign c697 = (a696 & b696) | (a696 & c696) | (b696 & c696);
  wire c_sub697;
  assign c_sub697 = (a696 & b_inv696) | (a696 & c696) | (b_inv696 & c696);
  wire s697, sub697, and697, or697;
  wire b_inv697;
  assign b_inv697 = ~b697;
  assign s697  = a697 ^ b697 ^ c697;
  assign sub697 = a697 ^ b_inv697 ^ c697;
  assign and697 = a697 & b697;
  assign or697  = a697 | b697;
  assign c698 = (a697 & b697) | (a697 & c697) | (b697 & c697);
  wire c_sub698;
  assign c_sub698 = (a697 & b_inv697) | (a697 & c697) | (b_inv697 & c697);
  wire s698, sub698, and698, or698;
  wire b_inv698;
  assign b_inv698 = ~b698;
  assign s698  = a698 ^ b698 ^ c698;
  assign sub698 = a698 ^ b_inv698 ^ c698;
  assign and698 = a698 & b698;
  assign or698  = a698 | b698;
  assign c699 = (a698 & b698) | (a698 & c698) | (b698 & c698);
  wire c_sub699;
  assign c_sub699 = (a698 & b_inv698) | (a698 & c698) | (b_inv698 & c698);
  wire s699, sub699, and699, or699;
  wire b_inv699;
  assign b_inv699 = ~b699;
  assign s699  = a699 ^ b699 ^ c699;
  assign sub699 = a699 ^ b_inv699 ^ c699;
  assign and699 = a699 & b699;
  assign or699  = a699 | b699;
  assign c700 = (a699 & b699) | (a699 & c699) | (b699 & c699);
  wire c_sub700;
  assign c_sub700 = (a699 & b_inv699) | (a699 & c699) | (b_inv699 & c699);
  wire s700, sub700, and700, or700;
  wire b_inv700;
  assign b_inv700 = ~b700;
  assign s700  = a700 ^ b700 ^ c700;
  assign sub700 = a700 ^ b_inv700 ^ c700;
  assign and700 = a700 & b700;
  assign or700  = a700 | b700;
  assign c701 = (a700 & b700) | (a700 & c700) | (b700 & c700);
  wire c_sub701;
  assign c_sub701 = (a700 & b_inv700) | (a700 & c700) | (b_inv700 & c700);
  wire s701, sub701, and701, or701;
  wire b_inv701;
  assign b_inv701 = ~b701;
  assign s701  = a701 ^ b701 ^ c701;
  assign sub701 = a701 ^ b_inv701 ^ c701;
  assign and701 = a701 & b701;
  assign or701  = a701 | b701;
  assign c702 = (a701 & b701) | (a701 & c701) | (b701 & c701);
  wire c_sub702;
  assign c_sub702 = (a701 & b_inv701) | (a701 & c701) | (b_inv701 & c701);
  wire s702, sub702, and702, or702;
  wire b_inv702;
  assign b_inv702 = ~b702;
  assign s702  = a702 ^ b702 ^ c702;
  assign sub702 = a702 ^ b_inv702 ^ c702;
  assign and702 = a702 & b702;
  assign or702  = a702 | b702;
  assign c703 = (a702 & b702) | (a702 & c702) | (b702 & c702);
  wire c_sub703;
  assign c_sub703 = (a702 & b_inv702) | (a702 & c702) | (b_inv702 & c702);
  wire s703, sub703, and703, or703;
  wire b_inv703;
  assign b_inv703 = ~b703;
  assign s703  = a703 ^ b703 ^ c703;
  assign sub703 = a703 ^ b_inv703 ^ c703;
  assign and703 = a703 & b703;
  assign or703  = a703 | b703;
  assign c704 = (a703 & b703) | (a703 & c703) | (b703 & c703);
  wire c_sub704;
  assign c_sub704 = (a703 & b_inv703) | (a703 & c703) | (b_inv703 & c703);
  wire s704, sub704, and704, or704;
  wire b_inv704;
  assign b_inv704 = ~b704;
  assign s704  = a704 ^ b704 ^ c704;
  assign sub704 = a704 ^ b_inv704 ^ c704;
  assign and704 = a704 & b704;
  assign or704  = a704 | b704;
  assign c705 = (a704 & b704) | (a704 & c704) | (b704 & c704);
  wire c_sub705;
  assign c_sub705 = (a704 & b_inv704) | (a704 & c704) | (b_inv704 & c704);
  wire s705, sub705, and705, or705;
  wire b_inv705;
  assign b_inv705 = ~b705;
  assign s705  = a705 ^ b705 ^ c705;
  assign sub705 = a705 ^ b_inv705 ^ c705;
  assign and705 = a705 & b705;
  assign or705  = a705 | b705;
  assign c706 = (a705 & b705) | (a705 & c705) | (b705 & c705);
  wire c_sub706;
  assign c_sub706 = (a705 & b_inv705) | (a705 & c705) | (b_inv705 & c705);
  wire s706, sub706, and706, or706;
  wire b_inv706;
  assign b_inv706 = ~b706;
  assign s706  = a706 ^ b706 ^ c706;
  assign sub706 = a706 ^ b_inv706 ^ c706;
  assign and706 = a706 & b706;
  assign or706  = a706 | b706;
  assign c707 = (a706 & b706) | (a706 & c706) | (b706 & c706);
  wire c_sub707;
  assign c_sub707 = (a706 & b_inv706) | (a706 & c706) | (b_inv706 & c706);
  wire s707, sub707, and707, or707;
  wire b_inv707;
  assign b_inv707 = ~b707;
  assign s707  = a707 ^ b707 ^ c707;
  assign sub707 = a707 ^ b_inv707 ^ c707;
  assign and707 = a707 & b707;
  assign or707  = a707 | b707;
  assign c708 = (a707 & b707) | (a707 & c707) | (b707 & c707);
  wire c_sub708;
  assign c_sub708 = (a707 & b_inv707) | (a707 & c707) | (b_inv707 & c707);
  wire s708, sub708, and708, or708;
  wire b_inv708;
  assign b_inv708 = ~b708;
  assign s708  = a708 ^ b708 ^ c708;
  assign sub708 = a708 ^ b_inv708 ^ c708;
  assign and708 = a708 & b708;
  assign or708  = a708 | b708;
  assign c709 = (a708 & b708) | (a708 & c708) | (b708 & c708);
  wire c_sub709;
  assign c_sub709 = (a708 & b_inv708) | (a708 & c708) | (b_inv708 & c708);
  wire s709, sub709, and709, or709;
  wire b_inv709;
  assign b_inv709 = ~b709;
  assign s709  = a709 ^ b709 ^ c709;
  assign sub709 = a709 ^ b_inv709 ^ c709;
  assign and709 = a709 & b709;
  assign or709  = a709 | b709;
  assign c710 = (a709 & b709) | (a709 & c709) | (b709 & c709);
  wire c_sub710;
  assign c_sub710 = (a709 & b_inv709) | (a709 & c709) | (b_inv709 & c709);
  wire s710, sub710, and710, or710;
  wire b_inv710;
  assign b_inv710 = ~b710;
  assign s710  = a710 ^ b710 ^ c710;
  assign sub710 = a710 ^ b_inv710 ^ c710;
  assign and710 = a710 & b710;
  assign or710  = a710 | b710;
  assign c711 = (a710 & b710) | (a710 & c710) | (b710 & c710);
  wire c_sub711;
  assign c_sub711 = (a710 & b_inv710) | (a710 & c710) | (b_inv710 & c710);
  wire s711, sub711, and711, or711;
  wire b_inv711;
  assign b_inv711 = ~b711;
  assign s711  = a711 ^ b711 ^ c711;
  assign sub711 = a711 ^ b_inv711 ^ c711;
  assign and711 = a711 & b711;
  assign or711  = a711 | b711;
  assign c712 = (a711 & b711) | (a711 & c711) | (b711 & c711);
  wire c_sub712;
  assign c_sub712 = (a711 & b_inv711) | (a711 & c711) | (b_inv711 & c711);
  wire s712, sub712, and712, or712;
  wire b_inv712;
  assign b_inv712 = ~b712;
  assign s712  = a712 ^ b712 ^ c712;
  assign sub712 = a712 ^ b_inv712 ^ c712;
  assign and712 = a712 & b712;
  assign or712  = a712 | b712;
  assign c713 = (a712 & b712) | (a712 & c712) | (b712 & c712);
  wire c_sub713;
  assign c_sub713 = (a712 & b_inv712) | (a712 & c712) | (b_inv712 & c712);
  wire s713, sub713, and713, or713;
  wire b_inv713;
  assign b_inv713 = ~b713;
  assign s713  = a713 ^ b713 ^ c713;
  assign sub713 = a713 ^ b_inv713 ^ c713;
  assign and713 = a713 & b713;
  assign or713  = a713 | b713;
  assign c714 = (a713 & b713) | (a713 & c713) | (b713 & c713);
  wire c_sub714;
  assign c_sub714 = (a713 & b_inv713) | (a713 & c713) | (b_inv713 & c713);
  wire s714, sub714, and714, or714;
  wire b_inv714;
  assign b_inv714 = ~b714;
  assign s714  = a714 ^ b714 ^ c714;
  assign sub714 = a714 ^ b_inv714 ^ c714;
  assign and714 = a714 & b714;
  assign or714  = a714 | b714;
  assign c715 = (a714 & b714) | (a714 & c714) | (b714 & c714);
  wire c_sub715;
  assign c_sub715 = (a714 & b_inv714) | (a714 & c714) | (b_inv714 & c714);
  wire s715, sub715, and715, or715;
  wire b_inv715;
  assign b_inv715 = ~b715;
  assign s715  = a715 ^ b715 ^ c715;
  assign sub715 = a715 ^ b_inv715 ^ c715;
  assign and715 = a715 & b715;
  assign or715  = a715 | b715;
  assign c716 = (a715 & b715) | (a715 & c715) | (b715 & c715);
  wire c_sub716;
  assign c_sub716 = (a715 & b_inv715) | (a715 & c715) | (b_inv715 & c715);
  wire s716, sub716, and716, or716;
  wire b_inv716;
  assign b_inv716 = ~b716;
  assign s716  = a716 ^ b716 ^ c716;
  assign sub716 = a716 ^ b_inv716 ^ c716;
  assign and716 = a716 & b716;
  assign or716  = a716 | b716;
  assign c717 = (a716 & b716) | (a716 & c716) | (b716 & c716);
  wire c_sub717;
  assign c_sub717 = (a716 & b_inv716) | (a716 & c716) | (b_inv716 & c716);
  wire s717, sub717, and717, or717;
  wire b_inv717;
  assign b_inv717 = ~b717;
  assign s717  = a717 ^ b717 ^ c717;
  assign sub717 = a717 ^ b_inv717 ^ c717;
  assign and717 = a717 & b717;
  assign or717  = a717 | b717;
  assign c718 = (a717 & b717) | (a717 & c717) | (b717 & c717);
  wire c_sub718;
  assign c_sub718 = (a717 & b_inv717) | (a717 & c717) | (b_inv717 & c717);
  wire s718, sub718, and718, or718;
  wire b_inv718;
  assign b_inv718 = ~b718;
  assign s718  = a718 ^ b718 ^ c718;
  assign sub718 = a718 ^ b_inv718 ^ c718;
  assign and718 = a718 & b718;
  assign or718  = a718 | b718;
  assign c719 = (a718 & b718) | (a718 & c718) | (b718 & c718);
  wire c_sub719;
  assign c_sub719 = (a718 & b_inv718) | (a718 & c718) | (b_inv718 & c718);
  wire s719, sub719, and719, or719;
  wire b_inv719;
  assign b_inv719 = ~b719;
  assign s719  = a719 ^ b719 ^ c719;
  assign sub719 = a719 ^ b_inv719 ^ c719;
  assign and719 = a719 & b719;
  assign or719  = a719 | b719;
  assign c720 = (a719 & b719) | (a719 & c719) | (b719 & c719);
  wire c_sub720;
  assign c_sub720 = (a719 & b_inv719) | (a719 & c719) | (b_inv719 & c719);
  wire s720, sub720, and720, or720;
  wire b_inv720;
  assign b_inv720 = ~b720;
  assign s720  = a720 ^ b720 ^ c720;
  assign sub720 = a720 ^ b_inv720 ^ c720;
  assign and720 = a720 & b720;
  assign or720  = a720 | b720;
  assign c721 = (a720 & b720) | (a720 & c720) | (b720 & c720);
  wire c_sub721;
  assign c_sub721 = (a720 & b_inv720) | (a720 & c720) | (b_inv720 & c720);
  wire s721, sub721, and721, or721;
  wire b_inv721;
  assign b_inv721 = ~b721;
  assign s721  = a721 ^ b721 ^ c721;
  assign sub721 = a721 ^ b_inv721 ^ c721;
  assign and721 = a721 & b721;
  assign or721  = a721 | b721;
  assign c722 = (a721 & b721) | (a721 & c721) | (b721 & c721);
  wire c_sub722;
  assign c_sub722 = (a721 & b_inv721) | (a721 & c721) | (b_inv721 & c721);
  wire s722, sub722, and722, or722;
  wire b_inv722;
  assign b_inv722 = ~b722;
  assign s722  = a722 ^ b722 ^ c722;
  assign sub722 = a722 ^ b_inv722 ^ c722;
  assign and722 = a722 & b722;
  assign or722  = a722 | b722;
  assign c723 = (a722 & b722) | (a722 & c722) | (b722 & c722);
  wire c_sub723;
  assign c_sub723 = (a722 & b_inv722) | (a722 & c722) | (b_inv722 & c722);
  wire s723, sub723, and723, or723;
  wire b_inv723;
  assign b_inv723 = ~b723;
  assign s723  = a723 ^ b723 ^ c723;
  assign sub723 = a723 ^ b_inv723 ^ c723;
  assign and723 = a723 & b723;
  assign or723  = a723 | b723;
  assign c724 = (a723 & b723) | (a723 & c723) | (b723 & c723);
  wire c_sub724;
  assign c_sub724 = (a723 & b_inv723) | (a723 & c723) | (b_inv723 & c723);
  wire s724, sub724, and724, or724;
  wire b_inv724;
  assign b_inv724 = ~b724;
  assign s724  = a724 ^ b724 ^ c724;
  assign sub724 = a724 ^ b_inv724 ^ c724;
  assign and724 = a724 & b724;
  assign or724  = a724 | b724;
  assign c725 = (a724 & b724) | (a724 & c724) | (b724 & c724);
  wire c_sub725;
  assign c_sub725 = (a724 & b_inv724) | (a724 & c724) | (b_inv724 & c724);
  wire s725, sub725, and725, or725;
  wire b_inv725;
  assign b_inv725 = ~b725;
  assign s725  = a725 ^ b725 ^ c725;
  assign sub725 = a725 ^ b_inv725 ^ c725;
  assign and725 = a725 & b725;
  assign or725  = a725 | b725;
  assign c726 = (a725 & b725) | (a725 & c725) | (b725 & c725);
  wire c_sub726;
  assign c_sub726 = (a725 & b_inv725) | (a725 & c725) | (b_inv725 & c725);
  wire s726, sub726, and726, or726;
  wire b_inv726;
  assign b_inv726 = ~b726;
  assign s726  = a726 ^ b726 ^ c726;
  assign sub726 = a726 ^ b_inv726 ^ c726;
  assign and726 = a726 & b726;
  assign or726  = a726 | b726;
  assign c727 = (a726 & b726) | (a726 & c726) | (b726 & c726);
  wire c_sub727;
  assign c_sub727 = (a726 & b_inv726) | (a726 & c726) | (b_inv726 & c726);
  wire s727, sub727, and727, or727;
  wire b_inv727;
  assign b_inv727 = ~b727;
  assign s727  = a727 ^ b727 ^ c727;
  assign sub727 = a727 ^ b_inv727 ^ c727;
  assign and727 = a727 & b727;
  assign or727  = a727 | b727;
  assign c728 = (a727 & b727) | (a727 & c727) | (b727 & c727);
  wire c_sub728;
  assign c_sub728 = (a727 & b_inv727) | (a727 & c727) | (b_inv727 & c727);
  wire s728, sub728, and728, or728;
  wire b_inv728;
  assign b_inv728 = ~b728;
  assign s728  = a728 ^ b728 ^ c728;
  assign sub728 = a728 ^ b_inv728 ^ c728;
  assign and728 = a728 & b728;
  assign or728  = a728 | b728;
  assign c729 = (a728 & b728) | (a728 & c728) | (b728 & c728);
  wire c_sub729;
  assign c_sub729 = (a728 & b_inv728) | (a728 & c728) | (b_inv728 & c728);
  wire s729, sub729, and729, or729;
  wire b_inv729;
  assign b_inv729 = ~b729;
  assign s729  = a729 ^ b729 ^ c729;
  assign sub729 = a729 ^ b_inv729 ^ c729;
  assign and729 = a729 & b729;
  assign or729  = a729 | b729;
  assign c730 = (a729 & b729) | (a729 & c729) | (b729 & c729);
  wire c_sub730;
  assign c_sub730 = (a729 & b_inv729) | (a729 & c729) | (b_inv729 & c729);
  wire s730, sub730, and730, or730;
  wire b_inv730;
  assign b_inv730 = ~b730;
  assign s730  = a730 ^ b730 ^ c730;
  assign sub730 = a730 ^ b_inv730 ^ c730;
  assign and730 = a730 & b730;
  assign or730  = a730 | b730;
  assign c731 = (a730 & b730) | (a730 & c730) | (b730 & c730);
  wire c_sub731;
  assign c_sub731 = (a730 & b_inv730) | (a730 & c730) | (b_inv730 & c730);
  wire s731, sub731, and731, or731;
  wire b_inv731;
  assign b_inv731 = ~b731;
  assign s731  = a731 ^ b731 ^ c731;
  assign sub731 = a731 ^ b_inv731 ^ c731;
  assign and731 = a731 & b731;
  assign or731  = a731 | b731;
  assign c732 = (a731 & b731) | (a731 & c731) | (b731 & c731);
  wire c_sub732;
  assign c_sub732 = (a731 & b_inv731) | (a731 & c731) | (b_inv731 & c731);
  wire s732, sub732, and732, or732;
  wire b_inv732;
  assign b_inv732 = ~b732;
  assign s732  = a732 ^ b732 ^ c732;
  assign sub732 = a732 ^ b_inv732 ^ c732;
  assign and732 = a732 & b732;
  assign or732  = a732 | b732;
  assign c733 = (a732 & b732) | (a732 & c732) | (b732 & c732);
  wire c_sub733;
  assign c_sub733 = (a732 & b_inv732) | (a732 & c732) | (b_inv732 & c732);
  wire s733, sub733, and733, or733;
  wire b_inv733;
  assign b_inv733 = ~b733;
  assign s733  = a733 ^ b733 ^ c733;
  assign sub733 = a733 ^ b_inv733 ^ c733;
  assign and733 = a733 & b733;
  assign or733  = a733 | b733;
  assign c734 = (a733 & b733) | (a733 & c733) | (b733 & c733);
  wire c_sub734;
  assign c_sub734 = (a733 & b_inv733) | (a733 & c733) | (b_inv733 & c733);
  wire s734, sub734, and734, or734;
  wire b_inv734;
  assign b_inv734 = ~b734;
  assign s734  = a734 ^ b734 ^ c734;
  assign sub734 = a734 ^ b_inv734 ^ c734;
  assign and734 = a734 & b734;
  assign or734  = a734 | b734;
  assign c735 = (a734 & b734) | (a734 & c734) | (b734 & c734);
  wire c_sub735;
  assign c_sub735 = (a734 & b_inv734) | (a734 & c734) | (b_inv734 & c734);
  wire s735, sub735, and735, or735;
  wire b_inv735;
  assign b_inv735 = ~b735;
  assign s735  = a735 ^ b735 ^ c735;
  assign sub735 = a735 ^ b_inv735 ^ c735;
  assign and735 = a735 & b735;
  assign or735  = a735 | b735;
  assign c736 = (a735 & b735) | (a735 & c735) | (b735 & c735);
  wire c_sub736;
  assign c_sub736 = (a735 & b_inv735) | (a735 & c735) | (b_inv735 & c735);
  wire s736, sub736, and736, or736;
  wire b_inv736;
  assign b_inv736 = ~b736;
  assign s736  = a736 ^ b736 ^ c736;
  assign sub736 = a736 ^ b_inv736 ^ c736;
  assign and736 = a736 & b736;
  assign or736  = a736 | b736;
  assign c737 = (a736 & b736) | (a736 & c736) | (b736 & c736);
  wire c_sub737;
  assign c_sub737 = (a736 & b_inv736) | (a736 & c736) | (b_inv736 & c736);
  wire s737, sub737, and737, or737;
  wire b_inv737;
  assign b_inv737 = ~b737;
  assign s737  = a737 ^ b737 ^ c737;
  assign sub737 = a737 ^ b_inv737 ^ c737;
  assign and737 = a737 & b737;
  assign or737  = a737 | b737;
  assign c738 = (a737 & b737) | (a737 & c737) | (b737 & c737);
  wire c_sub738;
  assign c_sub738 = (a737 & b_inv737) | (a737 & c737) | (b_inv737 & c737);
  wire s738, sub738, and738, or738;
  wire b_inv738;
  assign b_inv738 = ~b738;
  assign s738  = a738 ^ b738 ^ c738;
  assign sub738 = a738 ^ b_inv738 ^ c738;
  assign and738 = a738 & b738;
  assign or738  = a738 | b738;
  assign c739 = (a738 & b738) | (a738 & c738) | (b738 & c738);
  wire c_sub739;
  assign c_sub739 = (a738 & b_inv738) | (a738 & c738) | (b_inv738 & c738);
  wire s739, sub739, and739, or739;
  wire b_inv739;
  assign b_inv739 = ~b739;
  assign s739  = a739 ^ b739 ^ c739;
  assign sub739 = a739 ^ b_inv739 ^ c739;
  assign and739 = a739 & b739;
  assign or739  = a739 | b739;
  assign c740 = (a739 & b739) | (a739 & c739) | (b739 & c739);
  wire c_sub740;
  assign c_sub740 = (a739 & b_inv739) | (a739 & c739) | (b_inv739 & c739);
  wire s740, sub740, and740, or740;
  wire b_inv740;
  assign b_inv740 = ~b740;
  assign s740  = a740 ^ b740 ^ c740;
  assign sub740 = a740 ^ b_inv740 ^ c740;
  assign and740 = a740 & b740;
  assign or740  = a740 | b740;
  assign c741 = (a740 & b740) | (a740 & c740) | (b740 & c740);
  wire c_sub741;
  assign c_sub741 = (a740 & b_inv740) | (a740 & c740) | (b_inv740 & c740);
  wire s741, sub741, and741, or741;
  wire b_inv741;
  assign b_inv741 = ~b741;
  assign s741  = a741 ^ b741 ^ c741;
  assign sub741 = a741 ^ b_inv741 ^ c741;
  assign and741 = a741 & b741;
  assign or741  = a741 | b741;
  assign c742 = (a741 & b741) | (a741 & c741) | (b741 & c741);
  wire c_sub742;
  assign c_sub742 = (a741 & b_inv741) | (a741 & c741) | (b_inv741 & c741);
  wire s742, sub742, and742, or742;
  wire b_inv742;
  assign b_inv742 = ~b742;
  assign s742  = a742 ^ b742 ^ c742;
  assign sub742 = a742 ^ b_inv742 ^ c742;
  assign and742 = a742 & b742;
  assign or742  = a742 | b742;
  assign c743 = (a742 & b742) | (a742 & c742) | (b742 & c742);
  wire c_sub743;
  assign c_sub743 = (a742 & b_inv742) | (a742 & c742) | (b_inv742 & c742);
  wire s743, sub743, and743, or743;
  wire b_inv743;
  assign b_inv743 = ~b743;
  assign s743  = a743 ^ b743 ^ c743;
  assign sub743 = a743 ^ b_inv743 ^ c743;
  assign and743 = a743 & b743;
  assign or743  = a743 | b743;
  assign c744 = (a743 & b743) | (a743 & c743) | (b743 & c743);
  wire c_sub744;
  assign c_sub744 = (a743 & b_inv743) | (a743 & c743) | (b_inv743 & c743);
  wire s744, sub744, and744, or744;
  wire b_inv744;
  assign b_inv744 = ~b744;
  assign s744  = a744 ^ b744 ^ c744;
  assign sub744 = a744 ^ b_inv744 ^ c744;
  assign and744 = a744 & b744;
  assign or744  = a744 | b744;
  assign c745 = (a744 & b744) | (a744 & c744) | (b744 & c744);
  wire c_sub745;
  assign c_sub745 = (a744 & b_inv744) | (a744 & c744) | (b_inv744 & c744);
  wire s745, sub745, and745, or745;
  wire b_inv745;
  assign b_inv745 = ~b745;
  assign s745  = a745 ^ b745 ^ c745;
  assign sub745 = a745 ^ b_inv745 ^ c745;
  assign and745 = a745 & b745;
  assign or745  = a745 | b745;
  assign c746 = (a745 & b745) | (a745 & c745) | (b745 & c745);
  wire c_sub746;
  assign c_sub746 = (a745 & b_inv745) | (a745 & c745) | (b_inv745 & c745);
  wire s746, sub746, and746, or746;
  wire b_inv746;
  assign b_inv746 = ~b746;
  assign s746  = a746 ^ b746 ^ c746;
  assign sub746 = a746 ^ b_inv746 ^ c746;
  assign and746 = a746 & b746;
  assign or746  = a746 | b746;
  assign c747 = (a746 & b746) | (a746 & c746) | (b746 & c746);
  wire c_sub747;
  assign c_sub747 = (a746 & b_inv746) | (a746 & c746) | (b_inv746 & c746);
  wire s747, sub747, and747, or747;
  wire b_inv747;
  assign b_inv747 = ~b747;
  assign s747  = a747 ^ b747 ^ c747;
  assign sub747 = a747 ^ b_inv747 ^ c747;
  assign and747 = a747 & b747;
  assign or747  = a747 | b747;
  assign c748 = (a747 & b747) | (a747 & c747) | (b747 & c747);
  wire c_sub748;
  assign c_sub748 = (a747 & b_inv747) | (a747 & c747) | (b_inv747 & c747);
  wire s748, sub748, and748, or748;
  wire b_inv748;
  assign b_inv748 = ~b748;
  assign s748  = a748 ^ b748 ^ c748;
  assign sub748 = a748 ^ b_inv748 ^ c748;
  assign and748 = a748 & b748;
  assign or748  = a748 | b748;
  assign c749 = (a748 & b748) | (a748 & c748) | (b748 & c748);
  wire c_sub749;
  assign c_sub749 = (a748 & b_inv748) | (a748 & c748) | (b_inv748 & c748);
  wire s749, sub749, and749, or749;
  wire b_inv749;
  assign b_inv749 = ~b749;
  assign s749  = a749 ^ b749 ^ c749;
  assign sub749 = a749 ^ b_inv749 ^ c749;
  assign and749 = a749 & b749;
  assign or749  = a749 | b749;
  assign c750 = (a749 & b749) | (a749 & c749) | (b749 & c749);
  wire c_sub750;
  assign c_sub750 = (a749 & b_inv749) | (a749 & c749) | (b_inv749 & c749);
  wire s750, sub750, and750, or750;
  wire b_inv750;
  assign b_inv750 = ~b750;
  assign s750  = a750 ^ b750 ^ c750;
  assign sub750 = a750 ^ b_inv750 ^ c750;
  assign and750 = a750 & b750;
  assign or750  = a750 | b750;
  assign c751 = (a750 & b750) | (a750 & c750) | (b750 & c750);
  wire c_sub751;
  assign c_sub751 = (a750 & b_inv750) | (a750 & c750) | (b_inv750 & c750);
  wire s751, sub751, and751, or751;
  wire b_inv751;
  assign b_inv751 = ~b751;
  assign s751  = a751 ^ b751 ^ c751;
  assign sub751 = a751 ^ b_inv751 ^ c751;
  assign and751 = a751 & b751;
  assign or751  = a751 | b751;
  assign c752 = (a751 & b751) | (a751 & c751) | (b751 & c751);
  wire c_sub752;
  assign c_sub752 = (a751 & b_inv751) | (a751 & c751) | (b_inv751 & c751);
  wire s752, sub752, and752, or752;
  wire b_inv752;
  assign b_inv752 = ~b752;
  assign s752  = a752 ^ b752 ^ c752;
  assign sub752 = a752 ^ b_inv752 ^ c752;
  assign and752 = a752 & b752;
  assign or752  = a752 | b752;
  assign c753 = (a752 & b752) | (a752 & c752) | (b752 & c752);
  wire c_sub753;
  assign c_sub753 = (a752 & b_inv752) | (a752 & c752) | (b_inv752 & c752);
  wire s753, sub753, and753, or753;
  wire b_inv753;
  assign b_inv753 = ~b753;
  assign s753  = a753 ^ b753 ^ c753;
  assign sub753 = a753 ^ b_inv753 ^ c753;
  assign and753 = a753 & b753;
  assign or753  = a753 | b753;
  assign c754 = (a753 & b753) | (a753 & c753) | (b753 & c753);
  wire c_sub754;
  assign c_sub754 = (a753 & b_inv753) | (a753 & c753) | (b_inv753 & c753);
  wire s754, sub754, and754, or754;
  wire b_inv754;
  assign b_inv754 = ~b754;
  assign s754  = a754 ^ b754 ^ c754;
  assign sub754 = a754 ^ b_inv754 ^ c754;
  assign and754 = a754 & b754;
  assign or754  = a754 | b754;
  assign c755 = (a754 & b754) | (a754 & c754) | (b754 & c754);
  wire c_sub755;
  assign c_sub755 = (a754 & b_inv754) | (a754 & c754) | (b_inv754 & c754);
  wire s755, sub755, and755, or755;
  wire b_inv755;
  assign b_inv755 = ~b755;
  assign s755  = a755 ^ b755 ^ c755;
  assign sub755 = a755 ^ b_inv755 ^ c755;
  assign and755 = a755 & b755;
  assign or755  = a755 | b755;
  assign c756 = (a755 & b755) | (a755 & c755) | (b755 & c755);
  wire c_sub756;
  assign c_sub756 = (a755 & b_inv755) | (a755 & c755) | (b_inv755 & c755);
  wire s756, sub756, and756, or756;
  wire b_inv756;
  assign b_inv756 = ~b756;
  assign s756  = a756 ^ b756 ^ c756;
  assign sub756 = a756 ^ b_inv756 ^ c756;
  assign and756 = a756 & b756;
  assign or756  = a756 | b756;
  assign c757 = (a756 & b756) | (a756 & c756) | (b756 & c756);
  wire c_sub757;
  assign c_sub757 = (a756 & b_inv756) | (a756 & c756) | (b_inv756 & c756);
  wire s757, sub757, and757, or757;
  wire b_inv757;
  assign b_inv757 = ~b757;
  assign s757  = a757 ^ b757 ^ c757;
  assign sub757 = a757 ^ b_inv757 ^ c757;
  assign and757 = a757 & b757;
  assign or757  = a757 | b757;
  assign c758 = (a757 & b757) | (a757 & c757) | (b757 & c757);
  wire c_sub758;
  assign c_sub758 = (a757 & b_inv757) | (a757 & c757) | (b_inv757 & c757);
  wire s758, sub758, and758, or758;
  wire b_inv758;
  assign b_inv758 = ~b758;
  assign s758  = a758 ^ b758 ^ c758;
  assign sub758 = a758 ^ b_inv758 ^ c758;
  assign and758 = a758 & b758;
  assign or758  = a758 | b758;
  assign c759 = (a758 & b758) | (a758 & c758) | (b758 & c758);
  wire c_sub759;
  assign c_sub759 = (a758 & b_inv758) | (a758 & c758) | (b_inv758 & c758);
  wire s759, sub759, and759, or759;
  wire b_inv759;
  assign b_inv759 = ~b759;
  assign s759  = a759 ^ b759 ^ c759;
  assign sub759 = a759 ^ b_inv759 ^ c759;
  assign and759 = a759 & b759;
  assign or759  = a759 | b759;
  assign c760 = (a759 & b759) | (a759 & c759) | (b759 & c759);
  wire c_sub760;
  assign c_sub760 = (a759 & b_inv759) | (a759 & c759) | (b_inv759 & c759);
  wire s760, sub760, and760, or760;
  wire b_inv760;
  assign b_inv760 = ~b760;
  assign s760  = a760 ^ b760 ^ c760;
  assign sub760 = a760 ^ b_inv760 ^ c760;
  assign and760 = a760 & b760;
  assign or760  = a760 | b760;
  assign c761 = (a760 & b760) | (a760 & c760) | (b760 & c760);
  wire c_sub761;
  assign c_sub761 = (a760 & b_inv760) | (a760 & c760) | (b_inv760 & c760);
  wire s761, sub761, and761, or761;
  wire b_inv761;
  assign b_inv761 = ~b761;
  assign s761  = a761 ^ b761 ^ c761;
  assign sub761 = a761 ^ b_inv761 ^ c761;
  assign and761 = a761 & b761;
  assign or761  = a761 | b761;
  assign c762 = (a761 & b761) | (a761 & c761) | (b761 & c761);
  wire c_sub762;
  assign c_sub762 = (a761 & b_inv761) | (a761 & c761) | (b_inv761 & c761);
  wire s762, sub762, and762, or762;
  wire b_inv762;
  assign b_inv762 = ~b762;
  assign s762  = a762 ^ b762 ^ c762;
  assign sub762 = a762 ^ b_inv762 ^ c762;
  assign and762 = a762 & b762;
  assign or762  = a762 | b762;
  assign c763 = (a762 & b762) | (a762 & c762) | (b762 & c762);
  wire c_sub763;
  assign c_sub763 = (a762 & b_inv762) | (a762 & c762) | (b_inv762 & c762);
  wire s763, sub763, and763, or763;
  wire b_inv763;
  assign b_inv763 = ~b763;
  assign s763  = a763 ^ b763 ^ c763;
  assign sub763 = a763 ^ b_inv763 ^ c763;
  assign and763 = a763 & b763;
  assign or763  = a763 | b763;
  assign c764 = (a763 & b763) | (a763 & c763) | (b763 & c763);
  wire c_sub764;
  assign c_sub764 = (a763 & b_inv763) | (a763 & c763) | (b_inv763 & c763);
  wire s764, sub764, and764, or764;
  wire b_inv764;
  assign b_inv764 = ~b764;
  assign s764  = a764 ^ b764 ^ c764;
  assign sub764 = a764 ^ b_inv764 ^ c764;
  assign and764 = a764 & b764;
  assign or764  = a764 | b764;
  assign c765 = (a764 & b764) | (a764 & c764) | (b764 & c764);
  wire c_sub765;
  assign c_sub765 = (a764 & b_inv764) | (a764 & c764) | (b_inv764 & c764);
  wire s765, sub765, and765, or765;
  wire b_inv765;
  assign b_inv765 = ~b765;
  assign s765  = a765 ^ b765 ^ c765;
  assign sub765 = a765 ^ b_inv765 ^ c765;
  assign and765 = a765 & b765;
  assign or765  = a765 | b765;
  assign c766 = (a765 & b765) | (a765 & c765) | (b765 & c765);
  wire c_sub766;
  assign c_sub766 = (a765 & b_inv765) | (a765 & c765) | (b_inv765 & c765);
  wire s766, sub766, and766, or766;
  wire b_inv766;
  assign b_inv766 = ~b766;
  assign s766  = a766 ^ b766 ^ c766;
  assign sub766 = a766 ^ b_inv766 ^ c766;
  assign and766 = a766 & b766;
  assign or766  = a766 | b766;
  assign c767 = (a766 & b766) | (a766 & c766) | (b766 & c766);
  wire c_sub767;
  assign c_sub767 = (a766 & b_inv766) | (a766 & c766) | (b_inv766 & c766);
  wire s767, sub767, and767, or767;
  wire b_inv767;
  assign b_inv767 = ~b767;
  assign s767  = a767 ^ b767 ^ c767;
  assign sub767 = a767 ^ b_inv767 ^ c767;
  assign and767 = a767 & b767;
  assign or767  = a767 | b767;
  assign c768 = (a767 & b767) | (a767 & c767) | (b767 & c767);
  wire c_sub768;
  assign c_sub768 = (a767 & b_inv767) | (a767 & c767) | (b_inv767 & c767);
  wire s768, sub768, and768, or768;
  wire b_inv768;
  assign b_inv768 = ~b768;
  assign s768  = a768 ^ b768 ^ c768;
  assign sub768 = a768 ^ b_inv768 ^ c768;
  assign and768 = a768 & b768;
  assign or768  = a768 | b768;
  assign c769 = (a768 & b768) | (a768 & c768) | (b768 & c768);
  wire c_sub769;
  assign c_sub769 = (a768 & b_inv768) | (a768 & c768) | (b_inv768 & c768);
  wire s769, sub769, and769, or769;
  wire b_inv769;
  assign b_inv769 = ~b769;
  assign s769  = a769 ^ b769 ^ c769;
  assign sub769 = a769 ^ b_inv769 ^ c769;
  assign and769 = a769 & b769;
  assign or769  = a769 | b769;
  assign c770 = (a769 & b769) | (a769 & c769) | (b769 & c769);
  wire c_sub770;
  assign c_sub770 = (a769 & b_inv769) | (a769 & c769) | (b_inv769 & c769);
  wire s770, sub770, and770, or770;
  wire b_inv770;
  assign b_inv770 = ~b770;
  assign s770  = a770 ^ b770 ^ c770;
  assign sub770 = a770 ^ b_inv770 ^ c770;
  assign and770 = a770 & b770;
  assign or770  = a770 | b770;
  assign c771 = (a770 & b770) | (a770 & c770) | (b770 & c770);
  wire c_sub771;
  assign c_sub771 = (a770 & b_inv770) | (a770 & c770) | (b_inv770 & c770);
  wire s771, sub771, and771, or771;
  wire b_inv771;
  assign b_inv771 = ~b771;
  assign s771  = a771 ^ b771 ^ c771;
  assign sub771 = a771 ^ b_inv771 ^ c771;
  assign and771 = a771 & b771;
  assign or771  = a771 | b771;
  assign c772 = (a771 & b771) | (a771 & c771) | (b771 & c771);
  wire c_sub772;
  assign c_sub772 = (a771 & b_inv771) | (a771 & c771) | (b_inv771 & c771);
  wire s772, sub772, and772, or772;
  wire b_inv772;
  assign b_inv772 = ~b772;
  assign s772  = a772 ^ b772 ^ c772;
  assign sub772 = a772 ^ b_inv772 ^ c772;
  assign and772 = a772 & b772;
  assign or772  = a772 | b772;
  assign c773 = (a772 & b772) | (a772 & c772) | (b772 & c772);
  wire c_sub773;
  assign c_sub773 = (a772 & b_inv772) | (a772 & c772) | (b_inv772 & c772);
  wire s773, sub773, and773, or773;
  wire b_inv773;
  assign b_inv773 = ~b773;
  assign s773  = a773 ^ b773 ^ c773;
  assign sub773 = a773 ^ b_inv773 ^ c773;
  assign and773 = a773 & b773;
  assign or773  = a773 | b773;
  assign c774 = (a773 & b773) | (a773 & c773) | (b773 & c773);
  wire c_sub774;
  assign c_sub774 = (a773 & b_inv773) | (a773 & c773) | (b_inv773 & c773);
  wire s774, sub774, and774, or774;
  wire b_inv774;
  assign b_inv774 = ~b774;
  assign s774  = a774 ^ b774 ^ c774;
  assign sub774 = a774 ^ b_inv774 ^ c774;
  assign and774 = a774 & b774;
  assign or774  = a774 | b774;
  assign c775 = (a774 & b774) | (a774 & c774) | (b774 & c774);
  wire c_sub775;
  assign c_sub775 = (a774 & b_inv774) | (a774 & c774) | (b_inv774 & c774);
  wire s775, sub775, and775, or775;
  wire b_inv775;
  assign b_inv775 = ~b775;
  assign s775  = a775 ^ b775 ^ c775;
  assign sub775 = a775 ^ b_inv775 ^ c775;
  assign and775 = a775 & b775;
  assign or775  = a775 | b775;
  assign c776 = (a775 & b775) | (a775 & c775) | (b775 & c775);
  wire c_sub776;
  assign c_sub776 = (a775 & b_inv775) | (a775 & c775) | (b_inv775 & c775);
  wire s776, sub776, and776, or776;
  wire b_inv776;
  assign b_inv776 = ~b776;
  assign s776  = a776 ^ b776 ^ c776;
  assign sub776 = a776 ^ b_inv776 ^ c776;
  assign and776 = a776 & b776;
  assign or776  = a776 | b776;
  assign c777 = (a776 & b776) | (a776 & c776) | (b776 & c776);
  wire c_sub777;
  assign c_sub777 = (a776 & b_inv776) | (a776 & c776) | (b_inv776 & c776);
  wire s777, sub777, and777, or777;
  wire b_inv777;
  assign b_inv777 = ~b777;
  assign s777  = a777 ^ b777 ^ c777;
  assign sub777 = a777 ^ b_inv777 ^ c777;
  assign and777 = a777 & b777;
  assign or777  = a777 | b777;
  assign c778 = (a777 & b777) | (a777 & c777) | (b777 & c777);
  wire c_sub778;
  assign c_sub778 = (a777 & b_inv777) | (a777 & c777) | (b_inv777 & c777);
  wire s778, sub778, and778, or778;
  wire b_inv778;
  assign b_inv778 = ~b778;
  assign s778  = a778 ^ b778 ^ c778;
  assign sub778 = a778 ^ b_inv778 ^ c778;
  assign and778 = a778 & b778;
  assign or778  = a778 | b778;
  assign c779 = (a778 & b778) | (a778 & c778) | (b778 & c778);
  wire c_sub779;
  assign c_sub779 = (a778 & b_inv778) | (a778 & c778) | (b_inv778 & c778);
  wire s779, sub779, and779, or779;
  wire b_inv779;
  assign b_inv779 = ~b779;
  assign s779  = a779 ^ b779 ^ c779;
  assign sub779 = a779 ^ b_inv779 ^ c779;
  assign and779 = a779 & b779;
  assign or779  = a779 | b779;
  assign c780 = (a779 & b779) | (a779 & c779) | (b779 & c779);
  wire c_sub780;
  assign c_sub780 = (a779 & b_inv779) | (a779 & c779) | (b_inv779 & c779);
  wire s780, sub780, and780, or780;
  wire b_inv780;
  assign b_inv780 = ~b780;
  assign s780  = a780 ^ b780 ^ c780;
  assign sub780 = a780 ^ b_inv780 ^ c780;
  assign and780 = a780 & b780;
  assign or780  = a780 | b780;
  assign c781 = (a780 & b780) | (a780 & c780) | (b780 & c780);
  wire c_sub781;
  assign c_sub781 = (a780 & b_inv780) | (a780 & c780) | (b_inv780 & c780);
  wire s781, sub781, and781, or781;
  wire b_inv781;
  assign b_inv781 = ~b781;
  assign s781  = a781 ^ b781 ^ c781;
  assign sub781 = a781 ^ b_inv781 ^ c781;
  assign and781 = a781 & b781;
  assign or781  = a781 | b781;
  assign c782 = (a781 & b781) | (a781 & c781) | (b781 & c781);
  wire c_sub782;
  assign c_sub782 = (a781 & b_inv781) | (a781 & c781) | (b_inv781 & c781);
  wire s782, sub782, and782, or782;
  wire b_inv782;
  assign b_inv782 = ~b782;
  assign s782  = a782 ^ b782 ^ c782;
  assign sub782 = a782 ^ b_inv782 ^ c782;
  assign and782 = a782 & b782;
  assign or782  = a782 | b782;
  assign c783 = (a782 & b782) | (a782 & c782) | (b782 & c782);
  wire c_sub783;
  assign c_sub783 = (a782 & b_inv782) | (a782 & c782) | (b_inv782 & c782);
  wire s783, sub783, and783, or783;
  wire b_inv783;
  assign b_inv783 = ~b783;
  assign s783  = a783 ^ b783 ^ c783;
  assign sub783 = a783 ^ b_inv783 ^ c783;
  assign and783 = a783 & b783;
  assign or783  = a783 | b783;
  assign c784 = (a783 & b783) | (a783 & c783) | (b783 & c783);
  wire c_sub784;
  assign c_sub784 = (a783 & b_inv783) | (a783 & c783) | (b_inv783 & c783);
  wire s784, sub784, and784, or784;
  wire b_inv784;
  assign b_inv784 = ~b784;
  assign s784  = a784 ^ b784 ^ c784;
  assign sub784 = a784 ^ b_inv784 ^ c784;
  assign and784 = a784 & b784;
  assign or784  = a784 | b784;
  assign c785 = (a784 & b784) | (a784 & c784) | (b784 & c784);
  wire c_sub785;
  assign c_sub785 = (a784 & b_inv784) | (a784 & c784) | (b_inv784 & c784);
  wire s785, sub785, and785, or785;
  wire b_inv785;
  assign b_inv785 = ~b785;
  assign s785  = a785 ^ b785 ^ c785;
  assign sub785 = a785 ^ b_inv785 ^ c785;
  assign and785 = a785 & b785;
  assign or785  = a785 | b785;
  assign c786 = (a785 & b785) | (a785 & c785) | (b785 & c785);
  wire c_sub786;
  assign c_sub786 = (a785 & b_inv785) | (a785 & c785) | (b_inv785 & c785);
  wire s786, sub786, and786, or786;
  wire b_inv786;
  assign b_inv786 = ~b786;
  assign s786  = a786 ^ b786 ^ c786;
  assign sub786 = a786 ^ b_inv786 ^ c786;
  assign and786 = a786 & b786;
  assign or786  = a786 | b786;
  assign c787 = (a786 & b786) | (a786 & c786) | (b786 & c786);
  wire c_sub787;
  assign c_sub787 = (a786 & b_inv786) | (a786 & c786) | (b_inv786 & c786);
  wire s787, sub787, and787, or787;
  wire b_inv787;
  assign b_inv787 = ~b787;
  assign s787  = a787 ^ b787 ^ c787;
  assign sub787 = a787 ^ b_inv787 ^ c787;
  assign and787 = a787 & b787;
  assign or787  = a787 | b787;
  assign c788 = (a787 & b787) | (a787 & c787) | (b787 & c787);
  wire c_sub788;
  assign c_sub788 = (a787 & b_inv787) | (a787 & c787) | (b_inv787 & c787);
  wire s788, sub788, and788, or788;
  wire b_inv788;
  assign b_inv788 = ~b788;
  assign s788  = a788 ^ b788 ^ c788;
  assign sub788 = a788 ^ b_inv788 ^ c788;
  assign and788 = a788 & b788;
  assign or788  = a788 | b788;
  assign c789 = (a788 & b788) | (a788 & c788) | (b788 & c788);
  wire c_sub789;
  assign c_sub789 = (a788 & b_inv788) | (a788 & c788) | (b_inv788 & c788);
  wire s789, sub789, and789, or789;
  wire b_inv789;
  assign b_inv789 = ~b789;
  assign s789  = a789 ^ b789 ^ c789;
  assign sub789 = a789 ^ b_inv789 ^ c789;
  assign and789 = a789 & b789;
  assign or789  = a789 | b789;
  assign c790 = (a789 & b789) | (a789 & c789) | (b789 & c789);
  wire c_sub790;
  assign c_sub790 = (a789 & b_inv789) | (a789 & c789) | (b_inv789 & c789);
  wire s790, sub790, and790, or790;
  wire b_inv790;
  assign b_inv790 = ~b790;
  assign s790  = a790 ^ b790 ^ c790;
  assign sub790 = a790 ^ b_inv790 ^ c790;
  assign and790 = a790 & b790;
  assign or790  = a790 | b790;
  assign c791 = (a790 & b790) | (a790 & c790) | (b790 & c790);
  wire c_sub791;
  assign c_sub791 = (a790 & b_inv790) | (a790 & c790) | (b_inv790 & c790);
  wire s791, sub791, and791, or791;
  wire b_inv791;
  assign b_inv791 = ~b791;
  assign s791  = a791 ^ b791 ^ c791;
  assign sub791 = a791 ^ b_inv791 ^ c791;
  assign and791 = a791 & b791;
  assign or791  = a791 | b791;
  assign c792 = (a791 & b791) | (a791 & c791) | (b791 & c791);
  wire c_sub792;
  assign c_sub792 = (a791 & b_inv791) | (a791 & c791) | (b_inv791 & c791);
  wire s792, sub792, and792, or792;
  wire b_inv792;
  assign b_inv792 = ~b792;
  assign s792  = a792 ^ b792 ^ c792;
  assign sub792 = a792 ^ b_inv792 ^ c792;
  assign and792 = a792 & b792;
  assign or792  = a792 | b792;
  assign c793 = (a792 & b792) | (a792 & c792) | (b792 & c792);
  wire c_sub793;
  assign c_sub793 = (a792 & b_inv792) | (a792 & c792) | (b_inv792 & c792);
  wire s793, sub793, and793, or793;
  wire b_inv793;
  assign b_inv793 = ~b793;
  assign s793  = a793 ^ b793 ^ c793;
  assign sub793 = a793 ^ b_inv793 ^ c793;
  assign and793 = a793 & b793;
  assign or793  = a793 | b793;
  assign c794 = (a793 & b793) | (a793 & c793) | (b793 & c793);
  wire c_sub794;
  assign c_sub794 = (a793 & b_inv793) | (a793 & c793) | (b_inv793 & c793);
  wire s794, sub794, and794, or794;
  wire b_inv794;
  assign b_inv794 = ~b794;
  assign s794  = a794 ^ b794 ^ c794;
  assign sub794 = a794 ^ b_inv794 ^ c794;
  assign and794 = a794 & b794;
  assign or794  = a794 | b794;
  assign c795 = (a794 & b794) | (a794 & c794) | (b794 & c794);
  wire c_sub795;
  assign c_sub795 = (a794 & b_inv794) | (a794 & c794) | (b_inv794 & c794);
  wire s795, sub795, and795, or795;
  wire b_inv795;
  assign b_inv795 = ~b795;
  assign s795  = a795 ^ b795 ^ c795;
  assign sub795 = a795 ^ b_inv795 ^ c795;
  assign and795 = a795 & b795;
  assign or795  = a795 | b795;
  assign c796 = (a795 & b795) | (a795 & c795) | (b795 & c795);
  wire c_sub796;
  assign c_sub796 = (a795 & b_inv795) | (a795 & c795) | (b_inv795 & c795);
  wire s796, sub796, and796, or796;
  wire b_inv796;
  assign b_inv796 = ~b796;
  assign s796  = a796 ^ b796 ^ c796;
  assign sub796 = a796 ^ b_inv796 ^ c796;
  assign and796 = a796 & b796;
  assign or796  = a796 | b796;
  assign c797 = (a796 & b796) | (a796 & c796) | (b796 & c796);
  wire c_sub797;
  assign c_sub797 = (a796 & b_inv796) | (a796 & c796) | (b_inv796 & c796);
  wire s797, sub797, and797, or797;
  wire b_inv797;
  assign b_inv797 = ~b797;
  assign s797  = a797 ^ b797 ^ c797;
  assign sub797 = a797 ^ b_inv797 ^ c797;
  assign and797 = a797 & b797;
  assign or797  = a797 | b797;
  assign c798 = (a797 & b797) | (a797 & c797) | (b797 & c797);
  wire c_sub798;
  assign c_sub798 = (a797 & b_inv797) | (a797 & c797) | (b_inv797 & c797);
  wire s798, sub798, and798, or798;
  wire b_inv798;
  assign b_inv798 = ~b798;
  assign s798  = a798 ^ b798 ^ c798;
  assign sub798 = a798 ^ b_inv798 ^ c798;
  assign and798 = a798 & b798;
  assign or798  = a798 | b798;
  assign c799 = (a798 & b798) | (a798 & c798) | (b798 & c798);
  wire c_sub799;
  assign c_sub799 = (a798 & b_inv798) | (a798 & c798) | (b_inv798 & c798);
  wire s799, sub799, and799, or799;
  wire b_inv799;
  assign b_inv799 = ~b799;
  assign s799  = a799 ^ b799 ^ c799;
  assign sub799 = a799 ^ b_inv799 ^ c799;
  assign and799 = a799 & b799;
  assign or799  = a799 | b799;
  assign c800 = (a799 & b799) | (a799 & c799) | (b799 & c799);
  wire c_sub800;
  assign c_sub800 = (a799 & b_inv799) | (a799 & c799) | (b_inv799 & c799);
  wire s800, sub800, and800, or800;
  wire b_inv800;
  assign b_inv800 = ~b800;
  assign s800  = a800 ^ b800 ^ c800;
  assign sub800 = a800 ^ b_inv800 ^ c800;
  assign and800 = a800 & b800;
  assign or800  = a800 | b800;
  assign c801 = (a800 & b800) | (a800 & c800) | (b800 & c800);
  wire c_sub801;
  assign c_sub801 = (a800 & b_inv800) | (a800 & c800) | (b_inv800 & c800);
  wire s801, sub801, and801, or801;
  wire b_inv801;
  assign b_inv801 = ~b801;
  assign s801  = a801 ^ b801 ^ c801;
  assign sub801 = a801 ^ b_inv801 ^ c801;
  assign and801 = a801 & b801;
  assign or801  = a801 | b801;
  assign c802 = (a801 & b801) | (a801 & c801) | (b801 & c801);
  wire c_sub802;
  assign c_sub802 = (a801 & b_inv801) | (a801 & c801) | (b_inv801 & c801);
  wire s802, sub802, and802, or802;
  wire b_inv802;
  assign b_inv802 = ~b802;
  assign s802  = a802 ^ b802 ^ c802;
  assign sub802 = a802 ^ b_inv802 ^ c802;
  assign and802 = a802 & b802;
  assign or802  = a802 | b802;
  assign c803 = (a802 & b802) | (a802 & c802) | (b802 & c802);
  wire c_sub803;
  assign c_sub803 = (a802 & b_inv802) | (a802 & c802) | (b_inv802 & c802);
  wire s803, sub803, and803, or803;
  wire b_inv803;
  assign b_inv803 = ~b803;
  assign s803  = a803 ^ b803 ^ c803;
  assign sub803 = a803 ^ b_inv803 ^ c803;
  assign and803 = a803 & b803;
  assign or803  = a803 | b803;
  assign c804 = (a803 & b803) | (a803 & c803) | (b803 & c803);
  wire c_sub804;
  assign c_sub804 = (a803 & b_inv803) | (a803 & c803) | (b_inv803 & c803);
  wire s804, sub804, and804, or804;
  wire b_inv804;
  assign b_inv804 = ~b804;
  assign s804  = a804 ^ b804 ^ c804;
  assign sub804 = a804 ^ b_inv804 ^ c804;
  assign and804 = a804 & b804;
  assign or804  = a804 | b804;
  assign c805 = (a804 & b804) | (a804 & c804) | (b804 & c804);
  wire c_sub805;
  assign c_sub805 = (a804 & b_inv804) | (a804 & c804) | (b_inv804 & c804);
  wire s805, sub805, and805, or805;
  wire b_inv805;
  assign b_inv805 = ~b805;
  assign s805  = a805 ^ b805 ^ c805;
  assign sub805 = a805 ^ b_inv805 ^ c805;
  assign and805 = a805 & b805;
  assign or805  = a805 | b805;
  assign c806 = (a805 & b805) | (a805 & c805) | (b805 & c805);
  wire c_sub806;
  assign c_sub806 = (a805 & b_inv805) | (a805 & c805) | (b_inv805 & c805);
  wire s806, sub806, and806, or806;
  wire b_inv806;
  assign b_inv806 = ~b806;
  assign s806  = a806 ^ b806 ^ c806;
  assign sub806 = a806 ^ b_inv806 ^ c806;
  assign and806 = a806 & b806;
  assign or806  = a806 | b806;
  assign c807 = (a806 & b806) | (a806 & c806) | (b806 & c806);
  wire c_sub807;
  assign c_sub807 = (a806 & b_inv806) | (a806 & c806) | (b_inv806 & c806);
  wire s807, sub807, and807, or807;
  wire b_inv807;
  assign b_inv807 = ~b807;
  assign s807  = a807 ^ b807 ^ c807;
  assign sub807 = a807 ^ b_inv807 ^ c807;
  assign and807 = a807 & b807;
  assign or807  = a807 | b807;
  assign c808 = (a807 & b807) | (a807 & c807) | (b807 & c807);
  wire c_sub808;
  assign c_sub808 = (a807 & b_inv807) | (a807 & c807) | (b_inv807 & c807);
  wire s808, sub808, and808, or808;
  wire b_inv808;
  assign b_inv808 = ~b808;
  assign s808  = a808 ^ b808 ^ c808;
  assign sub808 = a808 ^ b_inv808 ^ c808;
  assign and808 = a808 & b808;
  assign or808  = a808 | b808;
  assign c809 = (a808 & b808) | (a808 & c808) | (b808 & c808);
  wire c_sub809;
  assign c_sub809 = (a808 & b_inv808) | (a808 & c808) | (b_inv808 & c808);
  wire s809, sub809, and809, or809;
  wire b_inv809;
  assign b_inv809 = ~b809;
  assign s809  = a809 ^ b809 ^ c809;
  assign sub809 = a809 ^ b_inv809 ^ c809;
  assign and809 = a809 & b809;
  assign or809  = a809 | b809;
  assign c810 = (a809 & b809) | (a809 & c809) | (b809 & c809);
  wire c_sub810;
  assign c_sub810 = (a809 & b_inv809) | (a809 & c809) | (b_inv809 & c809);
  wire s810, sub810, and810, or810;
  wire b_inv810;
  assign b_inv810 = ~b810;
  assign s810  = a810 ^ b810 ^ c810;
  assign sub810 = a810 ^ b_inv810 ^ c810;
  assign and810 = a810 & b810;
  assign or810  = a810 | b810;
  assign c811 = (a810 & b810) | (a810 & c810) | (b810 & c810);
  wire c_sub811;
  assign c_sub811 = (a810 & b_inv810) | (a810 & c810) | (b_inv810 & c810);
  wire s811, sub811, and811, or811;
  wire b_inv811;
  assign b_inv811 = ~b811;
  assign s811  = a811 ^ b811 ^ c811;
  assign sub811 = a811 ^ b_inv811 ^ c811;
  assign and811 = a811 & b811;
  assign or811  = a811 | b811;
  assign c812 = (a811 & b811) | (a811 & c811) | (b811 & c811);
  wire c_sub812;
  assign c_sub812 = (a811 & b_inv811) | (a811 & c811) | (b_inv811 & c811);
  wire s812, sub812, and812, or812;
  wire b_inv812;
  assign b_inv812 = ~b812;
  assign s812  = a812 ^ b812 ^ c812;
  assign sub812 = a812 ^ b_inv812 ^ c812;
  assign and812 = a812 & b812;
  assign or812  = a812 | b812;
  assign c813 = (a812 & b812) | (a812 & c812) | (b812 & c812);
  wire c_sub813;
  assign c_sub813 = (a812 & b_inv812) | (a812 & c812) | (b_inv812 & c812);
  wire s813, sub813, and813, or813;
  wire b_inv813;
  assign b_inv813 = ~b813;
  assign s813  = a813 ^ b813 ^ c813;
  assign sub813 = a813 ^ b_inv813 ^ c813;
  assign and813 = a813 & b813;
  assign or813  = a813 | b813;
  assign c814 = (a813 & b813) | (a813 & c813) | (b813 & c813);
  wire c_sub814;
  assign c_sub814 = (a813 & b_inv813) | (a813 & c813) | (b_inv813 & c813);
  wire s814, sub814, and814, or814;
  wire b_inv814;
  assign b_inv814 = ~b814;
  assign s814  = a814 ^ b814 ^ c814;
  assign sub814 = a814 ^ b_inv814 ^ c814;
  assign and814 = a814 & b814;
  assign or814  = a814 | b814;
  assign c815 = (a814 & b814) | (a814 & c814) | (b814 & c814);
  wire c_sub815;
  assign c_sub815 = (a814 & b_inv814) | (a814 & c814) | (b_inv814 & c814);
  wire s815, sub815, and815, or815;
  wire b_inv815;
  assign b_inv815 = ~b815;
  assign s815  = a815 ^ b815 ^ c815;
  assign sub815 = a815 ^ b_inv815 ^ c815;
  assign and815 = a815 & b815;
  assign or815  = a815 | b815;
  assign c816 = (a815 & b815) | (a815 & c815) | (b815 & c815);
  wire c_sub816;
  assign c_sub816 = (a815 & b_inv815) | (a815 & c815) | (b_inv815 & c815);
  wire s816, sub816, and816, or816;
  wire b_inv816;
  assign b_inv816 = ~b816;
  assign s816  = a816 ^ b816 ^ c816;
  assign sub816 = a816 ^ b_inv816 ^ c816;
  assign and816 = a816 & b816;
  assign or816  = a816 | b816;
  assign c817 = (a816 & b816) | (a816 & c816) | (b816 & c816);
  wire c_sub817;
  assign c_sub817 = (a816 & b_inv816) | (a816 & c816) | (b_inv816 & c816);
  wire s817, sub817, and817, or817;
  wire b_inv817;
  assign b_inv817 = ~b817;
  assign s817  = a817 ^ b817 ^ c817;
  assign sub817 = a817 ^ b_inv817 ^ c817;
  assign and817 = a817 & b817;
  assign or817  = a817 | b817;
  assign c818 = (a817 & b817) | (a817 & c817) | (b817 & c817);
  wire c_sub818;
  assign c_sub818 = (a817 & b_inv817) | (a817 & c817) | (b_inv817 & c817);
  wire s818, sub818, and818, or818;
  wire b_inv818;
  assign b_inv818 = ~b818;
  assign s818  = a818 ^ b818 ^ c818;
  assign sub818 = a818 ^ b_inv818 ^ c818;
  assign and818 = a818 & b818;
  assign or818  = a818 | b818;
  assign c819 = (a818 & b818) | (a818 & c818) | (b818 & c818);
  wire c_sub819;
  assign c_sub819 = (a818 & b_inv818) | (a818 & c818) | (b_inv818 & c818);
  wire s819, sub819, and819, or819;
  wire b_inv819;
  assign b_inv819 = ~b819;
  assign s819  = a819 ^ b819 ^ c819;
  assign sub819 = a819 ^ b_inv819 ^ c819;
  assign and819 = a819 & b819;
  assign or819  = a819 | b819;
  assign c820 = (a819 & b819) | (a819 & c819) | (b819 & c819);
  wire c_sub820;
  assign c_sub820 = (a819 & b_inv819) | (a819 & c819) | (b_inv819 & c819);
  wire s820, sub820, and820, or820;
  wire b_inv820;
  assign b_inv820 = ~b820;
  assign s820  = a820 ^ b820 ^ c820;
  assign sub820 = a820 ^ b_inv820 ^ c820;
  assign and820 = a820 & b820;
  assign or820  = a820 | b820;
  assign c821 = (a820 & b820) | (a820 & c820) | (b820 & c820);
  wire c_sub821;
  assign c_sub821 = (a820 & b_inv820) | (a820 & c820) | (b_inv820 & c820);
  wire s821, sub821, and821, or821;
  wire b_inv821;
  assign b_inv821 = ~b821;
  assign s821  = a821 ^ b821 ^ c821;
  assign sub821 = a821 ^ b_inv821 ^ c821;
  assign and821 = a821 & b821;
  assign or821  = a821 | b821;
  assign c822 = (a821 & b821) | (a821 & c821) | (b821 & c821);
  wire c_sub822;
  assign c_sub822 = (a821 & b_inv821) | (a821 & c821) | (b_inv821 & c821);
  wire s822, sub822, and822, or822;
  wire b_inv822;
  assign b_inv822 = ~b822;
  assign s822  = a822 ^ b822 ^ c822;
  assign sub822 = a822 ^ b_inv822 ^ c822;
  assign and822 = a822 & b822;
  assign or822  = a822 | b822;
  assign c823 = (a822 & b822) | (a822 & c822) | (b822 & c822);
  wire c_sub823;
  assign c_sub823 = (a822 & b_inv822) | (a822 & c822) | (b_inv822 & c822);
  wire s823, sub823, and823, or823;
  wire b_inv823;
  assign b_inv823 = ~b823;
  assign s823  = a823 ^ b823 ^ c823;
  assign sub823 = a823 ^ b_inv823 ^ c823;
  assign and823 = a823 & b823;
  assign or823  = a823 | b823;
  assign c824 = (a823 & b823) | (a823 & c823) | (b823 & c823);
  wire c_sub824;
  assign c_sub824 = (a823 & b_inv823) | (a823 & c823) | (b_inv823 & c823);
  wire s824, sub824, and824, or824;
  wire b_inv824;
  assign b_inv824 = ~b824;
  assign s824  = a824 ^ b824 ^ c824;
  assign sub824 = a824 ^ b_inv824 ^ c824;
  assign and824 = a824 & b824;
  assign or824  = a824 | b824;
  assign c825 = (a824 & b824) | (a824 & c824) | (b824 & c824);
  wire c_sub825;
  assign c_sub825 = (a824 & b_inv824) | (a824 & c824) | (b_inv824 & c824);
  wire s825, sub825, and825, or825;
  wire b_inv825;
  assign b_inv825 = ~b825;
  assign s825  = a825 ^ b825 ^ c825;
  assign sub825 = a825 ^ b_inv825 ^ c825;
  assign and825 = a825 & b825;
  assign or825  = a825 | b825;
  assign c826 = (a825 & b825) | (a825 & c825) | (b825 & c825);
  wire c_sub826;
  assign c_sub826 = (a825 & b_inv825) | (a825 & c825) | (b_inv825 & c825);
  wire s826, sub826, and826, or826;
  wire b_inv826;
  assign b_inv826 = ~b826;
  assign s826  = a826 ^ b826 ^ c826;
  assign sub826 = a826 ^ b_inv826 ^ c826;
  assign and826 = a826 & b826;
  assign or826  = a826 | b826;
  assign c827 = (a826 & b826) | (a826 & c826) | (b826 & c826);
  wire c_sub827;
  assign c_sub827 = (a826 & b_inv826) | (a826 & c826) | (b_inv826 & c826);
  wire s827, sub827, and827, or827;
  wire b_inv827;
  assign b_inv827 = ~b827;
  assign s827  = a827 ^ b827 ^ c827;
  assign sub827 = a827 ^ b_inv827 ^ c827;
  assign and827 = a827 & b827;
  assign or827  = a827 | b827;
  assign c828 = (a827 & b827) | (a827 & c827) | (b827 & c827);
  wire c_sub828;
  assign c_sub828 = (a827 & b_inv827) | (a827 & c827) | (b_inv827 & c827);
  wire s828, sub828, and828, or828;
  wire b_inv828;
  assign b_inv828 = ~b828;
  assign s828  = a828 ^ b828 ^ c828;
  assign sub828 = a828 ^ b_inv828 ^ c828;
  assign and828 = a828 & b828;
  assign or828  = a828 | b828;
  assign c829 = (a828 & b828) | (a828 & c828) | (b828 & c828);
  wire c_sub829;
  assign c_sub829 = (a828 & b_inv828) | (a828 & c828) | (b_inv828 & c828);
  wire s829, sub829, and829, or829;
  wire b_inv829;
  assign b_inv829 = ~b829;
  assign s829  = a829 ^ b829 ^ c829;
  assign sub829 = a829 ^ b_inv829 ^ c829;
  assign and829 = a829 & b829;
  assign or829  = a829 | b829;
  assign c830 = (a829 & b829) | (a829 & c829) | (b829 & c829);
  wire c_sub830;
  assign c_sub830 = (a829 & b_inv829) | (a829 & c829) | (b_inv829 & c829);
  wire s830, sub830, and830, or830;
  wire b_inv830;
  assign b_inv830 = ~b830;
  assign s830  = a830 ^ b830 ^ c830;
  assign sub830 = a830 ^ b_inv830 ^ c830;
  assign and830 = a830 & b830;
  assign or830  = a830 | b830;
  assign c831 = (a830 & b830) | (a830 & c830) | (b830 & c830);
  wire c_sub831;
  assign c_sub831 = (a830 & b_inv830) | (a830 & c830) | (b_inv830 & c830);
  wire s831, sub831, and831, or831;
  wire b_inv831;
  assign b_inv831 = ~b831;
  assign s831  = a831 ^ b831 ^ c831;
  assign sub831 = a831 ^ b_inv831 ^ c831;
  assign and831 = a831 & b831;
  assign or831  = a831 | b831;
  assign c832 = (a831 & b831) | (a831 & c831) | (b831 & c831);
  wire c_sub832;
  assign c_sub832 = (a831 & b_inv831) | (a831 & c831) | (b_inv831 & c831);
  wire s832, sub832, and832, or832;
  wire b_inv832;
  assign b_inv832 = ~b832;
  assign s832  = a832 ^ b832 ^ c832;
  assign sub832 = a832 ^ b_inv832 ^ c832;
  assign and832 = a832 & b832;
  assign or832  = a832 | b832;
  assign c833 = (a832 & b832) | (a832 & c832) | (b832 & c832);
  wire c_sub833;
  assign c_sub833 = (a832 & b_inv832) | (a832 & c832) | (b_inv832 & c832);
  wire s833, sub833, and833, or833;
  wire b_inv833;
  assign b_inv833 = ~b833;
  assign s833  = a833 ^ b833 ^ c833;
  assign sub833 = a833 ^ b_inv833 ^ c833;
  assign and833 = a833 & b833;
  assign or833  = a833 | b833;
  assign c834 = (a833 & b833) | (a833 & c833) | (b833 & c833);
  wire c_sub834;
  assign c_sub834 = (a833 & b_inv833) | (a833 & c833) | (b_inv833 & c833);
  wire s834, sub834, and834, or834;
  wire b_inv834;
  assign b_inv834 = ~b834;
  assign s834  = a834 ^ b834 ^ c834;
  assign sub834 = a834 ^ b_inv834 ^ c834;
  assign and834 = a834 & b834;
  assign or834  = a834 | b834;
  assign c835 = (a834 & b834) | (a834 & c834) | (b834 & c834);
  wire c_sub835;
  assign c_sub835 = (a834 & b_inv834) | (a834 & c834) | (b_inv834 & c834);
  wire s835, sub835, and835, or835;
  wire b_inv835;
  assign b_inv835 = ~b835;
  assign s835  = a835 ^ b835 ^ c835;
  assign sub835 = a835 ^ b_inv835 ^ c835;
  assign and835 = a835 & b835;
  assign or835  = a835 | b835;
  assign c836 = (a835 & b835) | (a835 & c835) | (b835 & c835);
  wire c_sub836;
  assign c_sub836 = (a835 & b_inv835) | (a835 & c835) | (b_inv835 & c835);
  wire s836, sub836, and836, or836;
  wire b_inv836;
  assign b_inv836 = ~b836;
  assign s836  = a836 ^ b836 ^ c836;
  assign sub836 = a836 ^ b_inv836 ^ c836;
  assign and836 = a836 & b836;
  assign or836  = a836 | b836;
  assign c837 = (a836 & b836) | (a836 & c836) | (b836 & c836);
  wire c_sub837;
  assign c_sub837 = (a836 & b_inv836) | (a836 & c836) | (b_inv836 & c836);
  wire s837, sub837, and837, or837;
  wire b_inv837;
  assign b_inv837 = ~b837;
  assign s837  = a837 ^ b837 ^ c837;
  assign sub837 = a837 ^ b_inv837 ^ c837;
  assign and837 = a837 & b837;
  assign or837  = a837 | b837;
  assign c838 = (a837 & b837) | (a837 & c837) | (b837 & c837);
  wire c_sub838;
  assign c_sub838 = (a837 & b_inv837) | (a837 & c837) | (b_inv837 & c837);
  wire s838, sub838, and838, or838;
  wire b_inv838;
  assign b_inv838 = ~b838;
  assign s838  = a838 ^ b838 ^ c838;
  assign sub838 = a838 ^ b_inv838 ^ c838;
  assign and838 = a838 & b838;
  assign or838  = a838 | b838;
  assign c839 = (a838 & b838) | (a838 & c838) | (b838 & c838);
  wire c_sub839;
  assign c_sub839 = (a838 & b_inv838) | (a838 & c838) | (b_inv838 & c838);
  wire s839, sub839, and839, or839;
  wire b_inv839;
  assign b_inv839 = ~b839;
  assign s839  = a839 ^ b839 ^ c839;
  assign sub839 = a839 ^ b_inv839 ^ c839;
  assign and839 = a839 & b839;
  assign or839  = a839 | b839;
  assign c840 = (a839 & b839) | (a839 & c839) | (b839 & c839);
  wire c_sub840;
  assign c_sub840 = (a839 & b_inv839) | (a839 & c839) | (b_inv839 & c839);
  wire s840, sub840, and840, or840;
  wire b_inv840;
  assign b_inv840 = ~b840;
  assign s840  = a840 ^ b840 ^ c840;
  assign sub840 = a840 ^ b_inv840 ^ c840;
  assign and840 = a840 & b840;
  assign or840  = a840 | b840;
  assign c841 = (a840 & b840) | (a840 & c840) | (b840 & c840);
  wire c_sub841;
  assign c_sub841 = (a840 & b_inv840) | (a840 & c840) | (b_inv840 & c840);
  wire s841, sub841, and841, or841;
  wire b_inv841;
  assign b_inv841 = ~b841;
  assign s841  = a841 ^ b841 ^ c841;
  assign sub841 = a841 ^ b_inv841 ^ c841;
  assign and841 = a841 & b841;
  assign or841  = a841 | b841;
  assign c842 = (a841 & b841) | (a841 & c841) | (b841 & c841);
  wire c_sub842;
  assign c_sub842 = (a841 & b_inv841) | (a841 & c841) | (b_inv841 & c841);
  wire s842, sub842, and842, or842;
  wire b_inv842;
  assign b_inv842 = ~b842;
  assign s842  = a842 ^ b842 ^ c842;
  assign sub842 = a842 ^ b_inv842 ^ c842;
  assign and842 = a842 & b842;
  assign or842  = a842 | b842;
  assign c843 = (a842 & b842) | (a842 & c842) | (b842 & c842);
  wire c_sub843;
  assign c_sub843 = (a842 & b_inv842) | (a842 & c842) | (b_inv842 & c842);
  wire s843, sub843, and843, or843;
  wire b_inv843;
  assign b_inv843 = ~b843;
  assign s843  = a843 ^ b843 ^ c843;
  assign sub843 = a843 ^ b_inv843 ^ c843;
  assign and843 = a843 & b843;
  assign or843  = a843 | b843;
  assign c844 = (a843 & b843) | (a843 & c843) | (b843 & c843);
  wire c_sub844;
  assign c_sub844 = (a843 & b_inv843) | (a843 & c843) | (b_inv843 & c843);
  wire s844, sub844, and844, or844;
  wire b_inv844;
  assign b_inv844 = ~b844;
  assign s844  = a844 ^ b844 ^ c844;
  assign sub844 = a844 ^ b_inv844 ^ c844;
  assign and844 = a844 & b844;
  assign or844  = a844 | b844;
  assign c845 = (a844 & b844) | (a844 & c844) | (b844 & c844);
  wire c_sub845;
  assign c_sub845 = (a844 & b_inv844) | (a844 & c844) | (b_inv844 & c844);
  wire s845, sub845, and845, or845;
  wire b_inv845;
  assign b_inv845 = ~b845;
  assign s845  = a845 ^ b845 ^ c845;
  assign sub845 = a845 ^ b_inv845 ^ c845;
  assign and845 = a845 & b845;
  assign or845  = a845 | b845;
  assign c846 = (a845 & b845) | (a845 & c845) | (b845 & c845);
  wire c_sub846;
  assign c_sub846 = (a845 & b_inv845) | (a845 & c845) | (b_inv845 & c845);
  wire s846, sub846, and846, or846;
  wire b_inv846;
  assign b_inv846 = ~b846;
  assign s846  = a846 ^ b846 ^ c846;
  assign sub846 = a846 ^ b_inv846 ^ c846;
  assign and846 = a846 & b846;
  assign or846  = a846 | b846;
  assign c847 = (a846 & b846) | (a846 & c846) | (b846 & c846);
  wire c_sub847;
  assign c_sub847 = (a846 & b_inv846) | (a846 & c846) | (b_inv846 & c846);
  wire s847, sub847, and847, or847;
  wire b_inv847;
  assign b_inv847 = ~b847;
  assign s847  = a847 ^ b847 ^ c847;
  assign sub847 = a847 ^ b_inv847 ^ c847;
  assign and847 = a847 & b847;
  assign or847  = a847 | b847;
  assign c848 = (a847 & b847) | (a847 & c847) | (b847 & c847);
  wire c_sub848;
  assign c_sub848 = (a847 & b_inv847) | (a847 & c847) | (b_inv847 & c847);
  wire s848, sub848, and848, or848;
  wire b_inv848;
  assign b_inv848 = ~b848;
  assign s848  = a848 ^ b848 ^ c848;
  assign sub848 = a848 ^ b_inv848 ^ c848;
  assign and848 = a848 & b848;
  assign or848  = a848 | b848;
  assign c849 = (a848 & b848) | (a848 & c848) | (b848 & c848);
  wire c_sub849;
  assign c_sub849 = (a848 & b_inv848) | (a848 & c848) | (b_inv848 & c848);
  wire s849, sub849, and849, or849;
  wire b_inv849;
  assign b_inv849 = ~b849;
  assign s849  = a849 ^ b849 ^ c849;
  assign sub849 = a849 ^ b_inv849 ^ c849;
  assign and849 = a849 & b849;
  assign or849  = a849 | b849;
  assign c850 = (a849 & b849) | (a849 & c849) | (b849 & c849);
  wire c_sub850;
  assign c_sub850 = (a849 & b_inv849) | (a849 & c849) | (b_inv849 & c849);
  wire s850, sub850, and850, or850;
  wire b_inv850;
  assign b_inv850 = ~b850;
  assign s850  = a850 ^ b850 ^ c850;
  assign sub850 = a850 ^ b_inv850 ^ c850;
  assign and850 = a850 & b850;
  assign or850  = a850 | b850;
  assign c851 = (a850 & b850) | (a850 & c850) | (b850 & c850);
  wire c_sub851;
  assign c_sub851 = (a850 & b_inv850) | (a850 & c850) | (b_inv850 & c850);
  wire s851, sub851, and851, or851;
  wire b_inv851;
  assign b_inv851 = ~b851;
  assign s851  = a851 ^ b851 ^ c851;
  assign sub851 = a851 ^ b_inv851 ^ c851;
  assign and851 = a851 & b851;
  assign or851  = a851 | b851;
  assign c852 = (a851 & b851) | (a851 & c851) | (b851 & c851);
  wire c_sub852;
  assign c_sub852 = (a851 & b_inv851) | (a851 & c851) | (b_inv851 & c851);
  wire s852, sub852, and852, or852;
  wire b_inv852;
  assign b_inv852 = ~b852;
  assign s852  = a852 ^ b852 ^ c852;
  assign sub852 = a852 ^ b_inv852 ^ c852;
  assign and852 = a852 & b852;
  assign or852  = a852 | b852;
  assign c853 = (a852 & b852) | (a852 & c852) | (b852 & c852);
  wire c_sub853;
  assign c_sub853 = (a852 & b_inv852) | (a852 & c852) | (b_inv852 & c852);
  wire s853, sub853, and853, or853;
  wire b_inv853;
  assign b_inv853 = ~b853;
  assign s853  = a853 ^ b853 ^ c853;
  assign sub853 = a853 ^ b_inv853 ^ c853;
  assign and853 = a853 & b853;
  assign or853  = a853 | b853;
  assign c854 = (a853 & b853) | (a853 & c853) | (b853 & c853);
  wire c_sub854;
  assign c_sub854 = (a853 & b_inv853) | (a853 & c853) | (b_inv853 & c853);
  wire s854, sub854, and854, or854;
  wire b_inv854;
  assign b_inv854 = ~b854;
  assign s854  = a854 ^ b854 ^ c854;
  assign sub854 = a854 ^ b_inv854 ^ c854;
  assign and854 = a854 & b854;
  assign or854  = a854 | b854;
  assign c855 = (a854 & b854) | (a854 & c854) | (b854 & c854);
  wire c_sub855;
  assign c_sub855 = (a854 & b_inv854) | (a854 & c854) | (b_inv854 & c854);
  wire s855, sub855, and855, or855;
  wire b_inv855;
  assign b_inv855 = ~b855;
  assign s855  = a855 ^ b855 ^ c855;
  assign sub855 = a855 ^ b_inv855 ^ c855;
  assign and855 = a855 & b855;
  assign or855  = a855 | b855;
  assign c856 = (a855 & b855) | (a855 & c855) | (b855 & c855);
  wire c_sub856;
  assign c_sub856 = (a855 & b_inv855) | (a855 & c855) | (b_inv855 & c855);
  wire s856, sub856, and856, or856;
  wire b_inv856;
  assign b_inv856 = ~b856;
  assign s856  = a856 ^ b856 ^ c856;
  assign sub856 = a856 ^ b_inv856 ^ c856;
  assign and856 = a856 & b856;
  assign or856  = a856 | b856;
  assign c857 = (a856 & b856) | (a856 & c856) | (b856 & c856);
  wire c_sub857;
  assign c_sub857 = (a856 & b_inv856) | (a856 & c856) | (b_inv856 & c856);
  wire s857, sub857, and857, or857;
  wire b_inv857;
  assign b_inv857 = ~b857;
  assign s857  = a857 ^ b857 ^ c857;
  assign sub857 = a857 ^ b_inv857 ^ c857;
  assign and857 = a857 & b857;
  assign or857  = a857 | b857;
  assign c858 = (a857 & b857) | (a857 & c857) | (b857 & c857);
  wire c_sub858;
  assign c_sub858 = (a857 & b_inv857) | (a857 & c857) | (b_inv857 & c857);
  wire s858, sub858, and858, or858;
  wire b_inv858;
  assign b_inv858 = ~b858;
  assign s858  = a858 ^ b858 ^ c858;
  assign sub858 = a858 ^ b_inv858 ^ c858;
  assign and858 = a858 & b858;
  assign or858  = a858 | b858;
  assign c859 = (a858 & b858) | (a858 & c858) | (b858 & c858);
  wire c_sub859;
  assign c_sub859 = (a858 & b_inv858) | (a858 & c858) | (b_inv858 & c858);
  wire s859, sub859, and859, or859;
  wire b_inv859;
  assign b_inv859 = ~b859;
  assign s859  = a859 ^ b859 ^ c859;
  assign sub859 = a859 ^ b_inv859 ^ c859;
  assign and859 = a859 & b859;
  assign or859  = a859 | b859;
  assign c860 = (a859 & b859) | (a859 & c859) | (b859 & c859);
  wire c_sub860;
  assign c_sub860 = (a859 & b_inv859) | (a859 & c859) | (b_inv859 & c859);
  wire s860, sub860, and860, or860;
  wire b_inv860;
  assign b_inv860 = ~b860;
  assign s860  = a860 ^ b860 ^ c860;
  assign sub860 = a860 ^ b_inv860 ^ c860;
  assign and860 = a860 & b860;
  assign or860  = a860 | b860;
  assign c861 = (a860 & b860) | (a860 & c860) | (b860 & c860);
  wire c_sub861;
  assign c_sub861 = (a860 & b_inv860) | (a860 & c860) | (b_inv860 & c860);
  wire s861, sub861, and861, or861;
  wire b_inv861;
  assign b_inv861 = ~b861;
  assign s861  = a861 ^ b861 ^ c861;
  assign sub861 = a861 ^ b_inv861 ^ c861;
  assign and861 = a861 & b861;
  assign or861  = a861 | b861;
  assign c862 = (a861 & b861) | (a861 & c861) | (b861 & c861);
  wire c_sub862;
  assign c_sub862 = (a861 & b_inv861) | (a861 & c861) | (b_inv861 & c861);
  wire s862, sub862, and862, or862;
  wire b_inv862;
  assign b_inv862 = ~b862;
  assign s862  = a862 ^ b862 ^ c862;
  assign sub862 = a862 ^ b_inv862 ^ c862;
  assign and862 = a862 & b862;
  assign or862  = a862 | b862;
  assign c863 = (a862 & b862) | (a862 & c862) | (b862 & c862);
  wire c_sub863;
  assign c_sub863 = (a862 & b_inv862) | (a862 & c862) | (b_inv862 & c862);
  wire s863, sub863, and863, or863;
  wire b_inv863;
  assign b_inv863 = ~b863;
  assign s863  = a863 ^ b863 ^ c863;
  assign sub863 = a863 ^ b_inv863 ^ c863;
  assign and863 = a863 & b863;
  assign or863  = a863 | b863;
  assign c864 = (a863 & b863) | (a863 & c863) | (b863 & c863);
  wire c_sub864;
  assign c_sub864 = (a863 & b_inv863) | (a863 & c863) | (b_inv863 & c863);
  wire s864, sub864, and864, or864;
  wire b_inv864;
  assign b_inv864 = ~b864;
  assign s864  = a864 ^ b864 ^ c864;
  assign sub864 = a864 ^ b_inv864 ^ c864;
  assign and864 = a864 & b864;
  assign or864  = a864 | b864;
  assign c865 = (a864 & b864) | (a864 & c864) | (b864 & c864);
  wire c_sub865;
  assign c_sub865 = (a864 & b_inv864) | (a864 & c864) | (b_inv864 & c864);
  wire s865, sub865, and865, or865;
  wire b_inv865;
  assign b_inv865 = ~b865;
  assign s865  = a865 ^ b865 ^ c865;
  assign sub865 = a865 ^ b_inv865 ^ c865;
  assign and865 = a865 & b865;
  assign or865  = a865 | b865;
  assign c866 = (a865 & b865) | (a865 & c865) | (b865 & c865);
  wire c_sub866;
  assign c_sub866 = (a865 & b_inv865) | (a865 & c865) | (b_inv865 & c865);
  wire s866, sub866, and866, or866;
  wire b_inv866;
  assign b_inv866 = ~b866;
  assign s866  = a866 ^ b866 ^ c866;
  assign sub866 = a866 ^ b_inv866 ^ c866;
  assign and866 = a866 & b866;
  assign or866  = a866 | b866;
  assign c867 = (a866 & b866) | (a866 & c866) | (b866 & c866);
  wire c_sub867;
  assign c_sub867 = (a866 & b_inv866) | (a866 & c866) | (b_inv866 & c866);
  wire s867, sub867, and867, or867;
  wire b_inv867;
  assign b_inv867 = ~b867;
  assign s867  = a867 ^ b867 ^ c867;
  assign sub867 = a867 ^ b_inv867 ^ c867;
  assign and867 = a867 & b867;
  assign or867  = a867 | b867;
  assign c868 = (a867 & b867) | (a867 & c867) | (b867 & c867);
  wire c_sub868;
  assign c_sub868 = (a867 & b_inv867) | (a867 & c867) | (b_inv867 & c867);
  wire s868, sub868, and868, or868;
  wire b_inv868;
  assign b_inv868 = ~b868;
  assign s868  = a868 ^ b868 ^ c868;
  assign sub868 = a868 ^ b_inv868 ^ c868;
  assign and868 = a868 & b868;
  assign or868  = a868 | b868;
  assign c869 = (a868 & b868) | (a868 & c868) | (b868 & c868);
  wire c_sub869;
  assign c_sub869 = (a868 & b_inv868) | (a868 & c868) | (b_inv868 & c868);
  wire s869, sub869, and869, or869;
  wire b_inv869;
  assign b_inv869 = ~b869;
  assign s869  = a869 ^ b869 ^ c869;
  assign sub869 = a869 ^ b_inv869 ^ c869;
  assign and869 = a869 & b869;
  assign or869  = a869 | b869;
  assign c870 = (a869 & b869) | (a869 & c869) | (b869 & c869);
  wire c_sub870;
  assign c_sub870 = (a869 & b_inv869) | (a869 & c869) | (b_inv869 & c869);
  wire s870, sub870, and870, or870;
  wire b_inv870;
  assign b_inv870 = ~b870;
  assign s870  = a870 ^ b870 ^ c870;
  assign sub870 = a870 ^ b_inv870 ^ c870;
  assign and870 = a870 & b870;
  assign or870  = a870 | b870;
  assign c871 = (a870 & b870) | (a870 & c870) | (b870 & c870);
  wire c_sub871;
  assign c_sub871 = (a870 & b_inv870) | (a870 & c870) | (b_inv870 & c870);
  wire s871, sub871, and871, or871;
  wire b_inv871;
  assign b_inv871 = ~b871;
  assign s871  = a871 ^ b871 ^ c871;
  assign sub871 = a871 ^ b_inv871 ^ c871;
  assign and871 = a871 & b871;
  assign or871  = a871 | b871;
  assign c872 = (a871 & b871) | (a871 & c871) | (b871 & c871);
  wire c_sub872;
  assign c_sub872 = (a871 & b_inv871) | (a871 & c871) | (b_inv871 & c871);
  wire s872, sub872, and872, or872;
  wire b_inv872;
  assign b_inv872 = ~b872;
  assign s872  = a872 ^ b872 ^ c872;
  assign sub872 = a872 ^ b_inv872 ^ c872;
  assign and872 = a872 & b872;
  assign or872  = a872 | b872;
  assign c873 = (a872 & b872) | (a872 & c872) | (b872 & c872);
  wire c_sub873;
  assign c_sub873 = (a872 & b_inv872) | (a872 & c872) | (b_inv872 & c872);
  wire s873, sub873, and873, or873;
  wire b_inv873;
  assign b_inv873 = ~b873;
  assign s873  = a873 ^ b873 ^ c873;
  assign sub873 = a873 ^ b_inv873 ^ c873;
  assign and873 = a873 & b873;
  assign or873  = a873 | b873;
  assign c874 = (a873 & b873) | (a873 & c873) | (b873 & c873);
  wire c_sub874;
  assign c_sub874 = (a873 & b_inv873) | (a873 & c873) | (b_inv873 & c873);
  wire s874, sub874, and874, or874;
  wire b_inv874;
  assign b_inv874 = ~b874;
  assign s874  = a874 ^ b874 ^ c874;
  assign sub874 = a874 ^ b_inv874 ^ c874;
  assign and874 = a874 & b874;
  assign or874  = a874 | b874;
  assign c875 = (a874 & b874) | (a874 & c874) | (b874 & c874);
  wire c_sub875;
  assign c_sub875 = (a874 & b_inv874) | (a874 & c874) | (b_inv874 & c874);
  wire s875, sub875, and875, or875;
  wire b_inv875;
  assign b_inv875 = ~b875;
  assign s875  = a875 ^ b875 ^ c875;
  assign sub875 = a875 ^ b_inv875 ^ c875;
  assign and875 = a875 & b875;
  assign or875  = a875 | b875;
  assign c876 = (a875 & b875) | (a875 & c875) | (b875 & c875);
  wire c_sub876;
  assign c_sub876 = (a875 & b_inv875) | (a875 & c875) | (b_inv875 & c875);
  wire s876, sub876, and876, or876;
  wire b_inv876;
  assign b_inv876 = ~b876;
  assign s876  = a876 ^ b876 ^ c876;
  assign sub876 = a876 ^ b_inv876 ^ c876;
  assign and876 = a876 & b876;
  assign or876  = a876 | b876;
  assign c877 = (a876 & b876) | (a876 & c876) | (b876 & c876);
  wire c_sub877;
  assign c_sub877 = (a876 & b_inv876) | (a876 & c876) | (b_inv876 & c876);
  wire s877, sub877, and877, or877;
  wire b_inv877;
  assign b_inv877 = ~b877;
  assign s877  = a877 ^ b877 ^ c877;
  assign sub877 = a877 ^ b_inv877 ^ c877;
  assign and877 = a877 & b877;
  assign or877  = a877 | b877;
  assign c878 = (a877 & b877) | (a877 & c877) | (b877 & c877);
  wire c_sub878;
  assign c_sub878 = (a877 & b_inv877) | (a877 & c877) | (b_inv877 & c877);
  wire s878, sub878, and878, or878;
  wire b_inv878;
  assign b_inv878 = ~b878;
  assign s878  = a878 ^ b878 ^ c878;
  assign sub878 = a878 ^ b_inv878 ^ c878;
  assign and878 = a878 & b878;
  assign or878  = a878 | b878;
  assign c879 = (a878 & b878) | (a878 & c878) | (b878 & c878);
  wire c_sub879;
  assign c_sub879 = (a878 & b_inv878) | (a878 & c878) | (b_inv878 & c878);
  wire s879, sub879, and879, or879;
  wire b_inv879;
  assign b_inv879 = ~b879;
  assign s879  = a879 ^ b879 ^ c879;
  assign sub879 = a879 ^ b_inv879 ^ c879;
  assign and879 = a879 & b879;
  assign or879  = a879 | b879;
  assign c880 = (a879 & b879) | (a879 & c879) | (b879 & c879);
  wire c_sub880;
  assign c_sub880 = (a879 & b_inv879) | (a879 & c879) | (b_inv879 & c879);
  wire s880, sub880, and880, or880;
  wire b_inv880;
  assign b_inv880 = ~b880;
  assign s880  = a880 ^ b880 ^ c880;
  assign sub880 = a880 ^ b_inv880 ^ c880;
  assign and880 = a880 & b880;
  assign or880  = a880 | b880;
  assign c881 = (a880 & b880) | (a880 & c880) | (b880 & c880);
  wire c_sub881;
  assign c_sub881 = (a880 & b_inv880) | (a880 & c880) | (b_inv880 & c880);
  wire s881, sub881, and881, or881;
  wire b_inv881;
  assign b_inv881 = ~b881;
  assign s881  = a881 ^ b881 ^ c881;
  assign sub881 = a881 ^ b_inv881 ^ c881;
  assign and881 = a881 & b881;
  assign or881  = a881 | b881;
  assign c882 = (a881 & b881) | (a881 & c881) | (b881 & c881);
  wire c_sub882;
  assign c_sub882 = (a881 & b_inv881) | (a881 & c881) | (b_inv881 & c881);
  wire s882, sub882, and882, or882;
  wire b_inv882;
  assign b_inv882 = ~b882;
  assign s882  = a882 ^ b882 ^ c882;
  assign sub882 = a882 ^ b_inv882 ^ c882;
  assign and882 = a882 & b882;
  assign or882  = a882 | b882;
  assign c883 = (a882 & b882) | (a882 & c882) | (b882 & c882);
  wire c_sub883;
  assign c_sub883 = (a882 & b_inv882) | (a882 & c882) | (b_inv882 & c882);
  wire s883, sub883, and883, or883;
  wire b_inv883;
  assign b_inv883 = ~b883;
  assign s883  = a883 ^ b883 ^ c883;
  assign sub883 = a883 ^ b_inv883 ^ c883;
  assign and883 = a883 & b883;
  assign or883  = a883 | b883;
  assign c884 = (a883 & b883) | (a883 & c883) | (b883 & c883);
  wire c_sub884;
  assign c_sub884 = (a883 & b_inv883) | (a883 & c883) | (b_inv883 & c883);
  wire s884, sub884, and884, or884;
  wire b_inv884;
  assign b_inv884 = ~b884;
  assign s884  = a884 ^ b884 ^ c884;
  assign sub884 = a884 ^ b_inv884 ^ c884;
  assign and884 = a884 & b884;
  assign or884  = a884 | b884;
  assign c885 = (a884 & b884) | (a884 & c884) | (b884 & c884);
  wire c_sub885;
  assign c_sub885 = (a884 & b_inv884) | (a884 & c884) | (b_inv884 & c884);
  wire s885, sub885, and885, or885;
  wire b_inv885;
  assign b_inv885 = ~b885;
  assign s885  = a885 ^ b885 ^ c885;
  assign sub885 = a885 ^ b_inv885 ^ c885;
  assign and885 = a885 & b885;
  assign or885  = a885 | b885;
  assign c886 = (a885 & b885) | (a885 & c885) | (b885 & c885);
  wire c_sub886;
  assign c_sub886 = (a885 & b_inv885) | (a885 & c885) | (b_inv885 & c885);
  wire s886, sub886, and886, or886;
  wire b_inv886;
  assign b_inv886 = ~b886;
  assign s886  = a886 ^ b886 ^ c886;
  assign sub886 = a886 ^ b_inv886 ^ c886;
  assign and886 = a886 & b886;
  assign or886  = a886 | b886;
  assign c887 = (a886 & b886) | (a886 & c886) | (b886 & c886);
  wire c_sub887;
  assign c_sub887 = (a886 & b_inv886) | (a886 & c886) | (b_inv886 & c886);
  wire s887, sub887, and887, or887;
  wire b_inv887;
  assign b_inv887 = ~b887;
  assign s887  = a887 ^ b887 ^ c887;
  assign sub887 = a887 ^ b_inv887 ^ c887;
  assign and887 = a887 & b887;
  assign or887  = a887 | b887;
  assign c888 = (a887 & b887) | (a887 & c887) | (b887 & c887);
  wire c_sub888;
  assign c_sub888 = (a887 & b_inv887) | (a887 & c887) | (b_inv887 & c887);
  wire s888, sub888, and888, or888;
  wire b_inv888;
  assign b_inv888 = ~b888;
  assign s888  = a888 ^ b888 ^ c888;
  assign sub888 = a888 ^ b_inv888 ^ c888;
  assign and888 = a888 & b888;
  assign or888  = a888 | b888;
  assign c889 = (a888 & b888) | (a888 & c888) | (b888 & c888);
  wire c_sub889;
  assign c_sub889 = (a888 & b_inv888) | (a888 & c888) | (b_inv888 & c888);
  wire s889, sub889, and889, or889;
  wire b_inv889;
  assign b_inv889 = ~b889;
  assign s889  = a889 ^ b889 ^ c889;
  assign sub889 = a889 ^ b_inv889 ^ c889;
  assign and889 = a889 & b889;
  assign or889  = a889 | b889;
  assign c890 = (a889 & b889) | (a889 & c889) | (b889 & c889);
  wire c_sub890;
  assign c_sub890 = (a889 & b_inv889) | (a889 & c889) | (b_inv889 & c889);
  wire s890, sub890, and890, or890;
  wire b_inv890;
  assign b_inv890 = ~b890;
  assign s890  = a890 ^ b890 ^ c890;
  assign sub890 = a890 ^ b_inv890 ^ c890;
  assign and890 = a890 & b890;
  assign or890  = a890 | b890;
  assign c891 = (a890 & b890) | (a890 & c890) | (b890 & c890);
  wire c_sub891;
  assign c_sub891 = (a890 & b_inv890) | (a890 & c890) | (b_inv890 & c890);
  wire s891, sub891, and891, or891;
  wire b_inv891;
  assign b_inv891 = ~b891;
  assign s891  = a891 ^ b891 ^ c891;
  assign sub891 = a891 ^ b_inv891 ^ c891;
  assign and891 = a891 & b891;
  assign or891  = a891 | b891;
  assign c892 = (a891 & b891) | (a891 & c891) | (b891 & c891);
  wire c_sub892;
  assign c_sub892 = (a891 & b_inv891) | (a891 & c891) | (b_inv891 & c891);
  wire s892, sub892, and892, or892;
  wire b_inv892;
  assign b_inv892 = ~b892;
  assign s892  = a892 ^ b892 ^ c892;
  assign sub892 = a892 ^ b_inv892 ^ c892;
  assign and892 = a892 & b892;
  assign or892  = a892 | b892;
  assign c893 = (a892 & b892) | (a892 & c892) | (b892 & c892);
  wire c_sub893;
  assign c_sub893 = (a892 & b_inv892) | (a892 & c892) | (b_inv892 & c892);
  wire s893, sub893, and893, or893;
  wire b_inv893;
  assign b_inv893 = ~b893;
  assign s893  = a893 ^ b893 ^ c893;
  assign sub893 = a893 ^ b_inv893 ^ c893;
  assign and893 = a893 & b893;
  assign or893  = a893 | b893;
  assign c894 = (a893 & b893) | (a893 & c893) | (b893 & c893);
  wire c_sub894;
  assign c_sub894 = (a893 & b_inv893) | (a893 & c893) | (b_inv893 & c893);
  wire s894, sub894, and894, or894;
  wire b_inv894;
  assign b_inv894 = ~b894;
  assign s894  = a894 ^ b894 ^ c894;
  assign sub894 = a894 ^ b_inv894 ^ c894;
  assign and894 = a894 & b894;
  assign or894  = a894 | b894;
  assign c895 = (a894 & b894) | (a894 & c894) | (b894 & c894);
  wire c_sub895;
  assign c_sub895 = (a894 & b_inv894) | (a894 & c894) | (b_inv894 & c894);
  wire s895, sub895, and895, or895;
  wire b_inv895;
  assign b_inv895 = ~b895;
  assign s895  = a895 ^ b895 ^ c895;
  assign sub895 = a895 ^ b_inv895 ^ c895;
  assign and895 = a895 & b895;
  assign or895  = a895 | b895;
  assign c896 = (a895 & b895) | (a895 & c895) | (b895 & c895);
  wire c_sub896;
  assign c_sub896 = (a895 & b_inv895) | (a895 & c895) | (b_inv895 & c895);
  wire s896, sub896, and896, or896;
  wire b_inv896;
  assign b_inv896 = ~b896;
  assign s896  = a896 ^ b896 ^ c896;
  assign sub896 = a896 ^ b_inv896 ^ c896;
  assign and896 = a896 & b896;
  assign or896  = a896 | b896;
  assign c897 = (a896 & b896) | (a896 & c896) | (b896 & c896);
  wire c_sub897;
  assign c_sub897 = (a896 & b_inv896) | (a896 & c896) | (b_inv896 & c896);
  wire s897, sub897, and897, or897;
  wire b_inv897;
  assign b_inv897 = ~b897;
  assign s897  = a897 ^ b897 ^ c897;
  assign sub897 = a897 ^ b_inv897 ^ c897;
  assign and897 = a897 & b897;
  assign or897  = a897 | b897;
  assign c898 = (a897 & b897) | (a897 & c897) | (b897 & c897);
  wire c_sub898;
  assign c_sub898 = (a897 & b_inv897) | (a897 & c897) | (b_inv897 & c897);
  wire s898, sub898, and898, or898;
  wire b_inv898;
  assign b_inv898 = ~b898;
  assign s898  = a898 ^ b898 ^ c898;
  assign sub898 = a898 ^ b_inv898 ^ c898;
  assign and898 = a898 & b898;
  assign or898  = a898 | b898;
  assign c899 = (a898 & b898) | (a898 & c898) | (b898 & c898);
  wire c_sub899;
  assign c_sub899 = (a898 & b_inv898) | (a898 & c898) | (b_inv898 & c898);
  wire s899, sub899, and899, or899;
  wire b_inv899;
  assign b_inv899 = ~b899;
  assign s899  = a899 ^ b899 ^ c899;
  assign sub899 = a899 ^ b_inv899 ^ c899;
  assign and899 = a899 & b899;
  assign or899  = a899 | b899;
  assign c900 = (a899 & b899) | (a899 & c899) | (b899 & c899);
  wire c_sub900;
  assign c_sub900 = (a899 & b_inv899) | (a899 & c899) | (b_inv899 & c899);
  wire s900, sub900, and900, or900;
  wire b_inv900;
  assign b_inv900 = ~b900;
  assign s900  = a900 ^ b900 ^ c900;
  assign sub900 = a900 ^ b_inv900 ^ c900;
  assign and900 = a900 & b900;
  assign or900  = a900 | b900;
  assign c901 = (a900 & b900) | (a900 & c900) | (b900 & c900);
  wire c_sub901;
  assign c_sub901 = (a900 & b_inv900) | (a900 & c900) | (b_inv900 & c900);
  wire s901, sub901, and901, or901;
  wire b_inv901;
  assign b_inv901 = ~b901;
  assign s901  = a901 ^ b901 ^ c901;
  assign sub901 = a901 ^ b_inv901 ^ c901;
  assign and901 = a901 & b901;
  assign or901  = a901 | b901;
  assign c902 = (a901 & b901) | (a901 & c901) | (b901 & c901);
  wire c_sub902;
  assign c_sub902 = (a901 & b_inv901) | (a901 & c901) | (b_inv901 & c901);
  wire s902, sub902, and902, or902;
  wire b_inv902;
  assign b_inv902 = ~b902;
  assign s902  = a902 ^ b902 ^ c902;
  assign sub902 = a902 ^ b_inv902 ^ c902;
  assign and902 = a902 & b902;
  assign or902  = a902 | b902;
  assign c903 = (a902 & b902) | (a902 & c902) | (b902 & c902);
  wire c_sub903;
  assign c_sub903 = (a902 & b_inv902) | (a902 & c902) | (b_inv902 & c902);
  wire s903, sub903, and903, or903;
  wire b_inv903;
  assign b_inv903 = ~b903;
  assign s903  = a903 ^ b903 ^ c903;
  assign sub903 = a903 ^ b_inv903 ^ c903;
  assign and903 = a903 & b903;
  assign or903  = a903 | b903;
  assign c904 = (a903 & b903) | (a903 & c903) | (b903 & c903);
  wire c_sub904;
  assign c_sub904 = (a903 & b_inv903) | (a903 & c903) | (b_inv903 & c903);
  wire s904, sub904, and904, or904;
  wire b_inv904;
  assign b_inv904 = ~b904;
  assign s904  = a904 ^ b904 ^ c904;
  assign sub904 = a904 ^ b_inv904 ^ c904;
  assign and904 = a904 & b904;
  assign or904  = a904 | b904;
  assign c905 = (a904 & b904) | (a904 & c904) | (b904 & c904);
  wire c_sub905;
  assign c_sub905 = (a904 & b_inv904) | (a904 & c904) | (b_inv904 & c904);
  wire s905, sub905, and905, or905;
  wire b_inv905;
  assign b_inv905 = ~b905;
  assign s905  = a905 ^ b905 ^ c905;
  assign sub905 = a905 ^ b_inv905 ^ c905;
  assign and905 = a905 & b905;
  assign or905  = a905 | b905;
  assign c906 = (a905 & b905) | (a905 & c905) | (b905 & c905);
  wire c_sub906;
  assign c_sub906 = (a905 & b_inv905) | (a905 & c905) | (b_inv905 & c905);
  wire s906, sub906, and906, or906;
  wire b_inv906;
  assign b_inv906 = ~b906;
  assign s906  = a906 ^ b906 ^ c906;
  assign sub906 = a906 ^ b_inv906 ^ c906;
  assign and906 = a906 & b906;
  assign or906  = a906 | b906;
  assign c907 = (a906 & b906) | (a906 & c906) | (b906 & c906);
  wire c_sub907;
  assign c_sub907 = (a906 & b_inv906) | (a906 & c906) | (b_inv906 & c906);
  wire s907, sub907, and907, or907;
  wire b_inv907;
  assign b_inv907 = ~b907;
  assign s907  = a907 ^ b907 ^ c907;
  assign sub907 = a907 ^ b_inv907 ^ c907;
  assign and907 = a907 & b907;
  assign or907  = a907 | b907;
  assign c908 = (a907 & b907) | (a907 & c907) | (b907 & c907);
  wire c_sub908;
  assign c_sub908 = (a907 & b_inv907) | (a907 & c907) | (b_inv907 & c907);
  wire s908, sub908, and908, or908;
  wire b_inv908;
  assign b_inv908 = ~b908;
  assign s908  = a908 ^ b908 ^ c908;
  assign sub908 = a908 ^ b_inv908 ^ c908;
  assign and908 = a908 & b908;
  assign or908  = a908 | b908;
  assign c909 = (a908 & b908) | (a908 & c908) | (b908 & c908);
  wire c_sub909;
  assign c_sub909 = (a908 & b_inv908) | (a908 & c908) | (b_inv908 & c908);
  wire s909, sub909, and909, or909;
  wire b_inv909;
  assign b_inv909 = ~b909;
  assign s909  = a909 ^ b909 ^ c909;
  assign sub909 = a909 ^ b_inv909 ^ c909;
  assign and909 = a909 & b909;
  assign or909  = a909 | b909;
  assign c910 = (a909 & b909) | (a909 & c909) | (b909 & c909);
  wire c_sub910;
  assign c_sub910 = (a909 & b_inv909) | (a909 & c909) | (b_inv909 & c909);
  wire s910, sub910, and910, or910;
  wire b_inv910;
  assign b_inv910 = ~b910;
  assign s910  = a910 ^ b910 ^ c910;
  assign sub910 = a910 ^ b_inv910 ^ c910;
  assign and910 = a910 & b910;
  assign or910  = a910 | b910;
  assign c911 = (a910 & b910) | (a910 & c910) | (b910 & c910);
  wire c_sub911;
  assign c_sub911 = (a910 & b_inv910) | (a910 & c910) | (b_inv910 & c910);
  wire s911, sub911, and911, or911;
  wire b_inv911;
  assign b_inv911 = ~b911;
  assign s911  = a911 ^ b911 ^ c911;
  assign sub911 = a911 ^ b_inv911 ^ c911;
  assign and911 = a911 & b911;
  assign or911  = a911 | b911;
  assign c912 = (a911 & b911) | (a911 & c911) | (b911 & c911);
  wire c_sub912;
  assign c_sub912 = (a911 & b_inv911) | (a911 & c911) | (b_inv911 & c911);
  wire s912, sub912, and912, or912;
  wire b_inv912;
  assign b_inv912 = ~b912;
  assign s912  = a912 ^ b912 ^ c912;
  assign sub912 = a912 ^ b_inv912 ^ c912;
  assign and912 = a912 & b912;
  assign or912  = a912 | b912;
  assign c913 = (a912 & b912) | (a912 & c912) | (b912 & c912);
  wire c_sub913;
  assign c_sub913 = (a912 & b_inv912) | (a912 & c912) | (b_inv912 & c912);
  wire s913, sub913, and913, or913;
  wire b_inv913;
  assign b_inv913 = ~b913;
  assign s913  = a913 ^ b913 ^ c913;
  assign sub913 = a913 ^ b_inv913 ^ c913;
  assign and913 = a913 & b913;
  assign or913  = a913 | b913;
  assign c914 = (a913 & b913) | (a913 & c913) | (b913 & c913);
  wire c_sub914;
  assign c_sub914 = (a913 & b_inv913) | (a913 & c913) | (b_inv913 & c913);
  wire s914, sub914, and914, or914;
  wire b_inv914;
  assign b_inv914 = ~b914;
  assign s914  = a914 ^ b914 ^ c914;
  assign sub914 = a914 ^ b_inv914 ^ c914;
  assign and914 = a914 & b914;
  assign or914  = a914 | b914;
  assign c915 = (a914 & b914) | (a914 & c914) | (b914 & c914);
  wire c_sub915;
  assign c_sub915 = (a914 & b_inv914) | (a914 & c914) | (b_inv914 & c914);
  wire s915, sub915, and915, or915;
  wire b_inv915;
  assign b_inv915 = ~b915;
  assign s915  = a915 ^ b915 ^ c915;
  assign sub915 = a915 ^ b_inv915 ^ c915;
  assign and915 = a915 & b915;
  assign or915  = a915 | b915;
  assign c916 = (a915 & b915) | (a915 & c915) | (b915 & c915);
  wire c_sub916;
  assign c_sub916 = (a915 & b_inv915) | (a915 & c915) | (b_inv915 & c915);
  wire s916, sub916, and916, or916;
  wire b_inv916;
  assign b_inv916 = ~b916;
  assign s916  = a916 ^ b916 ^ c916;
  assign sub916 = a916 ^ b_inv916 ^ c916;
  assign and916 = a916 & b916;
  assign or916  = a916 | b916;
  assign c917 = (a916 & b916) | (a916 & c916) | (b916 & c916);
  wire c_sub917;
  assign c_sub917 = (a916 & b_inv916) | (a916 & c916) | (b_inv916 & c916);
  wire s917, sub917, and917, or917;
  wire b_inv917;
  assign b_inv917 = ~b917;
  assign s917  = a917 ^ b917 ^ c917;
  assign sub917 = a917 ^ b_inv917 ^ c917;
  assign and917 = a917 & b917;
  assign or917  = a917 | b917;
  assign c918 = (a917 & b917) | (a917 & c917) | (b917 & c917);
  wire c_sub918;
  assign c_sub918 = (a917 & b_inv917) | (a917 & c917) | (b_inv917 & c917);
  wire s918, sub918, and918, or918;
  wire b_inv918;
  assign b_inv918 = ~b918;
  assign s918  = a918 ^ b918 ^ c918;
  assign sub918 = a918 ^ b_inv918 ^ c918;
  assign and918 = a918 & b918;
  assign or918  = a918 | b918;
  assign c919 = (a918 & b918) | (a918 & c918) | (b918 & c918);
  wire c_sub919;
  assign c_sub919 = (a918 & b_inv918) | (a918 & c918) | (b_inv918 & c918);
  wire s919, sub919, and919, or919;
  wire b_inv919;
  assign b_inv919 = ~b919;
  assign s919  = a919 ^ b919 ^ c919;
  assign sub919 = a919 ^ b_inv919 ^ c919;
  assign and919 = a919 & b919;
  assign or919  = a919 | b919;
  assign c920 = (a919 & b919) | (a919 & c919) | (b919 & c919);
  wire c_sub920;
  assign c_sub920 = (a919 & b_inv919) | (a919 & c919) | (b_inv919 & c919);
  wire s920, sub920, and920, or920;
  wire b_inv920;
  assign b_inv920 = ~b920;
  assign s920  = a920 ^ b920 ^ c920;
  assign sub920 = a920 ^ b_inv920 ^ c920;
  assign and920 = a920 & b920;
  assign or920  = a920 | b920;
  assign c921 = (a920 & b920) | (a920 & c920) | (b920 & c920);
  wire c_sub921;
  assign c_sub921 = (a920 & b_inv920) | (a920 & c920) | (b_inv920 & c920);
  wire s921, sub921, and921, or921;
  wire b_inv921;
  assign b_inv921 = ~b921;
  assign s921  = a921 ^ b921 ^ c921;
  assign sub921 = a921 ^ b_inv921 ^ c921;
  assign and921 = a921 & b921;
  assign or921  = a921 | b921;
  assign c922 = (a921 & b921) | (a921 & c921) | (b921 & c921);
  wire c_sub922;
  assign c_sub922 = (a921 & b_inv921) | (a921 & c921) | (b_inv921 & c921);
  wire s922, sub922, and922, or922;
  wire b_inv922;
  assign b_inv922 = ~b922;
  assign s922  = a922 ^ b922 ^ c922;
  assign sub922 = a922 ^ b_inv922 ^ c922;
  assign and922 = a922 & b922;
  assign or922  = a922 | b922;
  assign c923 = (a922 & b922) | (a922 & c922) | (b922 & c922);
  wire c_sub923;
  assign c_sub923 = (a922 & b_inv922) | (a922 & c922) | (b_inv922 & c922);
  wire s923, sub923, and923, or923;
  wire b_inv923;
  assign b_inv923 = ~b923;
  assign s923  = a923 ^ b923 ^ c923;
  assign sub923 = a923 ^ b_inv923 ^ c923;
  assign and923 = a923 & b923;
  assign or923  = a923 | b923;
  assign c924 = (a923 & b923) | (a923 & c923) | (b923 & c923);
  wire c_sub924;
  assign c_sub924 = (a923 & b_inv923) | (a923 & c923) | (b_inv923 & c923);
  wire s924, sub924, and924, or924;
  wire b_inv924;
  assign b_inv924 = ~b924;
  assign s924  = a924 ^ b924 ^ c924;
  assign sub924 = a924 ^ b_inv924 ^ c924;
  assign and924 = a924 & b924;
  assign or924  = a924 | b924;
  assign c925 = (a924 & b924) | (a924 & c924) | (b924 & c924);
  wire c_sub925;
  assign c_sub925 = (a924 & b_inv924) | (a924 & c924) | (b_inv924 & c924);
  wire s925, sub925, and925, or925;
  wire b_inv925;
  assign b_inv925 = ~b925;
  assign s925  = a925 ^ b925 ^ c925;
  assign sub925 = a925 ^ b_inv925 ^ c925;
  assign and925 = a925 & b925;
  assign or925  = a925 | b925;
  assign c926 = (a925 & b925) | (a925 & c925) | (b925 & c925);
  wire c_sub926;
  assign c_sub926 = (a925 & b_inv925) | (a925 & c925) | (b_inv925 & c925);
  wire s926, sub926, and926, or926;
  wire b_inv926;
  assign b_inv926 = ~b926;
  assign s926  = a926 ^ b926 ^ c926;
  assign sub926 = a926 ^ b_inv926 ^ c926;
  assign and926 = a926 & b926;
  assign or926  = a926 | b926;
  assign c927 = (a926 & b926) | (a926 & c926) | (b926 & c926);
  wire c_sub927;
  assign c_sub927 = (a926 & b_inv926) | (a926 & c926) | (b_inv926 & c926);
  wire s927, sub927, and927, or927;
  wire b_inv927;
  assign b_inv927 = ~b927;
  assign s927  = a927 ^ b927 ^ c927;
  assign sub927 = a927 ^ b_inv927 ^ c927;
  assign and927 = a927 & b927;
  assign or927  = a927 | b927;
  assign c928 = (a927 & b927) | (a927 & c927) | (b927 & c927);
  wire c_sub928;
  assign c_sub928 = (a927 & b_inv927) | (a927 & c927) | (b_inv927 & c927);
  wire s928, sub928, and928, or928;
  wire b_inv928;
  assign b_inv928 = ~b928;
  assign s928  = a928 ^ b928 ^ c928;
  assign sub928 = a928 ^ b_inv928 ^ c928;
  assign and928 = a928 & b928;
  assign or928  = a928 | b928;
  assign c929 = (a928 & b928) | (a928 & c928) | (b928 & c928);
  wire c_sub929;
  assign c_sub929 = (a928 & b_inv928) | (a928 & c928) | (b_inv928 & c928);
  wire s929, sub929, and929, or929;
  wire b_inv929;
  assign b_inv929 = ~b929;
  assign s929  = a929 ^ b929 ^ c929;
  assign sub929 = a929 ^ b_inv929 ^ c929;
  assign and929 = a929 & b929;
  assign or929  = a929 | b929;
  assign c930 = (a929 & b929) | (a929 & c929) | (b929 & c929);
  wire c_sub930;
  assign c_sub930 = (a929 & b_inv929) | (a929 & c929) | (b_inv929 & c929);
  wire s930, sub930, and930, or930;
  wire b_inv930;
  assign b_inv930 = ~b930;
  assign s930  = a930 ^ b930 ^ c930;
  assign sub930 = a930 ^ b_inv930 ^ c930;
  assign and930 = a930 & b930;
  assign or930  = a930 | b930;
  assign c931 = (a930 & b930) | (a930 & c930) | (b930 & c930);
  wire c_sub931;
  assign c_sub931 = (a930 & b_inv930) | (a930 & c930) | (b_inv930 & c930);
  wire s931, sub931, and931, or931;
  wire b_inv931;
  assign b_inv931 = ~b931;
  assign s931  = a931 ^ b931 ^ c931;
  assign sub931 = a931 ^ b_inv931 ^ c931;
  assign and931 = a931 & b931;
  assign or931  = a931 | b931;
  assign c932 = (a931 & b931) | (a931 & c931) | (b931 & c931);
  wire c_sub932;
  assign c_sub932 = (a931 & b_inv931) | (a931 & c931) | (b_inv931 & c931);
  wire s932, sub932, and932, or932;
  wire b_inv932;
  assign b_inv932 = ~b932;
  assign s932  = a932 ^ b932 ^ c932;
  assign sub932 = a932 ^ b_inv932 ^ c932;
  assign and932 = a932 & b932;
  assign or932  = a932 | b932;
  assign c933 = (a932 & b932) | (a932 & c932) | (b932 & c932);
  wire c_sub933;
  assign c_sub933 = (a932 & b_inv932) | (a932 & c932) | (b_inv932 & c932);
  wire s933, sub933, and933, or933;
  wire b_inv933;
  assign b_inv933 = ~b933;
  assign s933  = a933 ^ b933 ^ c933;
  assign sub933 = a933 ^ b_inv933 ^ c933;
  assign and933 = a933 & b933;
  assign or933  = a933 | b933;
  assign c934 = (a933 & b933) | (a933 & c933) | (b933 & c933);
  wire c_sub934;
  assign c_sub934 = (a933 & b_inv933) | (a933 & c933) | (b_inv933 & c933);
  wire s934, sub934, and934, or934;
  wire b_inv934;
  assign b_inv934 = ~b934;
  assign s934  = a934 ^ b934 ^ c934;
  assign sub934 = a934 ^ b_inv934 ^ c934;
  assign and934 = a934 & b934;
  assign or934  = a934 | b934;
  assign c935 = (a934 & b934) | (a934 & c934) | (b934 & c934);
  wire c_sub935;
  assign c_sub935 = (a934 & b_inv934) | (a934 & c934) | (b_inv934 & c934);
  wire s935, sub935, and935, or935;
  wire b_inv935;
  assign b_inv935 = ~b935;
  assign s935  = a935 ^ b935 ^ c935;
  assign sub935 = a935 ^ b_inv935 ^ c935;
  assign and935 = a935 & b935;
  assign or935  = a935 | b935;
  assign c936 = (a935 & b935) | (a935 & c935) | (b935 & c935);
  wire c_sub936;
  assign c_sub936 = (a935 & b_inv935) | (a935 & c935) | (b_inv935 & c935);
  wire s936, sub936, and936, or936;
  wire b_inv936;
  assign b_inv936 = ~b936;
  assign s936  = a936 ^ b936 ^ c936;
  assign sub936 = a936 ^ b_inv936 ^ c936;
  assign and936 = a936 & b936;
  assign or936  = a936 | b936;
  assign c937 = (a936 & b936) | (a936 & c936) | (b936 & c936);
  wire c_sub937;
  assign c_sub937 = (a936 & b_inv936) | (a936 & c936) | (b_inv936 & c936);
  wire s937, sub937, and937, or937;
  wire b_inv937;
  assign b_inv937 = ~b937;
  assign s937  = a937 ^ b937 ^ c937;
  assign sub937 = a937 ^ b_inv937 ^ c937;
  assign and937 = a937 & b937;
  assign or937  = a937 | b937;
  assign c938 = (a937 & b937) | (a937 & c937) | (b937 & c937);
  wire c_sub938;
  assign c_sub938 = (a937 & b_inv937) | (a937 & c937) | (b_inv937 & c937);
  wire s938, sub938, and938, or938;
  wire b_inv938;
  assign b_inv938 = ~b938;
  assign s938  = a938 ^ b938 ^ c938;
  assign sub938 = a938 ^ b_inv938 ^ c938;
  assign and938 = a938 & b938;
  assign or938  = a938 | b938;
  assign c939 = (a938 & b938) | (a938 & c938) | (b938 & c938);
  wire c_sub939;
  assign c_sub939 = (a938 & b_inv938) | (a938 & c938) | (b_inv938 & c938);
  wire s939, sub939, and939, or939;
  wire b_inv939;
  assign b_inv939 = ~b939;
  assign s939  = a939 ^ b939 ^ c939;
  assign sub939 = a939 ^ b_inv939 ^ c939;
  assign and939 = a939 & b939;
  assign or939  = a939 | b939;
  assign c940 = (a939 & b939) | (a939 & c939) | (b939 & c939);
  wire c_sub940;
  assign c_sub940 = (a939 & b_inv939) | (a939 & c939) | (b_inv939 & c939);
  wire s940, sub940, and940, or940;
  wire b_inv940;
  assign b_inv940 = ~b940;
  assign s940  = a940 ^ b940 ^ c940;
  assign sub940 = a940 ^ b_inv940 ^ c940;
  assign and940 = a940 & b940;
  assign or940  = a940 | b940;
  assign c941 = (a940 & b940) | (a940 & c940) | (b940 & c940);
  wire c_sub941;
  assign c_sub941 = (a940 & b_inv940) | (a940 & c940) | (b_inv940 & c940);
  wire s941, sub941, and941, or941;
  wire b_inv941;
  assign b_inv941 = ~b941;
  assign s941  = a941 ^ b941 ^ c941;
  assign sub941 = a941 ^ b_inv941 ^ c941;
  assign and941 = a941 & b941;
  assign or941  = a941 | b941;
  assign c942 = (a941 & b941) | (a941 & c941) | (b941 & c941);
  wire c_sub942;
  assign c_sub942 = (a941 & b_inv941) | (a941 & c941) | (b_inv941 & c941);
  wire s942, sub942, and942, or942;
  wire b_inv942;
  assign b_inv942 = ~b942;
  assign s942  = a942 ^ b942 ^ c942;
  assign sub942 = a942 ^ b_inv942 ^ c942;
  assign and942 = a942 & b942;
  assign or942  = a942 | b942;
  assign c943 = (a942 & b942) | (a942 & c942) | (b942 & c942);
  wire c_sub943;
  assign c_sub943 = (a942 & b_inv942) | (a942 & c942) | (b_inv942 & c942);
  wire s943, sub943, and943, or943;
  wire b_inv943;
  assign b_inv943 = ~b943;
  assign s943  = a943 ^ b943 ^ c943;
  assign sub943 = a943 ^ b_inv943 ^ c943;
  assign and943 = a943 & b943;
  assign or943  = a943 | b943;
  assign c944 = (a943 & b943) | (a943 & c943) | (b943 & c943);
  wire c_sub944;
  assign c_sub944 = (a943 & b_inv943) | (a943 & c943) | (b_inv943 & c943);
  wire s944, sub944, and944, or944;
  wire b_inv944;
  assign b_inv944 = ~b944;
  assign s944  = a944 ^ b944 ^ c944;
  assign sub944 = a944 ^ b_inv944 ^ c944;
  assign and944 = a944 & b944;
  assign or944  = a944 | b944;
  assign c945 = (a944 & b944) | (a944 & c944) | (b944 & c944);
  wire c_sub945;
  assign c_sub945 = (a944 & b_inv944) | (a944 & c944) | (b_inv944 & c944);
  wire s945, sub945, and945, or945;
  wire b_inv945;
  assign b_inv945 = ~b945;
  assign s945  = a945 ^ b945 ^ c945;
  assign sub945 = a945 ^ b_inv945 ^ c945;
  assign and945 = a945 & b945;
  assign or945  = a945 | b945;
  assign c946 = (a945 & b945) | (a945 & c945) | (b945 & c945);
  wire c_sub946;
  assign c_sub946 = (a945 & b_inv945) | (a945 & c945) | (b_inv945 & c945);
  wire s946, sub946, and946, or946;
  wire b_inv946;
  assign b_inv946 = ~b946;
  assign s946  = a946 ^ b946 ^ c946;
  assign sub946 = a946 ^ b_inv946 ^ c946;
  assign and946 = a946 & b946;
  assign or946  = a946 | b946;
  assign c947 = (a946 & b946) | (a946 & c946) | (b946 & c946);
  wire c_sub947;
  assign c_sub947 = (a946 & b_inv946) | (a946 & c946) | (b_inv946 & c946);
  wire s947, sub947, and947, or947;
  wire b_inv947;
  assign b_inv947 = ~b947;
  assign s947  = a947 ^ b947 ^ c947;
  assign sub947 = a947 ^ b_inv947 ^ c947;
  assign and947 = a947 & b947;
  assign or947  = a947 | b947;
  assign c948 = (a947 & b947) | (a947 & c947) | (b947 & c947);
  wire c_sub948;
  assign c_sub948 = (a947 & b_inv947) | (a947 & c947) | (b_inv947 & c947);
  wire s948, sub948, and948, or948;
  wire b_inv948;
  assign b_inv948 = ~b948;
  assign s948  = a948 ^ b948 ^ c948;
  assign sub948 = a948 ^ b_inv948 ^ c948;
  assign and948 = a948 & b948;
  assign or948  = a948 | b948;
  assign c949 = (a948 & b948) | (a948 & c948) | (b948 & c948);
  wire c_sub949;
  assign c_sub949 = (a948 & b_inv948) | (a948 & c948) | (b_inv948 & c948);
  wire s949, sub949, and949, or949;
  wire b_inv949;
  assign b_inv949 = ~b949;
  assign s949  = a949 ^ b949 ^ c949;
  assign sub949 = a949 ^ b_inv949 ^ c949;
  assign and949 = a949 & b949;
  assign or949  = a949 | b949;
  assign c950 = (a949 & b949) | (a949 & c949) | (b949 & c949);
  wire c_sub950;
  assign c_sub950 = (a949 & b_inv949) | (a949 & c949) | (b_inv949 & c949);
  wire s950, sub950, and950, or950;
  wire b_inv950;
  assign b_inv950 = ~b950;
  assign s950  = a950 ^ b950 ^ c950;
  assign sub950 = a950 ^ b_inv950 ^ c950;
  assign and950 = a950 & b950;
  assign or950  = a950 | b950;
  assign c951 = (a950 & b950) | (a950 & c950) | (b950 & c950);
  wire c_sub951;
  assign c_sub951 = (a950 & b_inv950) | (a950 & c950) | (b_inv950 & c950);
  wire s951, sub951, and951, or951;
  wire b_inv951;
  assign b_inv951 = ~b951;
  assign s951  = a951 ^ b951 ^ c951;
  assign sub951 = a951 ^ b_inv951 ^ c951;
  assign and951 = a951 & b951;
  assign or951  = a951 | b951;
  assign c952 = (a951 & b951) | (a951 & c951) | (b951 & c951);
  wire c_sub952;
  assign c_sub952 = (a951 & b_inv951) | (a951 & c951) | (b_inv951 & c951);
  wire s952, sub952, and952, or952;
  wire b_inv952;
  assign b_inv952 = ~b952;
  assign s952  = a952 ^ b952 ^ c952;
  assign sub952 = a952 ^ b_inv952 ^ c952;
  assign and952 = a952 & b952;
  assign or952  = a952 | b952;
  assign c953 = (a952 & b952) | (a952 & c952) | (b952 & c952);
  wire c_sub953;
  assign c_sub953 = (a952 & b_inv952) | (a952 & c952) | (b_inv952 & c952);
  wire s953, sub953, and953, or953;
  wire b_inv953;
  assign b_inv953 = ~b953;
  assign s953  = a953 ^ b953 ^ c953;
  assign sub953 = a953 ^ b_inv953 ^ c953;
  assign and953 = a953 & b953;
  assign or953  = a953 | b953;
  assign c954 = (a953 & b953) | (a953 & c953) | (b953 & c953);
  wire c_sub954;
  assign c_sub954 = (a953 & b_inv953) | (a953 & c953) | (b_inv953 & c953);
  wire s954, sub954, and954, or954;
  wire b_inv954;
  assign b_inv954 = ~b954;
  assign s954  = a954 ^ b954 ^ c954;
  assign sub954 = a954 ^ b_inv954 ^ c954;
  assign and954 = a954 & b954;
  assign or954  = a954 | b954;
  assign c955 = (a954 & b954) | (a954 & c954) | (b954 & c954);
  wire c_sub955;
  assign c_sub955 = (a954 & b_inv954) | (a954 & c954) | (b_inv954 & c954);
  wire s955, sub955, and955, or955;
  wire b_inv955;
  assign b_inv955 = ~b955;
  assign s955  = a955 ^ b955 ^ c955;
  assign sub955 = a955 ^ b_inv955 ^ c955;
  assign and955 = a955 & b955;
  assign or955  = a955 | b955;
  assign c956 = (a955 & b955) | (a955 & c955) | (b955 & c955);
  wire c_sub956;
  assign c_sub956 = (a955 & b_inv955) | (a955 & c955) | (b_inv955 & c955);
  wire s956, sub956, and956, or956;
  wire b_inv956;
  assign b_inv956 = ~b956;
  assign s956  = a956 ^ b956 ^ c956;
  assign sub956 = a956 ^ b_inv956 ^ c956;
  assign and956 = a956 & b956;
  assign or956  = a956 | b956;
  assign c957 = (a956 & b956) | (a956 & c956) | (b956 & c956);
  wire c_sub957;
  assign c_sub957 = (a956 & b_inv956) | (a956 & c956) | (b_inv956 & c956);
  wire s957, sub957, and957, or957;
  wire b_inv957;
  assign b_inv957 = ~b957;
  assign s957  = a957 ^ b957 ^ c957;
  assign sub957 = a957 ^ b_inv957 ^ c957;
  assign and957 = a957 & b957;
  assign or957  = a957 | b957;
  assign c958 = (a957 & b957) | (a957 & c957) | (b957 & c957);
  wire c_sub958;
  assign c_sub958 = (a957 & b_inv957) | (a957 & c957) | (b_inv957 & c957);
  wire s958, sub958, and958, or958;
  wire b_inv958;
  assign b_inv958 = ~b958;
  assign s958  = a958 ^ b958 ^ c958;
  assign sub958 = a958 ^ b_inv958 ^ c958;
  assign and958 = a958 & b958;
  assign or958  = a958 | b958;
  assign c959 = (a958 & b958) | (a958 & c958) | (b958 & c958);
  wire c_sub959;
  assign c_sub959 = (a958 & b_inv958) | (a958 & c958) | (b_inv958 & c958);
  wire s959, sub959, and959, or959;
  wire b_inv959;
  assign b_inv959 = ~b959;
  assign s959  = a959 ^ b959 ^ c959;
  assign sub959 = a959 ^ b_inv959 ^ c959;
  assign and959 = a959 & b959;
  assign or959  = a959 | b959;
  assign c960 = (a959 & b959) | (a959 & c959) | (b959 & c959);
  wire c_sub960;
  assign c_sub960 = (a959 & b_inv959) | (a959 & c959) | (b_inv959 & c959);
  wire s960, sub960, and960, or960;
  wire b_inv960;
  assign b_inv960 = ~b960;
  assign s960  = a960 ^ b960 ^ c960;
  assign sub960 = a960 ^ b_inv960 ^ c960;
  assign and960 = a960 & b960;
  assign or960  = a960 | b960;
  assign c961 = (a960 & b960) | (a960 & c960) | (b960 & c960);
  wire c_sub961;
  assign c_sub961 = (a960 & b_inv960) | (a960 & c960) | (b_inv960 & c960);
  wire s961, sub961, and961, or961;
  wire b_inv961;
  assign b_inv961 = ~b961;
  assign s961  = a961 ^ b961 ^ c961;
  assign sub961 = a961 ^ b_inv961 ^ c961;
  assign and961 = a961 & b961;
  assign or961  = a961 | b961;
  assign c962 = (a961 & b961) | (a961 & c961) | (b961 & c961);
  wire c_sub962;
  assign c_sub962 = (a961 & b_inv961) | (a961 & c961) | (b_inv961 & c961);
  wire s962, sub962, and962, or962;
  wire b_inv962;
  assign b_inv962 = ~b962;
  assign s962  = a962 ^ b962 ^ c962;
  assign sub962 = a962 ^ b_inv962 ^ c962;
  assign and962 = a962 & b962;
  assign or962  = a962 | b962;
  assign c963 = (a962 & b962) | (a962 & c962) | (b962 & c962);
  wire c_sub963;
  assign c_sub963 = (a962 & b_inv962) | (a962 & c962) | (b_inv962 & c962);
  wire s963, sub963, and963, or963;
  wire b_inv963;
  assign b_inv963 = ~b963;
  assign s963  = a963 ^ b963 ^ c963;
  assign sub963 = a963 ^ b_inv963 ^ c963;
  assign and963 = a963 & b963;
  assign or963  = a963 | b963;
  assign c964 = (a963 & b963) | (a963 & c963) | (b963 & c963);
  wire c_sub964;
  assign c_sub964 = (a963 & b_inv963) | (a963 & c963) | (b_inv963 & c963);
  wire s964, sub964, and964, or964;
  wire b_inv964;
  assign b_inv964 = ~b964;
  assign s964  = a964 ^ b964 ^ c964;
  assign sub964 = a964 ^ b_inv964 ^ c964;
  assign and964 = a964 & b964;
  assign or964  = a964 | b964;
  assign c965 = (a964 & b964) | (a964 & c964) | (b964 & c964);
  wire c_sub965;
  assign c_sub965 = (a964 & b_inv964) | (a964 & c964) | (b_inv964 & c964);
  wire s965, sub965, and965, or965;
  wire b_inv965;
  assign b_inv965 = ~b965;
  assign s965  = a965 ^ b965 ^ c965;
  assign sub965 = a965 ^ b_inv965 ^ c965;
  assign and965 = a965 & b965;
  assign or965  = a965 | b965;
  assign c966 = (a965 & b965) | (a965 & c965) | (b965 & c965);
  wire c_sub966;
  assign c_sub966 = (a965 & b_inv965) | (a965 & c965) | (b_inv965 & c965);
  wire s966, sub966, and966, or966;
  wire b_inv966;
  assign b_inv966 = ~b966;
  assign s966  = a966 ^ b966 ^ c966;
  assign sub966 = a966 ^ b_inv966 ^ c966;
  assign and966 = a966 & b966;
  assign or966  = a966 | b966;
  assign c967 = (a966 & b966) | (a966 & c966) | (b966 & c966);
  wire c_sub967;
  assign c_sub967 = (a966 & b_inv966) | (a966 & c966) | (b_inv966 & c966);
  wire s967, sub967, and967, or967;
  wire b_inv967;
  assign b_inv967 = ~b967;
  assign s967  = a967 ^ b967 ^ c967;
  assign sub967 = a967 ^ b_inv967 ^ c967;
  assign and967 = a967 & b967;
  assign or967  = a967 | b967;
  assign c968 = (a967 & b967) | (a967 & c967) | (b967 & c967);
  wire c_sub968;
  assign c_sub968 = (a967 & b_inv967) | (a967 & c967) | (b_inv967 & c967);
  wire s968, sub968, and968, or968;
  wire b_inv968;
  assign b_inv968 = ~b968;
  assign s968  = a968 ^ b968 ^ c968;
  assign sub968 = a968 ^ b_inv968 ^ c968;
  assign and968 = a968 & b968;
  assign or968  = a968 | b968;
  assign c969 = (a968 & b968) | (a968 & c968) | (b968 & c968);
  wire c_sub969;
  assign c_sub969 = (a968 & b_inv968) | (a968 & c968) | (b_inv968 & c968);
  wire s969, sub969, and969, or969;
  wire b_inv969;
  assign b_inv969 = ~b969;
  assign s969  = a969 ^ b969 ^ c969;
  assign sub969 = a969 ^ b_inv969 ^ c969;
  assign and969 = a969 & b969;
  assign or969  = a969 | b969;
  assign c970 = (a969 & b969) | (a969 & c969) | (b969 & c969);
  wire c_sub970;
  assign c_sub970 = (a969 & b_inv969) | (a969 & c969) | (b_inv969 & c969);
  wire s970, sub970, and970, or970;
  wire b_inv970;
  assign b_inv970 = ~b970;
  assign s970  = a970 ^ b970 ^ c970;
  assign sub970 = a970 ^ b_inv970 ^ c970;
  assign and970 = a970 & b970;
  assign or970  = a970 | b970;
  assign c971 = (a970 & b970) | (a970 & c970) | (b970 & c970);
  wire c_sub971;
  assign c_sub971 = (a970 & b_inv970) | (a970 & c970) | (b_inv970 & c970);
  wire s971, sub971, and971, or971;
  wire b_inv971;
  assign b_inv971 = ~b971;
  assign s971  = a971 ^ b971 ^ c971;
  assign sub971 = a971 ^ b_inv971 ^ c971;
  assign and971 = a971 & b971;
  assign or971  = a971 | b971;
  assign c972 = (a971 & b971) | (a971 & c971) | (b971 & c971);
  wire c_sub972;
  assign c_sub972 = (a971 & b_inv971) | (a971 & c971) | (b_inv971 & c971);
  wire s972, sub972, and972, or972;
  wire b_inv972;
  assign b_inv972 = ~b972;
  assign s972  = a972 ^ b972 ^ c972;
  assign sub972 = a972 ^ b_inv972 ^ c972;
  assign and972 = a972 & b972;
  assign or972  = a972 | b972;
  assign c973 = (a972 & b972) | (a972 & c972) | (b972 & c972);
  wire c_sub973;
  assign c_sub973 = (a972 & b_inv972) | (a972 & c972) | (b_inv972 & c972);
  wire s973, sub973, and973, or973;
  wire b_inv973;
  assign b_inv973 = ~b973;
  assign s973  = a973 ^ b973 ^ c973;
  assign sub973 = a973 ^ b_inv973 ^ c973;
  assign and973 = a973 & b973;
  assign or973  = a973 | b973;
  assign c974 = (a973 & b973) | (a973 & c973) | (b973 & c973);
  wire c_sub974;
  assign c_sub974 = (a973 & b_inv973) | (a973 & c973) | (b_inv973 & c973);
  wire s974, sub974, and974, or974;
  wire b_inv974;
  assign b_inv974 = ~b974;
  assign s974  = a974 ^ b974 ^ c974;
  assign sub974 = a974 ^ b_inv974 ^ c974;
  assign and974 = a974 & b974;
  assign or974  = a974 | b974;
  assign c975 = (a974 & b974) | (a974 & c974) | (b974 & c974);
  wire c_sub975;
  assign c_sub975 = (a974 & b_inv974) | (a974 & c974) | (b_inv974 & c974);
  wire s975, sub975, and975, or975;
  wire b_inv975;
  assign b_inv975 = ~b975;
  assign s975  = a975 ^ b975 ^ c975;
  assign sub975 = a975 ^ b_inv975 ^ c975;
  assign and975 = a975 & b975;
  assign or975  = a975 | b975;
  assign c976 = (a975 & b975) | (a975 & c975) | (b975 & c975);
  wire c_sub976;
  assign c_sub976 = (a975 & b_inv975) | (a975 & c975) | (b_inv975 & c975);
  wire s976, sub976, and976, or976;
  wire b_inv976;
  assign b_inv976 = ~b976;
  assign s976  = a976 ^ b976 ^ c976;
  assign sub976 = a976 ^ b_inv976 ^ c976;
  assign and976 = a976 & b976;
  assign or976  = a976 | b976;
  assign c977 = (a976 & b976) | (a976 & c976) | (b976 & c976);
  wire c_sub977;
  assign c_sub977 = (a976 & b_inv976) | (a976 & c976) | (b_inv976 & c976);
  wire s977, sub977, and977, or977;
  wire b_inv977;
  assign b_inv977 = ~b977;
  assign s977  = a977 ^ b977 ^ c977;
  assign sub977 = a977 ^ b_inv977 ^ c977;
  assign and977 = a977 & b977;
  assign or977  = a977 | b977;
  assign c978 = (a977 & b977) | (a977 & c977) | (b977 & c977);
  wire c_sub978;
  assign c_sub978 = (a977 & b_inv977) | (a977 & c977) | (b_inv977 & c977);
  wire s978, sub978, and978, or978;
  wire b_inv978;
  assign b_inv978 = ~b978;
  assign s978  = a978 ^ b978 ^ c978;
  assign sub978 = a978 ^ b_inv978 ^ c978;
  assign and978 = a978 & b978;
  assign or978  = a978 | b978;
  assign c979 = (a978 & b978) | (a978 & c978) | (b978 & c978);
  wire c_sub979;
  assign c_sub979 = (a978 & b_inv978) | (a978 & c978) | (b_inv978 & c978);
  wire s979, sub979, and979, or979;
  wire b_inv979;
  assign b_inv979 = ~b979;
  assign s979  = a979 ^ b979 ^ c979;
  assign sub979 = a979 ^ b_inv979 ^ c979;
  assign and979 = a979 & b979;
  assign or979  = a979 | b979;
  assign c980 = (a979 & b979) | (a979 & c979) | (b979 & c979);
  wire c_sub980;
  assign c_sub980 = (a979 & b_inv979) | (a979 & c979) | (b_inv979 & c979);
  wire s980, sub980, and980, or980;
  wire b_inv980;
  assign b_inv980 = ~b980;
  assign s980  = a980 ^ b980 ^ c980;
  assign sub980 = a980 ^ b_inv980 ^ c980;
  assign and980 = a980 & b980;
  assign or980  = a980 | b980;
  assign c981 = (a980 & b980) | (a980 & c980) | (b980 & c980);
  wire c_sub981;
  assign c_sub981 = (a980 & b_inv980) | (a980 & c980) | (b_inv980 & c980);
  wire s981, sub981, and981, or981;
  wire b_inv981;
  assign b_inv981 = ~b981;
  assign s981  = a981 ^ b981 ^ c981;
  assign sub981 = a981 ^ b_inv981 ^ c981;
  assign and981 = a981 & b981;
  assign or981  = a981 | b981;
  assign c982 = (a981 & b981) | (a981 & c981) | (b981 & c981);
  wire c_sub982;
  assign c_sub982 = (a981 & b_inv981) | (a981 & c981) | (b_inv981 & c981);
  wire s982, sub982, and982, or982;
  wire b_inv982;
  assign b_inv982 = ~b982;
  assign s982  = a982 ^ b982 ^ c982;
  assign sub982 = a982 ^ b_inv982 ^ c982;
  assign and982 = a982 & b982;
  assign or982  = a982 | b982;
  assign c983 = (a982 & b982) | (a982 & c982) | (b982 & c982);
  wire c_sub983;
  assign c_sub983 = (a982 & b_inv982) | (a982 & c982) | (b_inv982 & c982);
  wire s983, sub983, and983, or983;
  wire b_inv983;
  assign b_inv983 = ~b983;
  assign s983  = a983 ^ b983 ^ c983;
  assign sub983 = a983 ^ b_inv983 ^ c983;
  assign and983 = a983 & b983;
  assign or983  = a983 | b983;
  assign c984 = (a983 & b983) | (a983 & c983) | (b983 & c983);
  wire c_sub984;
  assign c_sub984 = (a983 & b_inv983) | (a983 & c983) | (b_inv983 & c983);
  wire s984, sub984, and984, or984;
  wire b_inv984;
  assign b_inv984 = ~b984;
  assign s984  = a984 ^ b984 ^ c984;
  assign sub984 = a984 ^ b_inv984 ^ c984;
  assign and984 = a984 & b984;
  assign or984  = a984 | b984;
  assign c985 = (a984 & b984) | (a984 & c984) | (b984 & c984);
  wire c_sub985;
  assign c_sub985 = (a984 & b_inv984) | (a984 & c984) | (b_inv984 & c984);
  wire s985, sub985, and985, or985;
  wire b_inv985;
  assign b_inv985 = ~b985;
  assign s985  = a985 ^ b985 ^ c985;
  assign sub985 = a985 ^ b_inv985 ^ c985;
  assign and985 = a985 & b985;
  assign or985  = a985 | b985;
  assign c986 = (a985 & b985) | (a985 & c985) | (b985 & c985);
  wire c_sub986;
  assign c_sub986 = (a985 & b_inv985) | (a985 & c985) | (b_inv985 & c985);
  wire s986, sub986, and986, or986;
  wire b_inv986;
  assign b_inv986 = ~b986;
  assign s986  = a986 ^ b986 ^ c986;
  assign sub986 = a986 ^ b_inv986 ^ c986;
  assign and986 = a986 & b986;
  assign or986  = a986 | b986;
  assign c987 = (a986 & b986) | (a986 & c986) | (b986 & c986);
  wire c_sub987;
  assign c_sub987 = (a986 & b_inv986) | (a986 & c986) | (b_inv986 & c986);
  wire s987, sub987, and987, or987;
  wire b_inv987;
  assign b_inv987 = ~b987;
  assign s987  = a987 ^ b987 ^ c987;
  assign sub987 = a987 ^ b_inv987 ^ c987;
  assign and987 = a987 & b987;
  assign or987  = a987 | b987;
  assign c988 = (a987 & b987) | (a987 & c987) | (b987 & c987);
  wire c_sub988;
  assign c_sub988 = (a987 & b_inv987) | (a987 & c987) | (b_inv987 & c987);
  wire s988, sub988, and988, or988;
  wire b_inv988;
  assign b_inv988 = ~b988;
  assign s988  = a988 ^ b988 ^ c988;
  assign sub988 = a988 ^ b_inv988 ^ c988;
  assign and988 = a988 & b988;
  assign or988  = a988 | b988;
  assign c989 = (a988 & b988) | (a988 & c988) | (b988 & c988);
  wire c_sub989;
  assign c_sub989 = (a988 & b_inv988) | (a988 & c988) | (b_inv988 & c988);
  wire s989, sub989, and989, or989;
  wire b_inv989;
  assign b_inv989 = ~b989;
  assign s989  = a989 ^ b989 ^ c989;
  assign sub989 = a989 ^ b_inv989 ^ c989;
  assign and989 = a989 & b989;
  assign or989  = a989 | b989;
  assign c990 = (a989 & b989) | (a989 & c989) | (b989 & c989);
  wire c_sub990;
  assign c_sub990 = (a989 & b_inv989) | (a989 & c989) | (b_inv989 & c989);
  wire s990, sub990, and990, or990;
  wire b_inv990;
  assign b_inv990 = ~b990;
  assign s990  = a990 ^ b990 ^ c990;
  assign sub990 = a990 ^ b_inv990 ^ c990;
  assign and990 = a990 & b990;
  assign or990  = a990 | b990;
  assign c991 = (a990 & b990) | (a990 & c990) | (b990 & c990);
  wire c_sub991;
  assign c_sub991 = (a990 & b_inv990) | (a990 & c990) | (b_inv990 & c990);
  wire s991, sub991, and991, or991;
  wire b_inv991;
  assign b_inv991 = ~b991;
  assign s991  = a991 ^ b991 ^ c991;
  assign sub991 = a991 ^ b_inv991 ^ c991;
  assign and991 = a991 & b991;
  assign or991  = a991 | b991;
  assign c992 = (a991 & b991) | (a991 & c991) | (b991 & c991);
  wire c_sub992;
  assign c_sub992 = (a991 & b_inv991) | (a991 & c991) | (b_inv991 & c991);
  wire s992, sub992, and992, or992;
  wire b_inv992;
  assign b_inv992 = ~b992;
  assign s992  = a992 ^ b992 ^ c992;
  assign sub992 = a992 ^ b_inv992 ^ c992;
  assign and992 = a992 & b992;
  assign or992  = a992 | b992;
  assign c993 = (a992 & b992) | (a992 & c992) | (b992 & c992);
  wire c_sub993;
  assign c_sub993 = (a992 & b_inv992) | (a992 & c992) | (b_inv992 & c992);
  wire s993, sub993, and993, or993;
  wire b_inv993;
  assign b_inv993 = ~b993;
  assign s993  = a993 ^ b993 ^ c993;
  assign sub993 = a993 ^ b_inv993 ^ c993;
  assign and993 = a993 & b993;
  assign or993  = a993 | b993;
  assign c994 = (a993 & b993) | (a993 & c993) | (b993 & c993);
  wire c_sub994;
  assign c_sub994 = (a993 & b_inv993) | (a993 & c993) | (b_inv993 & c993);
  wire s994, sub994, and994, or994;
  wire b_inv994;
  assign b_inv994 = ~b994;
  assign s994  = a994 ^ b994 ^ c994;
  assign sub994 = a994 ^ b_inv994 ^ c994;
  assign and994 = a994 & b994;
  assign or994  = a994 | b994;
  assign c995 = (a994 & b994) | (a994 & c994) | (b994 & c994);
  wire c_sub995;
  assign c_sub995 = (a994 & b_inv994) | (a994 & c994) | (b_inv994 & c994);
  wire s995, sub995, and995, or995;
  wire b_inv995;
  assign b_inv995 = ~b995;
  assign s995  = a995 ^ b995 ^ c995;
  assign sub995 = a995 ^ b_inv995 ^ c995;
  assign and995 = a995 & b995;
  assign or995  = a995 | b995;
  assign c996 = (a995 & b995) | (a995 & c995) | (b995 & c995);
  wire c_sub996;
  assign c_sub996 = (a995 & b_inv995) | (a995 & c995) | (b_inv995 & c995);
  wire s996, sub996, and996, or996;
  wire b_inv996;
  assign b_inv996 = ~b996;
  assign s996  = a996 ^ b996 ^ c996;
  assign sub996 = a996 ^ b_inv996 ^ c996;
  assign and996 = a996 & b996;
  assign or996  = a996 | b996;
  assign c997 = (a996 & b996) | (a996 & c996) | (b996 & c996);
  wire c_sub997;
  assign c_sub997 = (a996 & b_inv996) | (a996 & c996) | (b_inv996 & c996);
  wire s997, sub997, and997, or997;
  wire b_inv997;
  assign b_inv997 = ~b997;
  assign s997  = a997 ^ b997 ^ c997;
  assign sub997 = a997 ^ b_inv997 ^ c997;
  assign and997 = a997 & b997;
  assign or997  = a997 | b997;
  assign c998 = (a997 & b997) | (a997 & c997) | (b997 & c997);
  wire c_sub998;
  assign c_sub998 = (a997 & b_inv997) | (a997 & c997) | (b_inv997 & c997);
  wire s998, sub998, and998, or998;
  wire b_inv998;
  assign b_inv998 = ~b998;
  assign s998  = a998 ^ b998 ^ c998;
  assign sub998 = a998 ^ b_inv998 ^ c998;
  assign and998 = a998 & b998;
  assign or998  = a998 | b998;
  assign c999 = (a998 & b998) | (a998 & c998) | (b998 & c998);
  wire c_sub999;
  assign c_sub999 = (a998 & b_inv998) | (a998 & c998) | (b_inv998 & c998);
  wire s999, sub999, and999, or999;
  wire b_inv999;
  assign b_inv999 = ~b999;
  assign s999  = a999 ^ b999 ^ c999;
  assign sub999 = a999 ^ b_inv999 ^ c999;
  assign and999 = a999 & b999;
  assign or999  = a999 | b999;
  assign c1000 = (a999 & b999) | (a999 & c999) | (b999 & c999);
  wire c_sub1000;
  assign c_sub1000 = (a999 & b_inv999) | (a999 & c999) | (b_inv999 & c999);
  wire s1000, sub1000, and1000, or1000;
  wire b_inv1000;
  assign b_inv1000 = ~b1000;
  assign s1000  = a1000 ^ b1000 ^ c1000;
  assign sub1000 = a1000 ^ b_inv1000 ^ c1000;
  assign and1000 = a1000 & b1000;
  assign or1000  = a1000 | b1000;
  assign c1001 = (a1000 & b1000) | (a1000 & c1000) | (b1000 & c1000);
  wire c_sub1001;
  assign c_sub1001 = (a1000 & b_inv1000) | (a1000 & c1000) | (b_inv1000 & c1000);
  wire s1001, sub1001, and1001, or1001;
  wire b_inv1001;
  assign b_inv1001 = ~b1001;
  assign s1001  = a1001 ^ b1001 ^ c1001;
  assign sub1001 = a1001 ^ b_inv1001 ^ c1001;
  assign and1001 = a1001 & b1001;
  assign or1001  = a1001 | b1001;
  assign c1002 = (a1001 & b1001) | (a1001 & c1001) | (b1001 & c1001);
  wire c_sub1002;
  assign c_sub1002 = (a1001 & b_inv1001) | (a1001 & c1001) | (b_inv1001 & c1001);
  wire s1002, sub1002, and1002, or1002;
  wire b_inv1002;
  assign b_inv1002 = ~b1002;
  assign s1002  = a1002 ^ b1002 ^ c1002;
  assign sub1002 = a1002 ^ b_inv1002 ^ c1002;
  assign and1002 = a1002 & b1002;
  assign or1002  = a1002 | b1002;
  assign c1003 = (a1002 & b1002) | (a1002 & c1002) | (b1002 & c1002);
  wire c_sub1003;
  assign c_sub1003 = (a1002 & b_inv1002) | (a1002 & c1002) | (b_inv1002 & c1002);
  wire s1003, sub1003, and1003, or1003;
  wire b_inv1003;
  assign b_inv1003 = ~b1003;
  assign s1003  = a1003 ^ b1003 ^ c1003;
  assign sub1003 = a1003 ^ b_inv1003 ^ c1003;
  assign and1003 = a1003 & b1003;
  assign or1003  = a1003 | b1003;
  assign c1004 = (a1003 & b1003) | (a1003 & c1003) | (b1003 & c1003);
  wire c_sub1004;
  assign c_sub1004 = (a1003 & b_inv1003) | (a1003 & c1003) | (b_inv1003 & c1003);
  wire s1004, sub1004, and1004, or1004;
  wire b_inv1004;
  assign b_inv1004 = ~b1004;
  assign s1004  = a1004 ^ b1004 ^ c1004;
  assign sub1004 = a1004 ^ b_inv1004 ^ c1004;
  assign and1004 = a1004 & b1004;
  assign or1004  = a1004 | b1004;
  assign c1005 = (a1004 & b1004) | (a1004 & c1004) | (b1004 & c1004);
  wire c_sub1005;
  assign c_sub1005 = (a1004 & b_inv1004) | (a1004 & c1004) | (b_inv1004 & c1004);
  wire s1005, sub1005, and1005, or1005;
  wire b_inv1005;
  assign b_inv1005 = ~b1005;
  assign s1005  = a1005 ^ b1005 ^ c1005;
  assign sub1005 = a1005 ^ b_inv1005 ^ c1005;
  assign and1005 = a1005 & b1005;
  assign or1005  = a1005 | b1005;
  assign c1006 = (a1005 & b1005) | (a1005 & c1005) | (b1005 & c1005);
  wire c_sub1006;
  assign c_sub1006 = (a1005 & b_inv1005) | (a1005 & c1005) | (b_inv1005 & c1005);
  wire s1006, sub1006, and1006, or1006;
  wire b_inv1006;
  assign b_inv1006 = ~b1006;
  assign s1006  = a1006 ^ b1006 ^ c1006;
  assign sub1006 = a1006 ^ b_inv1006 ^ c1006;
  assign and1006 = a1006 & b1006;
  assign or1006  = a1006 | b1006;
  assign c1007 = (a1006 & b1006) | (a1006 & c1006) | (b1006 & c1006);
  wire c_sub1007;
  assign c_sub1007 = (a1006 & b_inv1006) | (a1006 & c1006) | (b_inv1006 & c1006);
  wire s1007, sub1007, and1007, or1007;
  wire b_inv1007;
  assign b_inv1007 = ~b1007;
  assign s1007  = a1007 ^ b1007 ^ c1007;
  assign sub1007 = a1007 ^ b_inv1007 ^ c1007;
  assign and1007 = a1007 & b1007;
  assign or1007  = a1007 | b1007;
  assign c1008 = (a1007 & b1007) | (a1007 & c1007) | (b1007 & c1007);
  wire c_sub1008;
  assign c_sub1008 = (a1007 & b_inv1007) | (a1007 & c1007) | (b_inv1007 & c1007);
  wire s1008, sub1008, and1008, or1008;
  wire b_inv1008;
  assign b_inv1008 = ~b1008;
  assign s1008  = a1008 ^ b1008 ^ c1008;
  assign sub1008 = a1008 ^ b_inv1008 ^ c1008;
  assign and1008 = a1008 & b1008;
  assign or1008  = a1008 | b1008;
  assign c1009 = (a1008 & b1008) | (a1008 & c1008) | (b1008 & c1008);
  wire c_sub1009;
  assign c_sub1009 = (a1008 & b_inv1008) | (a1008 & c1008) | (b_inv1008 & c1008);
  wire s1009, sub1009, and1009, or1009;
  wire b_inv1009;
  assign b_inv1009 = ~b1009;
  assign s1009  = a1009 ^ b1009 ^ c1009;
  assign sub1009 = a1009 ^ b_inv1009 ^ c1009;
  assign and1009 = a1009 & b1009;
  assign or1009  = a1009 | b1009;
  assign c1010 = (a1009 & b1009) | (a1009 & c1009) | (b1009 & c1009);
  wire c_sub1010;
  assign c_sub1010 = (a1009 & b_inv1009) | (a1009 & c1009) | (b_inv1009 & c1009);
  wire s1010, sub1010, and1010, or1010;
  wire b_inv1010;
  assign b_inv1010 = ~b1010;
  assign s1010  = a1010 ^ b1010 ^ c1010;
  assign sub1010 = a1010 ^ b_inv1010 ^ c1010;
  assign and1010 = a1010 & b1010;
  assign or1010  = a1010 | b1010;
  assign c1011 = (a1010 & b1010) | (a1010 & c1010) | (b1010 & c1010);
  wire c_sub1011;
  assign c_sub1011 = (a1010 & b_inv1010) | (a1010 & c1010) | (b_inv1010 & c1010);
  wire s1011, sub1011, and1011, or1011;
  wire b_inv1011;
  assign b_inv1011 = ~b1011;
  assign s1011  = a1011 ^ b1011 ^ c1011;
  assign sub1011 = a1011 ^ b_inv1011 ^ c1011;
  assign and1011 = a1011 & b1011;
  assign or1011  = a1011 | b1011;
  assign c1012 = (a1011 & b1011) | (a1011 & c1011) | (b1011 & c1011);
  wire c_sub1012;
  assign c_sub1012 = (a1011 & b_inv1011) | (a1011 & c1011) | (b_inv1011 & c1011);
  wire s1012, sub1012, and1012, or1012;
  wire b_inv1012;
  assign b_inv1012 = ~b1012;
  assign s1012  = a1012 ^ b1012 ^ c1012;
  assign sub1012 = a1012 ^ b_inv1012 ^ c1012;
  assign and1012 = a1012 & b1012;
  assign or1012  = a1012 | b1012;
  assign c1013 = (a1012 & b1012) | (a1012 & c1012) | (b1012 & c1012);
  wire c_sub1013;
  assign c_sub1013 = (a1012 & b_inv1012) | (a1012 & c1012) | (b_inv1012 & c1012);
  wire s1013, sub1013, and1013, or1013;
  wire b_inv1013;
  assign b_inv1013 = ~b1013;
  assign s1013  = a1013 ^ b1013 ^ c1013;
  assign sub1013 = a1013 ^ b_inv1013 ^ c1013;
  assign and1013 = a1013 & b1013;
  assign or1013  = a1013 | b1013;
  assign c1014 = (a1013 & b1013) | (a1013 & c1013) | (b1013 & c1013);
  wire c_sub1014;
  assign c_sub1014 = (a1013 & b_inv1013) | (a1013 & c1013) | (b_inv1013 & c1013);
  wire s1014, sub1014, and1014, or1014;
  wire b_inv1014;
  assign b_inv1014 = ~b1014;
  assign s1014  = a1014 ^ b1014 ^ c1014;
  assign sub1014 = a1014 ^ b_inv1014 ^ c1014;
  assign and1014 = a1014 & b1014;
  assign or1014  = a1014 | b1014;
  assign c1015 = (a1014 & b1014) | (a1014 & c1014) | (b1014 & c1014);
  wire c_sub1015;
  assign c_sub1015 = (a1014 & b_inv1014) | (a1014 & c1014) | (b_inv1014 & c1014);
  wire s1015, sub1015, and1015, or1015;
  wire b_inv1015;
  assign b_inv1015 = ~b1015;
  assign s1015  = a1015 ^ b1015 ^ c1015;
  assign sub1015 = a1015 ^ b_inv1015 ^ c1015;
  assign and1015 = a1015 & b1015;
  assign or1015  = a1015 | b1015;
  assign c1016 = (a1015 & b1015) | (a1015 & c1015) | (b1015 & c1015);
  wire c_sub1016;
  assign c_sub1016 = (a1015 & b_inv1015) | (a1015 & c1015) | (b_inv1015 & c1015);
  wire s1016, sub1016, and1016, or1016;
  wire b_inv1016;
  assign b_inv1016 = ~b1016;
  assign s1016  = a1016 ^ b1016 ^ c1016;
  assign sub1016 = a1016 ^ b_inv1016 ^ c1016;
  assign and1016 = a1016 & b1016;
  assign or1016  = a1016 | b1016;
  assign c1017 = (a1016 & b1016) | (a1016 & c1016) | (b1016 & c1016);
  wire c_sub1017;
  assign c_sub1017 = (a1016 & b_inv1016) | (a1016 & c1016) | (b_inv1016 & c1016);
  wire s1017, sub1017, and1017, or1017;
  wire b_inv1017;
  assign b_inv1017 = ~b1017;
  assign s1017  = a1017 ^ b1017 ^ c1017;
  assign sub1017 = a1017 ^ b_inv1017 ^ c1017;
  assign and1017 = a1017 & b1017;
  assign or1017  = a1017 | b1017;
  assign c1018 = (a1017 & b1017) | (a1017 & c1017) | (b1017 & c1017);
  wire c_sub1018;
  assign c_sub1018 = (a1017 & b_inv1017) | (a1017 & c1017) | (b_inv1017 & c1017);
  wire s1018, sub1018, and1018, or1018;
  wire b_inv1018;
  assign b_inv1018 = ~b1018;
  assign s1018  = a1018 ^ b1018 ^ c1018;
  assign sub1018 = a1018 ^ b_inv1018 ^ c1018;
  assign and1018 = a1018 & b1018;
  assign or1018  = a1018 | b1018;
  assign c1019 = (a1018 & b1018) | (a1018 & c1018) | (b1018 & c1018);
  wire c_sub1019;
  assign c_sub1019 = (a1018 & b_inv1018) | (a1018 & c1018) | (b_inv1018 & c1018);
  wire s1019, sub1019, and1019, or1019;
  wire b_inv1019;
  assign b_inv1019 = ~b1019;
  assign s1019  = a1019 ^ b1019 ^ c1019;
  assign sub1019 = a1019 ^ b_inv1019 ^ c1019;
  assign and1019 = a1019 & b1019;
  assign or1019  = a1019 | b1019;
  assign c1020 = (a1019 & b1019) | (a1019 & c1019) | (b1019 & c1019);
  wire c_sub1020;
  assign c_sub1020 = (a1019 & b_inv1019) | (a1019 & c1019) | (b_inv1019 & c1019);
  wire s1020, sub1020, and1020, or1020;
  wire b_inv1020;
  assign b_inv1020 = ~b1020;
  assign s1020  = a1020 ^ b1020 ^ c1020;
  assign sub1020 = a1020 ^ b_inv1020 ^ c1020;
  assign and1020 = a1020 & b1020;
  assign or1020  = a1020 | b1020;
  assign c1021 = (a1020 & b1020) | (a1020 & c1020) | (b1020 & c1020);
  wire c_sub1021;
  assign c_sub1021 = (a1020 & b_inv1020) | (a1020 & c1020) | (b_inv1020 & c1020);
  wire s1021, sub1021, and1021, or1021;
  wire b_inv1021;
  assign b_inv1021 = ~b1021;
  assign s1021  = a1021 ^ b1021 ^ c1021;
  assign sub1021 = a1021 ^ b_inv1021 ^ c1021;
  assign and1021 = a1021 & b1021;
  assign or1021  = a1021 | b1021;
  assign c1022 = (a1021 & b1021) | (a1021 & c1021) | (b1021 & c1021);
  wire c_sub1022;
  assign c_sub1022 = (a1021 & b_inv1021) | (a1021 & c1021) | (b_inv1021 & c1021);
  wire s1022, sub1022, and1022, or1022;
  wire b_inv1022;
  assign b_inv1022 = ~b1022;
  assign s1022  = a1022 ^ b1022 ^ c1022;
  assign sub1022 = a1022 ^ b_inv1022 ^ c1022;
  assign and1022 = a1022 & b1022;
  assign or1022  = a1022 | b1022;
  assign c1023 = (a1022 & b1022) | (a1022 & c1022) | (b1022 & c1022);
  wire c_sub1023;
  assign c_sub1023 = (a1022 & b_inv1022) | (a1022 & c1022) | (b_inv1022 & c1022);
  wire s1023, sub1023, and1023, or1023;
  wire b_inv1023;
  assign b_inv1023 = ~b1023;
  assign s1023  = a1023 ^ b1023 ^ c1023;
  assign sub1023 = a1023 ^ b_inv1023 ^ c1023;
  assign and1023 = a1023 & b1023;
  assign or1023  = a1023 | b1023;
  assign c1024 = (a1023 & b1023) | (a1023 & c1023) | (b1023 & c1023);
  wire c_sub1024;
  assign c_sub1024 = (a1023 & b_inv1023) | (a1023 & c1023) | (b_inv1023 & c1023);
  assign y0 = (add_sel & s0) | (sub_sel & sub0) | (and_sel & and0) | (or_sel & or0);
  assign y1 = (add_sel & s1) | (sub_sel & sub1) | (and_sel & and1) | (or_sel & or1);
  assign y2 = (add_sel & s2) | (sub_sel & sub2) | (and_sel & and2) | (or_sel & or2);
  assign y3 = (add_sel & s3) | (sub_sel & sub3) | (and_sel & and3) | (or_sel & or3);
  assign y4 = (add_sel & s4) | (sub_sel & sub4) | (and_sel & and4) | (or_sel & or4);
  assign y5 = (add_sel & s5) | (sub_sel & sub5) | (and_sel & and5) | (or_sel & or5);
  assign y6 = (add_sel & s6) | (sub_sel & sub6) | (and_sel & and6) | (or_sel & or6);
  assign y7 = (add_sel & s7) | (sub_sel & sub7) | (and_sel & and7) | (or_sel & or7);
  assign y8 = (add_sel & s8) | (sub_sel & sub8) | (and_sel & and8) | (or_sel & or8);
  assign y9 = (add_sel & s9) | (sub_sel & sub9) | (and_sel & and9) | (or_sel & or9);
  assign y10 = (add_sel & s10) | (sub_sel & sub10) | (and_sel & and10) | (or_sel & or10);
  assign y11 = (add_sel & s11) | (sub_sel & sub11) | (and_sel & and11) | (or_sel & or11);
  assign y12 = (add_sel & s12) | (sub_sel & sub12) | (and_sel & and12) | (or_sel & or12);
  assign y13 = (add_sel & s13) | (sub_sel & sub13) | (and_sel & and13) | (or_sel & or13);
  assign y14 = (add_sel & s14) | (sub_sel & sub14) | (and_sel & and14) | (or_sel & or14);
  assign y15 = (add_sel & s15) | (sub_sel & sub15) | (and_sel & and15) | (or_sel & or15);
  assign y16 = (add_sel & s16) | (sub_sel & sub16) | (and_sel & and16) | (or_sel & or16);
  assign y17 = (add_sel & s17) | (sub_sel & sub17) | (and_sel & and17) | (or_sel & or17);
  assign y18 = (add_sel & s18) | (sub_sel & sub18) | (and_sel & and18) | (or_sel & or18);
  assign y19 = (add_sel & s19) | (sub_sel & sub19) | (and_sel & and19) | (or_sel & or19);
  assign y20 = (add_sel & s20) | (sub_sel & sub20) | (and_sel & and20) | (or_sel & or20);
  assign y21 = (add_sel & s21) | (sub_sel & sub21) | (and_sel & and21) | (or_sel & or21);
  assign y22 = (add_sel & s22) | (sub_sel & sub22) | (and_sel & and22) | (or_sel & or22);
  assign y23 = (add_sel & s23) | (sub_sel & sub23) | (and_sel & and23) | (or_sel & or23);
  assign y24 = (add_sel & s24) | (sub_sel & sub24) | (and_sel & and24) | (or_sel & or24);
  assign y25 = (add_sel & s25) | (sub_sel & sub25) | (and_sel & and25) | (or_sel & or25);
  assign y26 = (add_sel & s26) | (sub_sel & sub26) | (and_sel & and26) | (or_sel & or26);
  assign y27 = (add_sel & s27) | (sub_sel & sub27) | (and_sel & and27) | (or_sel & or27);
  assign y28 = (add_sel & s28) | (sub_sel & sub28) | (and_sel & and28) | (or_sel & or28);
  assign y29 = (add_sel & s29) | (sub_sel & sub29) | (and_sel & and29) | (or_sel & or29);
  assign y30 = (add_sel & s30) | (sub_sel & sub30) | (and_sel & and30) | (or_sel & or30);
  assign y31 = (add_sel & s31) | (sub_sel & sub31) | (and_sel & and31) | (or_sel & or31);
  assign y32 = (add_sel & s32) | (sub_sel & sub32) | (and_sel & and32) | (or_sel & or32);
  assign y33 = (add_sel & s33) | (sub_sel & sub33) | (and_sel & and33) | (or_sel & or33);
  assign y34 = (add_sel & s34) | (sub_sel & sub34) | (and_sel & and34) | (or_sel & or34);
  assign y35 = (add_sel & s35) | (sub_sel & sub35) | (and_sel & and35) | (or_sel & or35);
  assign y36 = (add_sel & s36) | (sub_sel & sub36) | (and_sel & and36) | (or_sel & or36);
  assign y37 = (add_sel & s37) | (sub_sel & sub37) | (and_sel & and37) | (or_sel & or37);
  assign y38 = (add_sel & s38) | (sub_sel & sub38) | (and_sel & and38) | (or_sel & or38);
  assign y39 = (add_sel & s39) | (sub_sel & sub39) | (and_sel & and39) | (or_sel & or39);
  assign y40 = (add_sel & s40) | (sub_sel & sub40) | (and_sel & and40) | (or_sel & or40);
  assign y41 = (add_sel & s41) | (sub_sel & sub41) | (and_sel & and41) | (or_sel & or41);
  assign y42 = (add_sel & s42) | (sub_sel & sub42) | (and_sel & and42) | (or_sel & or42);
  assign y43 = (add_sel & s43) | (sub_sel & sub43) | (and_sel & and43) | (or_sel & or43);
  assign y44 = (add_sel & s44) | (sub_sel & sub44) | (and_sel & and44) | (or_sel & or44);
  assign y45 = (add_sel & s45) | (sub_sel & sub45) | (and_sel & and45) | (or_sel & or45);
  assign y46 = (add_sel & s46) | (sub_sel & sub46) | (and_sel & and46) | (or_sel & or46);
  assign y47 = (add_sel & s47) | (sub_sel & sub47) | (and_sel & and47) | (or_sel & or47);
  assign y48 = (add_sel & s48) | (sub_sel & sub48) | (and_sel & and48) | (or_sel & or48);
  assign y49 = (add_sel & s49) | (sub_sel & sub49) | (and_sel & and49) | (or_sel & or49);
  assign y50 = (add_sel & s50) | (sub_sel & sub50) | (and_sel & and50) | (or_sel & or50);
  assign y51 = (add_sel & s51) | (sub_sel & sub51) | (and_sel & and51) | (or_sel & or51);
  assign y52 = (add_sel & s52) | (sub_sel & sub52) | (and_sel & and52) | (or_sel & or52);
  assign y53 = (add_sel & s53) | (sub_sel & sub53) | (and_sel & and53) | (or_sel & or53);
  assign y54 = (add_sel & s54) | (sub_sel & sub54) | (and_sel & and54) | (or_sel & or54);
  assign y55 = (add_sel & s55) | (sub_sel & sub55) | (and_sel & and55) | (or_sel & or55);
  assign y56 = (add_sel & s56) | (sub_sel & sub56) | (and_sel & and56) | (or_sel & or56);
  assign y57 = (add_sel & s57) | (sub_sel & sub57) | (and_sel & and57) | (or_sel & or57);
  assign y58 = (add_sel & s58) | (sub_sel & sub58) | (and_sel & and58) | (or_sel & or58);
  assign y59 = (add_sel & s59) | (sub_sel & sub59) | (and_sel & and59) | (or_sel & or59);
  assign y60 = (add_sel & s60) | (sub_sel & sub60) | (and_sel & and60) | (or_sel & or60);
  assign y61 = (add_sel & s61) | (sub_sel & sub61) | (and_sel & and61) | (or_sel & or61);
  assign y62 = (add_sel & s62) | (sub_sel & sub62) | (and_sel & and62) | (or_sel & or62);
  assign y63 = (add_sel & s63) | (sub_sel & sub63) | (and_sel & and63) | (or_sel & or63);
  assign y64 = (add_sel & s64) | (sub_sel & sub64) | (and_sel & and64) | (or_sel & or64);
  assign y65 = (add_sel & s65) | (sub_sel & sub65) | (and_sel & and65) | (or_sel & or65);
  assign y66 = (add_sel & s66) | (sub_sel & sub66) | (and_sel & and66) | (or_sel & or66);
  assign y67 = (add_sel & s67) | (sub_sel & sub67) | (and_sel & and67) | (or_sel & or67);
  assign y68 = (add_sel & s68) | (sub_sel & sub68) | (and_sel & and68) | (or_sel & or68);
  assign y69 = (add_sel & s69) | (sub_sel & sub69) | (and_sel & and69) | (or_sel & or69);
  assign y70 = (add_sel & s70) | (sub_sel & sub70) | (and_sel & and70) | (or_sel & or70);
  assign y71 = (add_sel & s71) | (sub_sel & sub71) | (and_sel & and71) | (or_sel & or71);
  assign y72 = (add_sel & s72) | (sub_sel & sub72) | (and_sel & and72) | (or_sel & or72);
  assign y73 = (add_sel & s73) | (sub_sel & sub73) | (and_sel & and73) | (or_sel & or73);
  assign y74 = (add_sel & s74) | (sub_sel & sub74) | (and_sel & and74) | (or_sel & or74);
  assign y75 = (add_sel & s75) | (sub_sel & sub75) | (and_sel & and75) | (or_sel & or75);
  assign y76 = (add_sel & s76) | (sub_sel & sub76) | (and_sel & and76) | (or_sel & or76);
  assign y77 = (add_sel & s77) | (sub_sel & sub77) | (and_sel & and77) | (or_sel & or77);
  assign y78 = (add_sel & s78) | (sub_sel & sub78) | (and_sel & and78) | (or_sel & or78);
  assign y79 = (add_sel & s79) | (sub_sel & sub79) | (and_sel & and79) | (or_sel & or79);
  assign y80 = (add_sel & s80) | (sub_sel & sub80) | (and_sel & and80) | (or_sel & or80);
  assign y81 = (add_sel & s81) | (sub_sel & sub81) | (and_sel & and81) | (or_sel & or81);
  assign y82 = (add_sel & s82) | (sub_sel & sub82) | (and_sel & and82) | (or_sel & or82);
  assign y83 = (add_sel & s83) | (sub_sel & sub83) | (and_sel & and83) | (or_sel & or83);
  assign y84 = (add_sel & s84) | (sub_sel & sub84) | (and_sel & and84) | (or_sel & or84);
  assign y85 = (add_sel & s85) | (sub_sel & sub85) | (and_sel & and85) | (or_sel & or85);
  assign y86 = (add_sel & s86) | (sub_sel & sub86) | (and_sel & and86) | (or_sel & or86);
  assign y87 = (add_sel & s87) | (sub_sel & sub87) | (and_sel & and87) | (or_sel & or87);
  assign y88 = (add_sel & s88) | (sub_sel & sub88) | (and_sel & and88) | (or_sel & or88);
  assign y89 = (add_sel & s89) | (sub_sel & sub89) | (and_sel & and89) | (or_sel & or89);
  assign y90 = (add_sel & s90) | (sub_sel & sub90) | (and_sel & and90) | (or_sel & or90);
  assign y91 = (add_sel & s91) | (sub_sel & sub91) | (and_sel & and91) | (or_sel & or91);
  assign y92 = (add_sel & s92) | (sub_sel & sub92) | (and_sel & and92) | (or_sel & or92);
  assign y93 = (add_sel & s93) | (sub_sel & sub93) | (and_sel & and93) | (or_sel & or93);
  assign y94 = (add_sel & s94) | (sub_sel & sub94) | (and_sel & and94) | (or_sel & or94);
  assign y95 = (add_sel & s95) | (sub_sel & sub95) | (and_sel & and95) | (or_sel & or95);
  assign y96 = (add_sel & s96) | (sub_sel & sub96) | (and_sel & and96) | (or_sel & or96);
  assign y97 = (add_sel & s97) | (sub_sel & sub97) | (and_sel & and97) | (or_sel & or97);
  assign y98 = (add_sel & s98) | (sub_sel & sub98) | (and_sel & and98) | (or_sel & or98);
  assign y99 = (add_sel & s99) | (sub_sel & sub99) | (and_sel & and99) | (or_sel & or99);
  assign y100 = (add_sel & s100) | (sub_sel & sub100) | (and_sel & and100) | (or_sel & or100);
  assign y101 = (add_sel & s101) | (sub_sel & sub101) | (and_sel & and101) | (or_sel & or101);
  assign y102 = (add_sel & s102) | (sub_sel & sub102) | (and_sel & and102) | (or_sel & or102);
  assign y103 = (add_sel & s103) | (sub_sel & sub103) | (and_sel & and103) | (or_sel & or103);
  assign y104 = (add_sel & s104) | (sub_sel & sub104) | (and_sel & and104) | (or_sel & or104);
  assign y105 = (add_sel & s105) | (sub_sel & sub105) | (and_sel & and105) | (or_sel & or105);
  assign y106 = (add_sel & s106) | (sub_sel & sub106) | (and_sel & and106) | (or_sel & or106);
  assign y107 = (add_sel & s107) | (sub_sel & sub107) | (and_sel & and107) | (or_sel & or107);
  assign y108 = (add_sel & s108) | (sub_sel & sub108) | (and_sel & and108) | (or_sel & or108);
  assign y109 = (add_sel & s109) | (sub_sel & sub109) | (and_sel & and109) | (or_sel & or109);
  assign y110 = (add_sel & s110) | (sub_sel & sub110) | (and_sel & and110) | (or_sel & or110);
  assign y111 = (add_sel & s111) | (sub_sel & sub111) | (and_sel & and111) | (or_sel & or111);
  assign y112 = (add_sel & s112) | (sub_sel & sub112) | (and_sel & and112) | (or_sel & or112);
  assign y113 = (add_sel & s113) | (sub_sel & sub113) | (and_sel & and113) | (or_sel & or113);
  assign y114 = (add_sel & s114) | (sub_sel & sub114) | (and_sel & and114) | (or_sel & or114);
  assign y115 = (add_sel & s115) | (sub_sel & sub115) | (and_sel & and115) | (or_sel & or115);
  assign y116 = (add_sel & s116) | (sub_sel & sub116) | (and_sel & and116) | (or_sel & or116);
  assign y117 = (add_sel & s117) | (sub_sel & sub117) | (and_sel & and117) | (or_sel & or117);
  assign y118 = (add_sel & s118) | (sub_sel & sub118) | (and_sel & and118) | (or_sel & or118);
  assign y119 = (add_sel & s119) | (sub_sel & sub119) | (and_sel & and119) | (or_sel & or119);
  assign y120 = (add_sel & s120) | (sub_sel & sub120) | (and_sel & and120) | (or_sel & or120);
  assign y121 = (add_sel & s121) | (sub_sel & sub121) | (and_sel & and121) | (or_sel & or121);
  assign y122 = (add_sel & s122) | (sub_sel & sub122) | (and_sel & and122) | (or_sel & or122);
  assign y123 = (add_sel & s123) | (sub_sel & sub123) | (and_sel & and123) | (or_sel & or123);
  assign y124 = (add_sel & s124) | (sub_sel & sub124) | (and_sel & and124) | (or_sel & or124);
  assign y125 = (add_sel & s125) | (sub_sel & sub125) | (and_sel & and125) | (or_sel & or125);
  assign y126 = (add_sel & s126) | (sub_sel & sub126) | (and_sel & and126) | (or_sel & or126);
  assign y127 = (add_sel & s127) | (sub_sel & sub127) | (and_sel & and127) | (or_sel & or127);
  assign y128 = (add_sel & s128) | (sub_sel & sub128) | (and_sel & and128) | (or_sel & or128);
  assign y129 = (add_sel & s129) | (sub_sel & sub129) | (and_sel & and129) | (or_sel & or129);
  assign y130 = (add_sel & s130) | (sub_sel & sub130) | (and_sel & and130) | (or_sel & or130);
  assign y131 = (add_sel & s131) | (sub_sel & sub131) | (and_sel & and131) | (or_sel & or131);
  assign y132 = (add_sel & s132) | (sub_sel & sub132) | (and_sel & and132) | (or_sel & or132);
  assign y133 = (add_sel & s133) | (sub_sel & sub133) | (and_sel & and133) | (or_sel & or133);
  assign y134 = (add_sel & s134) | (sub_sel & sub134) | (and_sel & and134) | (or_sel & or134);
  assign y135 = (add_sel & s135) | (sub_sel & sub135) | (and_sel & and135) | (or_sel & or135);
  assign y136 = (add_sel & s136) | (sub_sel & sub136) | (and_sel & and136) | (or_sel & or136);
  assign y137 = (add_sel & s137) | (sub_sel & sub137) | (and_sel & and137) | (or_sel & or137);
  assign y138 = (add_sel & s138) | (sub_sel & sub138) | (and_sel & and138) | (or_sel & or138);
  assign y139 = (add_sel & s139) | (sub_sel & sub139) | (and_sel & and139) | (or_sel & or139);
  assign y140 = (add_sel & s140) | (sub_sel & sub140) | (and_sel & and140) | (or_sel & or140);
  assign y141 = (add_sel & s141) | (sub_sel & sub141) | (and_sel & and141) | (or_sel & or141);
  assign y142 = (add_sel & s142) | (sub_sel & sub142) | (and_sel & and142) | (or_sel & or142);
  assign y143 = (add_sel & s143) | (sub_sel & sub143) | (and_sel & and143) | (or_sel & or143);
  assign y144 = (add_sel & s144) | (sub_sel & sub144) | (and_sel & and144) | (or_sel & or144);
  assign y145 = (add_sel & s145) | (sub_sel & sub145) | (and_sel & and145) | (or_sel & or145);
  assign y146 = (add_sel & s146) | (sub_sel & sub146) | (and_sel & and146) | (or_sel & or146);
  assign y147 = (add_sel & s147) | (sub_sel & sub147) | (and_sel & and147) | (or_sel & or147);
  assign y148 = (add_sel & s148) | (sub_sel & sub148) | (and_sel & and148) | (or_sel & or148);
  assign y149 = (add_sel & s149) | (sub_sel & sub149) | (and_sel & and149) | (or_sel & or149);
  assign y150 = (add_sel & s150) | (sub_sel & sub150) | (and_sel & and150) | (or_sel & or150);
  assign y151 = (add_sel & s151) | (sub_sel & sub151) | (and_sel & and151) | (or_sel & or151);
  assign y152 = (add_sel & s152) | (sub_sel & sub152) | (and_sel & and152) | (or_sel & or152);
  assign y153 = (add_sel & s153) | (sub_sel & sub153) | (and_sel & and153) | (or_sel & or153);
  assign y154 = (add_sel & s154) | (sub_sel & sub154) | (and_sel & and154) | (or_sel & or154);
  assign y155 = (add_sel & s155) | (sub_sel & sub155) | (and_sel & and155) | (or_sel & or155);
  assign y156 = (add_sel & s156) | (sub_sel & sub156) | (and_sel & and156) | (or_sel & or156);
  assign y157 = (add_sel & s157) | (sub_sel & sub157) | (and_sel & and157) | (or_sel & or157);
  assign y158 = (add_sel & s158) | (sub_sel & sub158) | (and_sel & and158) | (or_sel & or158);
  assign y159 = (add_sel & s159) | (sub_sel & sub159) | (and_sel & and159) | (or_sel & or159);
  assign y160 = (add_sel & s160) | (sub_sel & sub160) | (and_sel & and160) | (or_sel & or160);
  assign y161 = (add_sel & s161) | (sub_sel & sub161) | (and_sel & and161) | (or_sel & or161);
  assign y162 = (add_sel & s162) | (sub_sel & sub162) | (and_sel & and162) | (or_sel & or162);
  assign y163 = (add_sel & s163) | (sub_sel & sub163) | (and_sel & and163) | (or_sel & or163);
  assign y164 = (add_sel & s164) | (sub_sel & sub164) | (and_sel & and164) | (or_sel & or164);
  assign y165 = (add_sel & s165) | (sub_sel & sub165) | (and_sel & and165) | (or_sel & or165);
  assign y166 = (add_sel & s166) | (sub_sel & sub166) | (and_sel & and166) | (or_sel & or166);
  assign y167 = (add_sel & s167) | (sub_sel & sub167) | (and_sel & and167) | (or_sel & or167);
  assign y168 = (add_sel & s168) | (sub_sel & sub168) | (and_sel & and168) | (or_sel & or168);
  assign y169 = (add_sel & s169) | (sub_sel & sub169) | (and_sel & and169) | (or_sel & or169);
  assign y170 = (add_sel & s170) | (sub_sel & sub170) | (and_sel & and170) | (or_sel & or170);
  assign y171 = (add_sel & s171) | (sub_sel & sub171) | (and_sel & and171) | (or_sel & or171);
  assign y172 = (add_sel & s172) | (sub_sel & sub172) | (and_sel & and172) | (or_sel & or172);
  assign y173 = (add_sel & s173) | (sub_sel & sub173) | (and_sel & and173) | (or_sel & or173);
  assign y174 = (add_sel & s174) | (sub_sel & sub174) | (and_sel & and174) | (or_sel & or174);
  assign y175 = (add_sel & s175) | (sub_sel & sub175) | (and_sel & and175) | (or_sel & or175);
  assign y176 = (add_sel & s176) | (sub_sel & sub176) | (and_sel & and176) | (or_sel & or176);
  assign y177 = (add_sel & s177) | (sub_sel & sub177) | (and_sel & and177) | (or_sel & or177);
  assign y178 = (add_sel & s178) | (sub_sel & sub178) | (and_sel & and178) | (or_sel & or178);
  assign y179 = (add_sel & s179) | (sub_sel & sub179) | (and_sel & and179) | (or_sel & or179);
  assign y180 = (add_sel & s180) | (sub_sel & sub180) | (and_sel & and180) | (or_sel & or180);
  assign y181 = (add_sel & s181) | (sub_sel & sub181) | (and_sel & and181) | (or_sel & or181);
  assign y182 = (add_sel & s182) | (sub_sel & sub182) | (and_sel & and182) | (or_sel & or182);
  assign y183 = (add_sel & s183) | (sub_sel & sub183) | (and_sel & and183) | (or_sel & or183);
  assign y184 = (add_sel & s184) | (sub_sel & sub184) | (and_sel & and184) | (or_sel & or184);
  assign y185 = (add_sel & s185) | (sub_sel & sub185) | (and_sel & and185) | (or_sel & or185);
  assign y186 = (add_sel & s186) | (sub_sel & sub186) | (and_sel & and186) | (or_sel & or186);
  assign y187 = (add_sel & s187) | (sub_sel & sub187) | (and_sel & and187) | (or_sel & or187);
  assign y188 = (add_sel & s188) | (sub_sel & sub188) | (and_sel & and188) | (or_sel & or188);
  assign y189 = (add_sel & s189) | (sub_sel & sub189) | (and_sel & and189) | (or_sel & or189);
  assign y190 = (add_sel & s190) | (sub_sel & sub190) | (and_sel & and190) | (or_sel & or190);
  assign y191 = (add_sel & s191) | (sub_sel & sub191) | (and_sel & and191) | (or_sel & or191);
  assign y192 = (add_sel & s192) | (sub_sel & sub192) | (and_sel & and192) | (or_sel & or192);
  assign y193 = (add_sel & s193) | (sub_sel & sub193) | (and_sel & and193) | (or_sel & or193);
  assign y194 = (add_sel & s194) | (sub_sel & sub194) | (and_sel & and194) | (or_sel & or194);
  assign y195 = (add_sel & s195) | (sub_sel & sub195) | (and_sel & and195) | (or_sel & or195);
  assign y196 = (add_sel & s196) | (sub_sel & sub196) | (and_sel & and196) | (or_sel & or196);
  assign y197 = (add_sel & s197) | (sub_sel & sub197) | (and_sel & and197) | (or_sel & or197);
  assign y198 = (add_sel & s198) | (sub_sel & sub198) | (and_sel & and198) | (or_sel & or198);
  assign y199 = (add_sel & s199) | (sub_sel & sub199) | (and_sel & and199) | (or_sel & or199);
  assign y200 = (add_sel & s200) | (sub_sel & sub200) | (and_sel & and200) | (or_sel & or200);
  assign y201 = (add_sel & s201) | (sub_sel & sub201) | (and_sel & and201) | (or_sel & or201);
  assign y202 = (add_sel & s202) | (sub_sel & sub202) | (and_sel & and202) | (or_sel & or202);
  assign y203 = (add_sel & s203) | (sub_sel & sub203) | (and_sel & and203) | (or_sel & or203);
  assign y204 = (add_sel & s204) | (sub_sel & sub204) | (and_sel & and204) | (or_sel & or204);
  assign y205 = (add_sel & s205) | (sub_sel & sub205) | (and_sel & and205) | (or_sel & or205);
  assign y206 = (add_sel & s206) | (sub_sel & sub206) | (and_sel & and206) | (or_sel & or206);
  assign y207 = (add_sel & s207) | (sub_sel & sub207) | (and_sel & and207) | (or_sel & or207);
  assign y208 = (add_sel & s208) | (sub_sel & sub208) | (and_sel & and208) | (or_sel & or208);
  assign y209 = (add_sel & s209) | (sub_sel & sub209) | (and_sel & and209) | (or_sel & or209);
  assign y210 = (add_sel & s210) | (sub_sel & sub210) | (and_sel & and210) | (or_sel & or210);
  assign y211 = (add_sel & s211) | (sub_sel & sub211) | (and_sel & and211) | (or_sel & or211);
  assign y212 = (add_sel & s212) | (sub_sel & sub212) | (and_sel & and212) | (or_sel & or212);
  assign y213 = (add_sel & s213) | (sub_sel & sub213) | (and_sel & and213) | (or_sel & or213);
  assign y214 = (add_sel & s214) | (sub_sel & sub214) | (and_sel & and214) | (or_sel & or214);
  assign y215 = (add_sel & s215) | (sub_sel & sub215) | (and_sel & and215) | (or_sel & or215);
  assign y216 = (add_sel & s216) | (sub_sel & sub216) | (and_sel & and216) | (or_sel & or216);
  assign y217 = (add_sel & s217) | (sub_sel & sub217) | (and_sel & and217) | (or_sel & or217);
  assign y218 = (add_sel & s218) | (sub_sel & sub218) | (and_sel & and218) | (or_sel & or218);
  assign y219 = (add_sel & s219) | (sub_sel & sub219) | (and_sel & and219) | (or_sel & or219);
  assign y220 = (add_sel & s220) | (sub_sel & sub220) | (and_sel & and220) | (or_sel & or220);
  assign y221 = (add_sel & s221) | (sub_sel & sub221) | (and_sel & and221) | (or_sel & or221);
  assign y222 = (add_sel & s222) | (sub_sel & sub222) | (and_sel & and222) | (or_sel & or222);
  assign y223 = (add_sel & s223) | (sub_sel & sub223) | (and_sel & and223) | (or_sel & or223);
  assign y224 = (add_sel & s224) | (sub_sel & sub224) | (and_sel & and224) | (or_sel & or224);
  assign y225 = (add_sel & s225) | (sub_sel & sub225) | (and_sel & and225) | (or_sel & or225);
  assign y226 = (add_sel & s226) | (sub_sel & sub226) | (and_sel & and226) | (or_sel & or226);
  assign y227 = (add_sel & s227) | (sub_sel & sub227) | (and_sel & and227) | (or_sel & or227);
  assign y228 = (add_sel & s228) | (sub_sel & sub228) | (and_sel & and228) | (or_sel & or228);
  assign y229 = (add_sel & s229) | (sub_sel & sub229) | (and_sel & and229) | (or_sel & or229);
  assign y230 = (add_sel & s230) | (sub_sel & sub230) | (and_sel & and230) | (or_sel & or230);
  assign y231 = (add_sel & s231) | (sub_sel & sub231) | (and_sel & and231) | (or_sel & or231);
  assign y232 = (add_sel & s232) | (sub_sel & sub232) | (and_sel & and232) | (or_sel & or232);
  assign y233 = (add_sel & s233) | (sub_sel & sub233) | (and_sel & and233) | (or_sel & or233);
  assign y234 = (add_sel & s234) | (sub_sel & sub234) | (and_sel & and234) | (or_sel & or234);
  assign y235 = (add_sel & s235) | (sub_sel & sub235) | (and_sel & and235) | (or_sel & or235);
  assign y236 = (add_sel & s236) | (sub_sel & sub236) | (and_sel & and236) | (or_sel & or236);
  assign y237 = (add_sel & s237) | (sub_sel & sub237) | (and_sel & and237) | (or_sel & or237);
  assign y238 = (add_sel & s238) | (sub_sel & sub238) | (and_sel & and238) | (or_sel & or238);
  assign y239 = (add_sel & s239) | (sub_sel & sub239) | (and_sel & and239) | (or_sel & or239);
  assign y240 = (add_sel & s240) | (sub_sel & sub240) | (and_sel & and240) | (or_sel & or240);
  assign y241 = (add_sel & s241) | (sub_sel & sub241) | (and_sel & and241) | (or_sel & or241);
  assign y242 = (add_sel & s242) | (sub_sel & sub242) | (and_sel & and242) | (or_sel & or242);
  assign y243 = (add_sel & s243) | (sub_sel & sub243) | (and_sel & and243) | (or_sel & or243);
  assign y244 = (add_sel & s244) | (sub_sel & sub244) | (and_sel & and244) | (or_sel & or244);
  assign y245 = (add_sel & s245) | (sub_sel & sub245) | (and_sel & and245) | (or_sel & or245);
  assign y246 = (add_sel & s246) | (sub_sel & sub246) | (and_sel & and246) | (or_sel & or246);
  assign y247 = (add_sel & s247) | (sub_sel & sub247) | (and_sel & and247) | (or_sel & or247);
  assign y248 = (add_sel & s248) | (sub_sel & sub248) | (and_sel & and248) | (or_sel & or248);
  assign y249 = (add_sel & s249) | (sub_sel & sub249) | (and_sel & and249) | (or_sel & or249);
  assign y250 = (add_sel & s250) | (sub_sel & sub250) | (and_sel & and250) | (or_sel & or250);
  assign y251 = (add_sel & s251) | (sub_sel & sub251) | (and_sel & and251) | (or_sel & or251);
  assign y252 = (add_sel & s252) | (sub_sel & sub252) | (and_sel & and252) | (or_sel & or252);
  assign y253 = (add_sel & s253) | (sub_sel & sub253) | (and_sel & and253) | (or_sel & or253);
  assign y254 = (add_sel & s254) | (sub_sel & sub254) | (and_sel & and254) | (or_sel & or254);
  assign y255 = (add_sel & s255) | (sub_sel & sub255) | (and_sel & and255) | (or_sel & or255);
  assign y256 = (add_sel & s256) | (sub_sel & sub256) | (and_sel & and256) | (or_sel & or256);
  assign y257 = (add_sel & s257) | (sub_sel & sub257) | (and_sel & and257) | (or_sel & or257);
  assign y258 = (add_sel & s258) | (sub_sel & sub258) | (and_sel & and258) | (or_sel & or258);
  assign y259 = (add_sel & s259) | (sub_sel & sub259) | (and_sel & and259) | (or_sel & or259);
  assign y260 = (add_sel & s260) | (sub_sel & sub260) | (and_sel & and260) | (or_sel & or260);
  assign y261 = (add_sel & s261) | (sub_sel & sub261) | (and_sel & and261) | (or_sel & or261);
  assign y262 = (add_sel & s262) | (sub_sel & sub262) | (and_sel & and262) | (or_sel & or262);
  assign y263 = (add_sel & s263) | (sub_sel & sub263) | (and_sel & and263) | (or_sel & or263);
  assign y264 = (add_sel & s264) | (sub_sel & sub264) | (and_sel & and264) | (or_sel & or264);
  assign y265 = (add_sel & s265) | (sub_sel & sub265) | (and_sel & and265) | (or_sel & or265);
  assign y266 = (add_sel & s266) | (sub_sel & sub266) | (and_sel & and266) | (or_sel & or266);
  assign y267 = (add_sel & s267) | (sub_sel & sub267) | (and_sel & and267) | (or_sel & or267);
  assign y268 = (add_sel & s268) | (sub_sel & sub268) | (and_sel & and268) | (or_sel & or268);
  assign y269 = (add_sel & s269) | (sub_sel & sub269) | (and_sel & and269) | (or_sel & or269);
  assign y270 = (add_sel & s270) | (sub_sel & sub270) | (and_sel & and270) | (or_sel & or270);
  assign y271 = (add_sel & s271) | (sub_sel & sub271) | (and_sel & and271) | (or_sel & or271);
  assign y272 = (add_sel & s272) | (sub_sel & sub272) | (and_sel & and272) | (or_sel & or272);
  assign y273 = (add_sel & s273) | (sub_sel & sub273) | (and_sel & and273) | (or_sel & or273);
  assign y274 = (add_sel & s274) | (sub_sel & sub274) | (and_sel & and274) | (or_sel & or274);
  assign y275 = (add_sel & s275) | (sub_sel & sub275) | (and_sel & and275) | (or_sel & or275);
  assign y276 = (add_sel & s276) | (sub_sel & sub276) | (and_sel & and276) | (or_sel & or276);
  assign y277 = (add_sel & s277) | (sub_sel & sub277) | (and_sel & and277) | (or_sel & or277);
  assign y278 = (add_sel & s278) | (sub_sel & sub278) | (and_sel & and278) | (or_sel & or278);
  assign y279 = (add_sel & s279) | (sub_sel & sub279) | (and_sel & and279) | (or_sel & or279);
  assign y280 = (add_sel & s280) | (sub_sel & sub280) | (and_sel & and280) | (or_sel & or280);
  assign y281 = (add_sel & s281) | (sub_sel & sub281) | (and_sel & and281) | (or_sel & or281);
  assign y282 = (add_sel & s282) | (sub_sel & sub282) | (and_sel & and282) | (or_sel & or282);
  assign y283 = (add_sel & s283) | (sub_sel & sub283) | (and_sel & and283) | (or_sel & or283);
  assign y284 = (add_sel & s284) | (sub_sel & sub284) | (and_sel & and284) | (or_sel & or284);
  assign y285 = (add_sel & s285) | (sub_sel & sub285) | (and_sel & and285) | (or_sel & or285);
  assign y286 = (add_sel & s286) | (sub_sel & sub286) | (and_sel & and286) | (or_sel & or286);
  assign y287 = (add_sel & s287) | (sub_sel & sub287) | (and_sel & and287) | (or_sel & or287);
  assign y288 = (add_sel & s288) | (sub_sel & sub288) | (and_sel & and288) | (or_sel & or288);
  assign y289 = (add_sel & s289) | (sub_sel & sub289) | (and_sel & and289) | (or_sel & or289);
  assign y290 = (add_sel & s290) | (sub_sel & sub290) | (and_sel & and290) | (or_sel & or290);
  assign y291 = (add_sel & s291) | (sub_sel & sub291) | (and_sel & and291) | (or_sel & or291);
  assign y292 = (add_sel & s292) | (sub_sel & sub292) | (and_sel & and292) | (or_sel & or292);
  assign y293 = (add_sel & s293) | (sub_sel & sub293) | (and_sel & and293) | (or_sel & or293);
  assign y294 = (add_sel & s294) | (sub_sel & sub294) | (and_sel & and294) | (or_sel & or294);
  assign y295 = (add_sel & s295) | (sub_sel & sub295) | (and_sel & and295) | (or_sel & or295);
  assign y296 = (add_sel & s296) | (sub_sel & sub296) | (and_sel & and296) | (or_sel & or296);
  assign y297 = (add_sel & s297) | (sub_sel & sub297) | (and_sel & and297) | (or_sel & or297);
  assign y298 = (add_sel & s298) | (sub_sel & sub298) | (and_sel & and298) | (or_sel & or298);
  assign y299 = (add_sel & s299) | (sub_sel & sub299) | (and_sel & and299) | (or_sel & or299);
  assign y300 = (add_sel & s300) | (sub_sel & sub300) | (and_sel & and300) | (or_sel & or300);
  assign y301 = (add_sel & s301) | (sub_sel & sub301) | (and_sel & and301) | (or_sel & or301);
  assign y302 = (add_sel & s302) | (sub_sel & sub302) | (and_sel & and302) | (or_sel & or302);
  assign y303 = (add_sel & s303) | (sub_sel & sub303) | (and_sel & and303) | (or_sel & or303);
  assign y304 = (add_sel & s304) | (sub_sel & sub304) | (and_sel & and304) | (or_sel & or304);
  assign y305 = (add_sel & s305) | (sub_sel & sub305) | (and_sel & and305) | (or_sel & or305);
  assign y306 = (add_sel & s306) | (sub_sel & sub306) | (and_sel & and306) | (or_sel & or306);
  assign y307 = (add_sel & s307) | (sub_sel & sub307) | (and_sel & and307) | (or_sel & or307);
  assign y308 = (add_sel & s308) | (sub_sel & sub308) | (and_sel & and308) | (or_sel & or308);
  assign y309 = (add_sel & s309) | (sub_sel & sub309) | (and_sel & and309) | (or_sel & or309);
  assign y310 = (add_sel & s310) | (sub_sel & sub310) | (and_sel & and310) | (or_sel & or310);
  assign y311 = (add_sel & s311) | (sub_sel & sub311) | (and_sel & and311) | (or_sel & or311);
  assign y312 = (add_sel & s312) | (sub_sel & sub312) | (and_sel & and312) | (or_sel & or312);
  assign y313 = (add_sel & s313) | (sub_sel & sub313) | (and_sel & and313) | (or_sel & or313);
  assign y314 = (add_sel & s314) | (sub_sel & sub314) | (and_sel & and314) | (or_sel & or314);
  assign y315 = (add_sel & s315) | (sub_sel & sub315) | (and_sel & and315) | (or_sel & or315);
  assign y316 = (add_sel & s316) | (sub_sel & sub316) | (and_sel & and316) | (or_sel & or316);
  assign y317 = (add_sel & s317) | (sub_sel & sub317) | (and_sel & and317) | (or_sel & or317);
  assign y318 = (add_sel & s318) | (sub_sel & sub318) | (and_sel & and318) | (or_sel & or318);
  assign y319 = (add_sel & s319) | (sub_sel & sub319) | (and_sel & and319) | (or_sel & or319);
  assign y320 = (add_sel & s320) | (sub_sel & sub320) | (and_sel & and320) | (or_sel & or320);
  assign y321 = (add_sel & s321) | (sub_sel & sub321) | (and_sel & and321) | (or_sel & or321);
  assign y322 = (add_sel & s322) | (sub_sel & sub322) | (and_sel & and322) | (or_sel & or322);
  assign y323 = (add_sel & s323) | (sub_sel & sub323) | (and_sel & and323) | (or_sel & or323);
  assign y324 = (add_sel & s324) | (sub_sel & sub324) | (and_sel & and324) | (or_sel & or324);
  assign y325 = (add_sel & s325) | (sub_sel & sub325) | (and_sel & and325) | (or_sel & or325);
  assign y326 = (add_sel & s326) | (sub_sel & sub326) | (and_sel & and326) | (or_sel & or326);
  assign y327 = (add_sel & s327) | (sub_sel & sub327) | (and_sel & and327) | (or_sel & or327);
  assign y328 = (add_sel & s328) | (sub_sel & sub328) | (and_sel & and328) | (or_sel & or328);
  assign y329 = (add_sel & s329) | (sub_sel & sub329) | (and_sel & and329) | (or_sel & or329);
  assign y330 = (add_sel & s330) | (sub_sel & sub330) | (and_sel & and330) | (or_sel & or330);
  assign y331 = (add_sel & s331) | (sub_sel & sub331) | (and_sel & and331) | (or_sel & or331);
  assign y332 = (add_sel & s332) | (sub_sel & sub332) | (and_sel & and332) | (or_sel & or332);
  assign y333 = (add_sel & s333) | (sub_sel & sub333) | (and_sel & and333) | (or_sel & or333);
  assign y334 = (add_sel & s334) | (sub_sel & sub334) | (and_sel & and334) | (or_sel & or334);
  assign y335 = (add_sel & s335) | (sub_sel & sub335) | (and_sel & and335) | (or_sel & or335);
  assign y336 = (add_sel & s336) | (sub_sel & sub336) | (and_sel & and336) | (or_sel & or336);
  assign y337 = (add_sel & s337) | (sub_sel & sub337) | (and_sel & and337) | (or_sel & or337);
  assign y338 = (add_sel & s338) | (sub_sel & sub338) | (and_sel & and338) | (or_sel & or338);
  assign y339 = (add_sel & s339) | (sub_sel & sub339) | (and_sel & and339) | (or_sel & or339);
  assign y340 = (add_sel & s340) | (sub_sel & sub340) | (and_sel & and340) | (or_sel & or340);
  assign y341 = (add_sel & s341) | (sub_sel & sub341) | (and_sel & and341) | (or_sel & or341);
  assign y342 = (add_sel & s342) | (sub_sel & sub342) | (and_sel & and342) | (or_sel & or342);
  assign y343 = (add_sel & s343) | (sub_sel & sub343) | (and_sel & and343) | (or_sel & or343);
  assign y344 = (add_sel & s344) | (sub_sel & sub344) | (and_sel & and344) | (or_sel & or344);
  assign y345 = (add_sel & s345) | (sub_sel & sub345) | (and_sel & and345) | (or_sel & or345);
  assign y346 = (add_sel & s346) | (sub_sel & sub346) | (and_sel & and346) | (or_sel & or346);
  assign y347 = (add_sel & s347) | (sub_sel & sub347) | (and_sel & and347) | (or_sel & or347);
  assign y348 = (add_sel & s348) | (sub_sel & sub348) | (and_sel & and348) | (or_sel & or348);
  assign y349 = (add_sel & s349) | (sub_sel & sub349) | (and_sel & and349) | (or_sel & or349);
  assign y350 = (add_sel & s350) | (sub_sel & sub350) | (and_sel & and350) | (or_sel & or350);
  assign y351 = (add_sel & s351) | (sub_sel & sub351) | (and_sel & and351) | (or_sel & or351);
  assign y352 = (add_sel & s352) | (sub_sel & sub352) | (and_sel & and352) | (or_sel & or352);
  assign y353 = (add_sel & s353) | (sub_sel & sub353) | (and_sel & and353) | (or_sel & or353);
  assign y354 = (add_sel & s354) | (sub_sel & sub354) | (and_sel & and354) | (or_sel & or354);
  assign y355 = (add_sel & s355) | (sub_sel & sub355) | (and_sel & and355) | (or_sel & or355);
  assign y356 = (add_sel & s356) | (sub_sel & sub356) | (and_sel & and356) | (or_sel & or356);
  assign y357 = (add_sel & s357) | (sub_sel & sub357) | (and_sel & and357) | (or_sel & or357);
  assign y358 = (add_sel & s358) | (sub_sel & sub358) | (and_sel & and358) | (or_sel & or358);
  assign y359 = (add_sel & s359) | (sub_sel & sub359) | (and_sel & and359) | (or_sel & or359);
  assign y360 = (add_sel & s360) | (sub_sel & sub360) | (and_sel & and360) | (or_sel & or360);
  assign y361 = (add_sel & s361) | (sub_sel & sub361) | (and_sel & and361) | (or_sel & or361);
  assign y362 = (add_sel & s362) | (sub_sel & sub362) | (and_sel & and362) | (or_sel & or362);
  assign y363 = (add_sel & s363) | (sub_sel & sub363) | (and_sel & and363) | (or_sel & or363);
  assign y364 = (add_sel & s364) | (sub_sel & sub364) | (and_sel & and364) | (or_sel & or364);
  assign y365 = (add_sel & s365) | (sub_sel & sub365) | (and_sel & and365) | (or_sel & or365);
  assign y366 = (add_sel & s366) | (sub_sel & sub366) | (and_sel & and366) | (or_sel & or366);
  assign y367 = (add_sel & s367) | (sub_sel & sub367) | (and_sel & and367) | (or_sel & or367);
  assign y368 = (add_sel & s368) | (sub_sel & sub368) | (and_sel & and368) | (or_sel & or368);
  assign y369 = (add_sel & s369) | (sub_sel & sub369) | (and_sel & and369) | (or_sel & or369);
  assign y370 = (add_sel & s370) | (sub_sel & sub370) | (and_sel & and370) | (or_sel & or370);
  assign y371 = (add_sel & s371) | (sub_sel & sub371) | (and_sel & and371) | (or_sel & or371);
  assign y372 = (add_sel & s372) | (sub_sel & sub372) | (and_sel & and372) | (or_sel & or372);
  assign y373 = (add_sel & s373) | (sub_sel & sub373) | (and_sel & and373) | (or_sel & or373);
  assign y374 = (add_sel & s374) | (sub_sel & sub374) | (and_sel & and374) | (or_sel & or374);
  assign y375 = (add_sel & s375) | (sub_sel & sub375) | (and_sel & and375) | (or_sel & or375);
  assign y376 = (add_sel & s376) | (sub_sel & sub376) | (and_sel & and376) | (or_sel & or376);
  assign y377 = (add_sel & s377) | (sub_sel & sub377) | (and_sel & and377) | (or_sel & or377);
  assign y378 = (add_sel & s378) | (sub_sel & sub378) | (and_sel & and378) | (or_sel & or378);
  assign y379 = (add_sel & s379) | (sub_sel & sub379) | (and_sel & and379) | (or_sel & or379);
  assign y380 = (add_sel & s380) | (sub_sel & sub380) | (and_sel & and380) | (or_sel & or380);
  assign y381 = (add_sel & s381) | (sub_sel & sub381) | (and_sel & and381) | (or_sel & or381);
  assign y382 = (add_sel & s382) | (sub_sel & sub382) | (and_sel & and382) | (or_sel & or382);
  assign y383 = (add_sel & s383) | (sub_sel & sub383) | (and_sel & and383) | (or_sel & or383);
  assign y384 = (add_sel & s384) | (sub_sel & sub384) | (and_sel & and384) | (or_sel & or384);
  assign y385 = (add_sel & s385) | (sub_sel & sub385) | (and_sel & and385) | (or_sel & or385);
  assign y386 = (add_sel & s386) | (sub_sel & sub386) | (and_sel & and386) | (or_sel & or386);
  assign y387 = (add_sel & s387) | (sub_sel & sub387) | (and_sel & and387) | (or_sel & or387);
  assign y388 = (add_sel & s388) | (sub_sel & sub388) | (and_sel & and388) | (or_sel & or388);
  assign y389 = (add_sel & s389) | (sub_sel & sub389) | (and_sel & and389) | (or_sel & or389);
  assign y390 = (add_sel & s390) | (sub_sel & sub390) | (and_sel & and390) | (or_sel & or390);
  assign y391 = (add_sel & s391) | (sub_sel & sub391) | (and_sel & and391) | (or_sel & or391);
  assign y392 = (add_sel & s392) | (sub_sel & sub392) | (and_sel & and392) | (or_sel & or392);
  assign y393 = (add_sel & s393) | (sub_sel & sub393) | (and_sel & and393) | (or_sel & or393);
  assign y394 = (add_sel & s394) | (sub_sel & sub394) | (and_sel & and394) | (or_sel & or394);
  assign y395 = (add_sel & s395) | (sub_sel & sub395) | (and_sel & and395) | (or_sel & or395);
  assign y396 = (add_sel & s396) | (sub_sel & sub396) | (and_sel & and396) | (or_sel & or396);
  assign y397 = (add_sel & s397) | (sub_sel & sub397) | (and_sel & and397) | (or_sel & or397);
  assign y398 = (add_sel & s398) | (sub_sel & sub398) | (and_sel & and398) | (or_sel & or398);
  assign y399 = (add_sel & s399) | (sub_sel & sub399) | (and_sel & and399) | (or_sel & or399);
  assign y400 = (add_sel & s400) | (sub_sel & sub400) | (and_sel & and400) | (or_sel & or400);
  assign y401 = (add_sel & s401) | (sub_sel & sub401) | (and_sel & and401) | (or_sel & or401);
  assign y402 = (add_sel & s402) | (sub_sel & sub402) | (and_sel & and402) | (or_sel & or402);
  assign y403 = (add_sel & s403) | (sub_sel & sub403) | (and_sel & and403) | (or_sel & or403);
  assign y404 = (add_sel & s404) | (sub_sel & sub404) | (and_sel & and404) | (or_sel & or404);
  assign y405 = (add_sel & s405) | (sub_sel & sub405) | (and_sel & and405) | (or_sel & or405);
  assign y406 = (add_sel & s406) | (sub_sel & sub406) | (and_sel & and406) | (or_sel & or406);
  assign y407 = (add_sel & s407) | (sub_sel & sub407) | (and_sel & and407) | (or_sel & or407);
  assign y408 = (add_sel & s408) | (sub_sel & sub408) | (and_sel & and408) | (or_sel & or408);
  assign y409 = (add_sel & s409) | (sub_sel & sub409) | (and_sel & and409) | (or_sel & or409);
  assign y410 = (add_sel & s410) | (sub_sel & sub410) | (and_sel & and410) | (or_sel & or410);
  assign y411 = (add_sel & s411) | (sub_sel & sub411) | (and_sel & and411) | (or_sel & or411);
  assign y412 = (add_sel & s412) | (sub_sel & sub412) | (and_sel & and412) | (or_sel & or412);
  assign y413 = (add_sel & s413) | (sub_sel & sub413) | (and_sel & and413) | (or_sel & or413);
  assign y414 = (add_sel & s414) | (sub_sel & sub414) | (and_sel & and414) | (or_sel & or414);
  assign y415 = (add_sel & s415) | (sub_sel & sub415) | (and_sel & and415) | (or_sel & or415);
  assign y416 = (add_sel & s416) | (sub_sel & sub416) | (and_sel & and416) | (or_sel & or416);
  assign y417 = (add_sel & s417) | (sub_sel & sub417) | (and_sel & and417) | (or_sel & or417);
  assign y418 = (add_sel & s418) | (sub_sel & sub418) | (and_sel & and418) | (or_sel & or418);
  assign y419 = (add_sel & s419) | (sub_sel & sub419) | (and_sel & and419) | (or_sel & or419);
  assign y420 = (add_sel & s420) | (sub_sel & sub420) | (and_sel & and420) | (or_sel & or420);
  assign y421 = (add_sel & s421) | (sub_sel & sub421) | (and_sel & and421) | (or_sel & or421);
  assign y422 = (add_sel & s422) | (sub_sel & sub422) | (and_sel & and422) | (or_sel & or422);
  assign y423 = (add_sel & s423) | (sub_sel & sub423) | (and_sel & and423) | (or_sel & or423);
  assign y424 = (add_sel & s424) | (sub_sel & sub424) | (and_sel & and424) | (or_sel & or424);
  assign y425 = (add_sel & s425) | (sub_sel & sub425) | (and_sel & and425) | (or_sel & or425);
  assign y426 = (add_sel & s426) | (sub_sel & sub426) | (and_sel & and426) | (or_sel & or426);
  assign y427 = (add_sel & s427) | (sub_sel & sub427) | (and_sel & and427) | (or_sel & or427);
  assign y428 = (add_sel & s428) | (sub_sel & sub428) | (and_sel & and428) | (or_sel & or428);
  assign y429 = (add_sel & s429) | (sub_sel & sub429) | (and_sel & and429) | (or_sel & or429);
  assign y430 = (add_sel & s430) | (sub_sel & sub430) | (and_sel & and430) | (or_sel & or430);
  assign y431 = (add_sel & s431) | (sub_sel & sub431) | (and_sel & and431) | (or_sel & or431);
  assign y432 = (add_sel & s432) | (sub_sel & sub432) | (and_sel & and432) | (or_sel & or432);
  assign y433 = (add_sel & s433) | (sub_sel & sub433) | (and_sel & and433) | (or_sel & or433);
  assign y434 = (add_sel & s434) | (sub_sel & sub434) | (and_sel & and434) | (or_sel & or434);
  assign y435 = (add_sel & s435) | (sub_sel & sub435) | (and_sel & and435) | (or_sel & or435);
  assign y436 = (add_sel & s436) | (sub_sel & sub436) | (and_sel & and436) | (or_sel & or436);
  assign y437 = (add_sel & s437) | (sub_sel & sub437) | (and_sel & and437) | (or_sel & or437);
  assign y438 = (add_sel & s438) | (sub_sel & sub438) | (and_sel & and438) | (or_sel & or438);
  assign y439 = (add_sel & s439) | (sub_sel & sub439) | (and_sel & and439) | (or_sel & or439);
  assign y440 = (add_sel & s440) | (sub_sel & sub440) | (and_sel & and440) | (or_sel & or440);
  assign y441 = (add_sel & s441) | (sub_sel & sub441) | (and_sel & and441) | (or_sel & or441);
  assign y442 = (add_sel & s442) | (sub_sel & sub442) | (and_sel & and442) | (or_sel & or442);
  assign y443 = (add_sel & s443) | (sub_sel & sub443) | (and_sel & and443) | (or_sel & or443);
  assign y444 = (add_sel & s444) | (sub_sel & sub444) | (and_sel & and444) | (or_sel & or444);
  assign y445 = (add_sel & s445) | (sub_sel & sub445) | (and_sel & and445) | (or_sel & or445);
  assign y446 = (add_sel & s446) | (sub_sel & sub446) | (and_sel & and446) | (or_sel & or446);
  assign y447 = (add_sel & s447) | (sub_sel & sub447) | (and_sel & and447) | (or_sel & or447);
  assign y448 = (add_sel & s448) | (sub_sel & sub448) | (and_sel & and448) | (or_sel & or448);
  assign y449 = (add_sel & s449) | (sub_sel & sub449) | (and_sel & and449) | (or_sel & or449);
  assign y450 = (add_sel & s450) | (sub_sel & sub450) | (and_sel & and450) | (or_sel & or450);
  assign y451 = (add_sel & s451) | (sub_sel & sub451) | (and_sel & and451) | (or_sel & or451);
  assign y452 = (add_sel & s452) | (sub_sel & sub452) | (and_sel & and452) | (or_sel & or452);
  assign y453 = (add_sel & s453) | (sub_sel & sub453) | (and_sel & and453) | (or_sel & or453);
  assign y454 = (add_sel & s454) | (sub_sel & sub454) | (and_sel & and454) | (or_sel & or454);
  assign y455 = (add_sel & s455) | (sub_sel & sub455) | (and_sel & and455) | (or_sel & or455);
  assign y456 = (add_sel & s456) | (sub_sel & sub456) | (and_sel & and456) | (or_sel & or456);
  assign y457 = (add_sel & s457) | (sub_sel & sub457) | (and_sel & and457) | (or_sel & or457);
  assign y458 = (add_sel & s458) | (sub_sel & sub458) | (and_sel & and458) | (or_sel & or458);
  assign y459 = (add_sel & s459) | (sub_sel & sub459) | (and_sel & and459) | (or_sel & or459);
  assign y460 = (add_sel & s460) | (sub_sel & sub460) | (and_sel & and460) | (or_sel & or460);
  assign y461 = (add_sel & s461) | (sub_sel & sub461) | (and_sel & and461) | (or_sel & or461);
  assign y462 = (add_sel & s462) | (sub_sel & sub462) | (and_sel & and462) | (or_sel & or462);
  assign y463 = (add_sel & s463) | (sub_sel & sub463) | (and_sel & and463) | (or_sel & or463);
  assign y464 = (add_sel & s464) | (sub_sel & sub464) | (and_sel & and464) | (or_sel & or464);
  assign y465 = (add_sel & s465) | (sub_sel & sub465) | (and_sel & and465) | (or_sel & or465);
  assign y466 = (add_sel & s466) | (sub_sel & sub466) | (and_sel & and466) | (or_sel & or466);
  assign y467 = (add_sel & s467) | (sub_sel & sub467) | (and_sel & and467) | (or_sel & or467);
  assign y468 = (add_sel & s468) | (sub_sel & sub468) | (and_sel & and468) | (or_sel & or468);
  assign y469 = (add_sel & s469) | (sub_sel & sub469) | (and_sel & and469) | (or_sel & or469);
  assign y470 = (add_sel & s470) | (sub_sel & sub470) | (and_sel & and470) | (or_sel & or470);
  assign y471 = (add_sel & s471) | (sub_sel & sub471) | (and_sel & and471) | (or_sel & or471);
  assign y472 = (add_sel & s472) | (sub_sel & sub472) | (and_sel & and472) | (or_sel & or472);
  assign y473 = (add_sel & s473) | (sub_sel & sub473) | (and_sel & and473) | (or_sel & or473);
  assign y474 = (add_sel & s474) | (sub_sel & sub474) | (and_sel & and474) | (or_sel & or474);
  assign y475 = (add_sel & s475) | (sub_sel & sub475) | (and_sel & and475) | (or_sel & or475);
  assign y476 = (add_sel & s476) | (sub_sel & sub476) | (and_sel & and476) | (or_sel & or476);
  assign y477 = (add_sel & s477) | (sub_sel & sub477) | (and_sel & and477) | (or_sel & or477);
  assign y478 = (add_sel & s478) | (sub_sel & sub478) | (and_sel & and478) | (or_sel & or478);
  assign y479 = (add_sel & s479) | (sub_sel & sub479) | (and_sel & and479) | (or_sel & or479);
  assign y480 = (add_sel & s480) | (sub_sel & sub480) | (and_sel & and480) | (or_sel & or480);
  assign y481 = (add_sel & s481) | (sub_sel & sub481) | (and_sel & and481) | (or_sel & or481);
  assign y482 = (add_sel & s482) | (sub_sel & sub482) | (and_sel & and482) | (or_sel & or482);
  assign y483 = (add_sel & s483) | (sub_sel & sub483) | (and_sel & and483) | (or_sel & or483);
  assign y484 = (add_sel & s484) | (sub_sel & sub484) | (and_sel & and484) | (or_sel & or484);
  assign y485 = (add_sel & s485) | (sub_sel & sub485) | (and_sel & and485) | (or_sel & or485);
  assign y486 = (add_sel & s486) | (sub_sel & sub486) | (and_sel & and486) | (or_sel & or486);
  assign y487 = (add_sel & s487) | (sub_sel & sub487) | (and_sel & and487) | (or_sel & or487);
  assign y488 = (add_sel & s488) | (sub_sel & sub488) | (and_sel & and488) | (or_sel & or488);
  assign y489 = (add_sel & s489) | (sub_sel & sub489) | (and_sel & and489) | (or_sel & or489);
  assign y490 = (add_sel & s490) | (sub_sel & sub490) | (and_sel & and490) | (or_sel & or490);
  assign y491 = (add_sel & s491) | (sub_sel & sub491) | (and_sel & and491) | (or_sel & or491);
  assign y492 = (add_sel & s492) | (sub_sel & sub492) | (and_sel & and492) | (or_sel & or492);
  assign y493 = (add_sel & s493) | (sub_sel & sub493) | (and_sel & and493) | (or_sel & or493);
  assign y494 = (add_sel & s494) | (sub_sel & sub494) | (and_sel & and494) | (or_sel & or494);
  assign y495 = (add_sel & s495) | (sub_sel & sub495) | (and_sel & and495) | (or_sel & or495);
  assign y496 = (add_sel & s496) | (sub_sel & sub496) | (and_sel & and496) | (or_sel & or496);
  assign y497 = (add_sel & s497) | (sub_sel & sub497) | (and_sel & and497) | (or_sel & or497);
  assign y498 = (add_sel & s498) | (sub_sel & sub498) | (and_sel & and498) | (or_sel & or498);
  assign y499 = (add_sel & s499) | (sub_sel & sub499) | (and_sel & and499) | (or_sel & or499);
  assign y500 = (add_sel & s500) | (sub_sel & sub500) | (and_sel & and500) | (or_sel & or500);
  assign y501 = (add_sel & s501) | (sub_sel & sub501) | (and_sel & and501) | (or_sel & or501);
  assign y502 = (add_sel & s502) | (sub_sel & sub502) | (and_sel & and502) | (or_sel & or502);
  assign y503 = (add_sel & s503) | (sub_sel & sub503) | (and_sel & and503) | (or_sel & or503);
  assign y504 = (add_sel & s504) | (sub_sel & sub504) | (and_sel & and504) | (or_sel & or504);
  assign y505 = (add_sel & s505) | (sub_sel & sub505) | (and_sel & and505) | (or_sel & or505);
  assign y506 = (add_sel & s506) | (sub_sel & sub506) | (and_sel & and506) | (or_sel & or506);
  assign y507 = (add_sel & s507) | (sub_sel & sub507) | (and_sel & and507) | (or_sel & or507);
  assign y508 = (add_sel & s508) | (sub_sel & sub508) | (and_sel & and508) | (or_sel & or508);
  assign y509 = (add_sel & s509) | (sub_sel & sub509) | (and_sel & and509) | (or_sel & or509);
  assign y510 = (add_sel & s510) | (sub_sel & sub510) | (and_sel & and510) | (or_sel & or510);
  assign y511 = (add_sel & s511) | (sub_sel & sub511) | (and_sel & and511) | (or_sel & or511);
  assign y512 = (add_sel & s512) | (sub_sel & sub512) | (and_sel & and512) | (or_sel & or512);
  assign y513 = (add_sel & s513) | (sub_sel & sub513) | (and_sel & and513) | (or_sel & or513);
  assign y514 = (add_sel & s514) | (sub_sel & sub514) | (and_sel & and514) | (or_sel & or514);
  assign y515 = (add_sel & s515) | (sub_sel & sub515) | (and_sel & and515) | (or_sel & or515);
  assign y516 = (add_sel & s516) | (sub_sel & sub516) | (and_sel & and516) | (or_sel & or516);
  assign y517 = (add_sel & s517) | (sub_sel & sub517) | (and_sel & and517) | (or_sel & or517);
  assign y518 = (add_sel & s518) | (sub_sel & sub518) | (and_sel & and518) | (or_sel & or518);
  assign y519 = (add_sel & s519) | (sub_sel & sub519) | (and_sel & and519) | (or_sel & or519);
  assign y520 = (add_sel & s520) | (sub_sel & sub520) | (and_sel & and520) | (or_sel & or520);
  assign y521 = (add_sel & s521) | (sub_sel & sub521) | (and_sel & and521) | (or_sel & or521);
  assign y522 = (add_sel & s522) | (sub_sel & sub522) | (and_sel & and522) | (or_sel & or522);
  assign y523 = (add_sel & s523) | (sub_sel & sub523) | (and_sel & and523) | (or_sel & or523);
  assign y524 = (add_sel & s524) | (sub_sel & sub524) | (and_sel & and524) | (or_sel & or524);
  assign y525 = (add_sel & s525) | (sub_sel & sub525) | (and_sel & and525) | (or_sel & or525);
  assign y526 = (add_sel & s526) | (sub_sel & sub526) | (and_sel & and526) | (or_sel & or526);
  assign y527 = (add_sel & s527) | (sub_sel & sub527) | (and_sel & and527) | (or_sel & or527);
  assign y528 = (add_sel & s528) | (sub_sel & sub528) | (and_sel & and528) | (or_sel & or528);
  assign y529 = (add_sel & s529) | (sub_sel & sub529) | (and_sel & and529) | (or_sel & or529);
  assign y530 = (add_sel & s530) | (sub_sel & sub530) | (and_sel & and530) | (or_sel & or530);
  assign y531 = (add_sel & s531) | (sub_sel & sub531) | (and_sel & and531) | (or_sel & or531);
  assign y532 = (add_sel & s532) | (sub_sel & sub532) | (and_sel & and532) | (or_sel & or532);
  assign y533 = (add_sel & s533) | (sub_sel & sub533) | (and_sel & and533) | (or_sel & or533);
  assign y534 = (add_sel & s534) | (sub_sel & sub534) | (and_sel & and534) | (or_sel & or534);
  assign y535 = (add_sel & s535) | (sub_sel & sub535) | (and_sel & and535) | (or_sel & or535);
  assign y536 = (add_sel & s536) | (sub_sel & sub536) | (and_sel & and536) | (or_sel & or536);
  assign y537 = (add_sel & s537) | (sub_sel & sub537) | (and_sel & and537) | (or_sel & or537);
  assign y538 = (add_sel & s538) | (sub_sel & sub538) | (and_sel & and538) | (or_sel & or538);
  assign y539 = (add_sel & s539) | (sub_sel & sub539) | (and_sel & and539) | (or_sel & or539);
  assign y540 = (add_sel & s540) | (sub_sel & sub540) | (and_sel & and540) | (or_sel & or540);
  assign y541 = (add_sel & s541) | (sub_sel & sub541) | (and_sel & and541) | (or_sel & or541);
  assign y542 = (add_sel & s542) | (sub_sel & sub542) | (and_sel & and542) | (or_sel & or542);
  assign y543 = (add_sel & s543) | (sub_sel & sub543) | (and_sel & and543) | (or_sel & or543);
  assign y544 = (add_sel & s544) | (sub_sel & sub544) | (and_sel & and544) | (or_sel & or544);
  assign y545 = (add_sel & s545) | (sub_sel & sub545) | (and_sel & and545) | (or_sel & or545);
  assign y546 = (add_sel & s546) | (sub_sel & sub546) | (and_sel & and546) | (or_sel & or546);
  assign y547 = (add_sel & s547) | (sub_sel & sub547) | (and_sel & and547) | (or_sel & or547);
  assign y548 = (add_sel & s548) | (sub_sel & sub548) | (and_sel & and548) | (or_sel & or548);
  assign y549 = (add_sel & s549) | (sub_sel & sub549) | (and_sel & and549) | (or_sel & or549);
  assign y550 = (add_sel & s550) | (sub_sel & sub550) | (and_sel & and550) | (or_sel & or550);
  assign y551 = (add_sel & s551) | (sub_sel & sub551) | (and_sel & and551) | (or_sel & or551);
  assign y552 = (add_sel & s552) | (sub_sel & sub552) | (and_sel & and552) | (or_sel & or552);
  assign y553 = (add_sel & s553) | (sub_sel & sub553) | (and_sel & and553) | (or_sel & or553);
  assign y554 = (add_sel & s554) | (sub_sel & sub554) | (and_sel & and554) | (or_sel & or554);
  assign y555 = (add_sel & s555) | (sub_sel & sub555) | (and_sel & and555) | (or_sel & or555);
  assign y556 = (add_sel & s556) | (sub_sel & sub556) | (and_sel & and556) | (or_sel & or556);
  assign y557 = (add_sel & s557) | (sub_sel & sub557) | (and_sel & and557) | (or_sel & or557);
  assign y558 = (add_sel & s558) | (sub_sel & sub558) | (and_sel & and558) | (or_sel & or558);
  assign y559 = (add_sel & s559) | (sub_sel & sub559) | (and_sel & and559) | (or_sel & or559);
  assign y560 = (add_sel & s560) | (sub_sel & sub560) | (and_sel & and560) | (or_sel & or560);
  assign y561 = (add_sel & s561) | (sub_sel & sub561) | (and_sel & and561) | (or_sel & or561);
  assign y562 = (add_sel & s562) | (sub_sel & sub562) | (and_sel & and562) | (or_sel & or562);
  assign y563 = (add_sel & s563) | (sub_sel & sub563) | (and_sel & and563) | (or_sel & or563);
  assign y564 = (add_sel & s564) | (sub_sel & sub564) | (and_sel & and564) | (or_sel & or564);
  assign y565 = (add_sel & s565) | (sub_sel & sub565) | (and_sel & and565) | (or_sel & or565);
  assign y566 = (add_sel & s566) | (sub_sel & sub566) | (and_sel & and566) | (or_sel & or566);
  assign y567 = (add_sel & s567) | (sub_sel & sub567) | (and_sel & and567) | (or_sel & or567);
  assign y568 = (add_sel & s568) | (sub_sel & sub568) | (and_sel & and568) | (or_sel & or568);
  assign y569 = (add_sel & s569) | (sub_sel & sub569) | (and_sel & and569) | (or_sel & or569);
  assign y570 = (add_sel & s570) | (sub_sel & sub570) | (and_sel & and570) | (or_sel & or570);
  assign y571 = (add_sel & s571) | (sub_sel & sub571) | (and_sel & and571) | (or_sel & or571);
  assign y572 = (add_sel & s572) | (sub_sel & sub572) | (and_sel & and572) | (or_sel & or572);
  assign y573 = (add_sel & s573) | (sub_sel & sub573) | (and_sel & and573) | (or_sel & or573);
  assign y574 = (add_sel & s574) | (sub_sel & sub574) | (and_sel & and574) | (or_sel & or574);
  assign y575 = (add_sel & s575) | (sub_sel & sub575) | (and_sel & and575) | (or_sel & or575);
  assign y576 = (add_sel & s576) | (sub_sel & sub576) | (and_sel & and576) | (or_sel & or576);
  assign y577 = (add_sel & s577) | (sub_sel & sub577) | (and_sel & and577) | (or_sel & or577);
  assign y578 = (add_sel & s578) | (sub_sel & sub578) | (and_sel & and578) | (or_sel & or578);
  assign y579 = (add_sel & s579) | (sub_sel & sub579) | (and_sel & and579) | (or_sel & or579);
  assign y580 = (add_sel & s580) | (sub_sel & sub580) | (and_sel & and580) | (or_sel & or580);
  assign y581 = (add_sel & s581) | (sub_sel & sub581) | (and_sel & and581) | (or_sel & or581);
  assign y582 = (add_sel & s582) | (sub_sel & sub582) | (and_sel & and582) | (or_sel & or582);
  assign y583 = (add_sel & s583) | (sub_sel & sub583) | (and_sel & and583) | (or_sel & or583);
  assign y584 = (add_sel & s584) | (sub_sel & sub584) | (and_sel & and584) | (or_sel & or584);
  assign y585 = (add_sel & s585) | (sub_sel & sub585) | (and_sel & and585) | (or_sel & or585);
  assign y586 = (add_sel & s586) | (sub_sel & sub586) | (and_sel & and586) | (or_sel & or586);
  assign y587 = (add_sel & s587) | (sub_sel & sub587) | (and_sel & and587) | (or_sel & or587);
  assign y588 = (add_sel & s588) | (sub_sel & sub588) | (and_sel & and588) | (or_sel & or588);
  assign y589 = (add_sel & s589) | (sub_sel & sub589) | (and_sel & and589) | (or_sel & or589);
  assign y590 = (add_sel & s590) | (sub_sel & sub590) | (and_sel & and590) | (or_sel & or590);
  assign y591 = (add_sel & s591) | (sub_sel & sub591) | (and_sel & and591) | (or_sel & or591);
  assign y592 = (add_sel & s592) | (sub_sel & sub592) | (and_sel & and592) | (or_sel & or592);
  assign y593 = (add_sel & s593) | (sub_sel & sub593) | (and_sel & and593) | (or_sel & or593);
  assign y594 = (add_sel & s594) | (sub_sel & sub594) | (and_sel & and594) | (or_sel & or594);
  assign y595 = (add_sel & s595) | (sub_sel & sub595) | (and_sel & and595) | (or_sel & or595);
  assign y596 = (add_sel & s596) | (sub_sel & sub596) | (and_sel & and596) | (or_sel & or596);
  assign y597 = (add_sel & s597) | (sub_sel & sub597) | (and_sel & and597) | (or_sel & or597);
  assign y598 = (add_sel & s598) | (sub_sel & sub598) | (and_sel & and598) | (or_sel & or598);
  assign y599 = (add_sel & s599) | (sub_sel & sub599) | (and_sel & and599) | (or_sel & or599);
  assign y600 = (add_sel & s600) | (sub_sel & sub600) | (and_sel & and600) | (or_sel & or600);
  assign y601 = (add_sel & s601) | (sub_sel & sub601) | (and_sel & and601) | (or_sel & or601);
  assign y602 = (add_sel & s602) | (sub_sel & sub602) | (and_sel & and602) | (or_sel & or602);
  assign y603 = (add_sel & s603) | (sub_sel & sub603) | (and_sel & and603) | (or_sel & or603);
  assign y604 = (add_sel & s604) | (sub_sel & sub604) | (and_sel & and604) | (or_sel & or604);
  assign y605 = (add_sel & s605) | (sub_sel & sub605) | (and_sel & and605) | (or_sel & or605);
  assign y606 = (add_sel & s606) | (sub_sel & sub606) | (and_sel & and606) | (or_sel & or606);
  assign y607 = (add_sel & s607) | (sub_sel & sub607) | (and_sel & and607) | (or_sel & or607);
  assign y608 = (add_sel & s608) | (sub_sel & sub608) | (and_sel & and608) | (or_sel & or608);
  assign y609 = (add_sel & s609) | (sub_sel & sub609) | (and_sel & and609) | (or_sel & or609);
  assign y610 = (add_sel & s610) | (sub_sel & sub610) | (and_sel & and610) | (or_sel & or610);
  assign y611 = (add_sel & s611) | (sub_sel & sub611) | (and_sel & and611) | (or_sel & or611);
  assign y612 = (add_sel & s612) | (sub_sel & sub612) | (and_sel & and612) | (or_sel & or612);
  assign y613 = (add_sel & s613) | (sub_sel & sub613) | (and_sel & and613) | (or_sel & or613);
  assign y614 = (add_sel & s614) | (sub_sel & sub614) | (and_sel & and614) | (or_sel & or614);
  assign y615 = (add_sel & s615) | (sub_sel & sub615) | (and_sel & and615) | (or_sel & or615);
  assign y616 = (add_sel & s616) | (sub_sel & sub616) | (and_sel & and616) | (or_sel & or616);
  assign y617 = (add_sel & s617) | (sub_sel & sub617) | (and_sel & and617) | (or_sel & or617);
  assign y618 = (add_sel & s618) | (sub_sel & sub618) | (and_sel & and618) | (or_sel & or618);
  assign y619 = (add_sel & s619) | (sub_sel & sub619) | (and_sel & and619) | (or_sel & or619);
  assign y620 = (add_sel & s620) | (sub_sel & sub620) | (and_sel & and620) | (or_sel & or620);
  assign y621 = (add_sel & s621) | (sub_sel & sub621) | (and_sel & and621) | (or_sel & or621);
  assign y622 = (add_sel & s622) | (sub_sel & sub622) | (and_sel & and622) | (or_sel & or622);
  assign y623 = (add_sel & s623) | (sub_sel & sub623) | (and_sel & and623) | (or_sel & or623);
  assign y624 = (add_sel & s624) | (sub_sel & sub624) | (and_sel & and624) | (or_sel & or624);
  assign y625 = (add_sel & s625) | (sub_sel & sub625) | (and_sel & and625) | (or_sel & or625);
  assign y626 = (add_sel & s626) | (sub_sel & sub626) | (and_sel & and626) | (or_sel & or626);
  assign y627 = (add_sel & s627) | (sub_sel & sub627) | (and_sel & and627) | (or_sel & or627);
  assign y628 = (add_sel & s628) | (sub_sel & sub628) | (and_sel & and628) | (or_sel & or628);
  assign y629 = (add_sel & s629) | (sub_sel & sub629) | (and_sel & and629) | (or_sel & or629);
  assign y630 = (add_sel & s630) | (sub_sel & sub630) | (and_sel & and630) | (or_sel & or630);
  assign y631 = (add_sel & s631) | (sub_sel & sub631) | (and_sel & and631) | (or_sel & or631);
  assign y632 = (add_sel & s632) | (sub_sel & sub632) | (and_sel & and632) | (or_sel & or632);
  assign y633 = (add_sel & s633) | (sub_sel & sub633) | (and_sel & and633) | (or_sel & or633);
  assign y634 = (add_sel & s634) | (sub_sel & sub634) | (and_sel & and634) | (or_sel & or634);
  assign y635 = (add_sel & s635) | (sub_sel & sub635) | (and_sel & and635) | (or_sel & or635);
  assign y636 = (add_sel & s636) | (sub_sel & sub636) | (and_sel & and636) | (or_sel & or636);
  assign y637 = (add_sel & s637) | (sub_sel & sub637) | (and_sel & and637) | (or_sel & or637);
  assign y638 = (add_sel & s638) | (sub_sel & sub638) | (and_sel & and638) | (or_sel & or638);
  assign y639 = (add_sel & s639) | (sub_sel & sub639) | (and_sel & and639) | (or_sel & or639);
  assign y640 = (add_sel & s640) | (sub_sel & sub640) | (and_sel & and640) | (or_sel & or640);
  assign y641 = (add_sel & s641) | (sub_sel & sub641) | (and_sel & and641) | (or_sel & or641);
  assign y642 = (add_sel & s642) | (sub_sel & sub642) | (and_sel & and642) | (or_sel & or642);
  assign y643 = (add_sel & s643) | (sub_sel & sub643) | (and_sel & and643) | (or_sel & or643);
  assign y644 = (add_sel & s644) | (sub_sel & sub644) | (and_sel & and644) | (or_sel & or644);
  assign y645 = (add_sel & s645) | (sub_sel & sub645) | (and_sel & and645) | (or_sel & or645);
  assign y646 = (add_sel & s646) | (sub_sel & sub646) | (and_sel & and646) | (or_sel & or646);
  assign y647 = (add_sel & s647) | (sub_sel & sub647) | (and_sel & and647) | (or_sel & or647);
  assign y648 = (add_sel & s648) | (sub_sel & sub648) | (and_sel & and648) | (or_sel & or648);
  assign y649 = (add_sel & s649) | (sub_sel & sub649) | (and_sel & and649) | (or_sel & or649);
  assign y650 = (add_sel & s650) | (sub_sel & sub650) | (and_sel & and650) | (or_sel & or650);
  assign y651 = (add_sel & s651) | (sub_sel & sub651) | (and_sel & and651) | (or_sel & or651);
  assign y652 = (add_sel & s652) | (sub_sel & sub652) | (and_sel & and652) | (or_sel & or652);
  assign y653 = (add_sel & s653) | (sub_sel & sub653) | (and_sel & and653) | (or_sel & or653);
  assign y654 = (add_sel & s654) | (sub_sel & sub654) | (and_sel & and654) | (or_sel & or654);
  assign y655 = (add_sel & s655) | (sub_sel & sub655) | (and_sel & and655) | (or_sel & or655);
  assign y656 = (add_sel & s656) | (sub_sel & sub656) | (and_sel & and656) | (or_sel & or656);
  assign y657 = (add_sel & s657) | (sub_sel & sub657) | (and_sel & and657) | (or_sel & or657);
  assign y658 = (add_sel & s658) | (sub_sel & sub658) | (and_sel & and658) | (or_sel & or658);
  assign y659 = (add_sel & s659) | (sub_sel & sub659) | (and_sel & and659) | (or_sel & or659);
  assign y660 = (add_sel & s660) | (sub_sel & sub660) | (and_sel & and660) | (or_sel & or660);
  assign y661 = (add_sel & s661) | (sub_sel & sub661) | (and_sel & and661) | (or_sel & or661);
  assign y662 = (add_sel & s662) | (sub_sel & sub662) | (and_sel & and662) | (or_sel & or662);
  assign y663 = (add_sel & s663) | (sub_sel & sub663) | (and_sel & and663) | (or_sel & or663);
  assign y664 = (add_sel & s664) | (sub_sel & sub664) | (and_sel & and664) | (or_sel & or664);
  assign y665 = (add_sel & s665) | (sub_sel & sub665) | (and_sel & and665) | (or_sel & or665);
  assign y666 = (add_sel & s666) | (sub_sel & sub666) | (and_sel & and666) | (or_sel & or666);
  assign y667 = (add_sel & s667) | (sub_sel & sub667) | (and_sel & and667) | (or_sel & or667);
  assign y668 = (add_sel & s668) | (sub_sel & sub668) | (and_sel & and668) | (or_sel & or668);
  assign y669 = (add_sel & s669) | (sub_sel & sub669) | (and_sel & and669) | (or_sel & or669);
  assign y670 = (add_sel & s670) | (sub_sel & sub670) | (and_sel & and670) | (or_sel & or670);
  assign y671 = (add_sel & s671) | (sub_sel & sub671) | (and_sel & and671) | (or_sel & or671);
  assign y672 = (add_sel & s672) | (sub_sel & sub672) | (and_sel & and672) | (or_sel & or672);
  assign y673 = (add_sel & s673) | (sub_sel & sub673) | (and_sel & and673) | (or_sel & or673);
  assign y674 = (add_sel & s674) | (sub_sel & sub674) | (and_sel & and674) | (or_sel & or674);
  assign y675 = (add_sel & s675) | (sub_sel & sub675) | (and_sel & and675) | (or_sel & or675);
  assign y676 = (add_sel & s676) | (sub_sel & sub676) | (and_sel & and676) | (or_sel & or676);
  assign y677 = (add_sel & s677) | (sub_sel & sub677) | (and_sel & and677) | (or_sel & or677);
  assign y678 = (add_sel & s678) | (sub_sel & sub678) | (and_sel & and678) | (or_sel & or678);
  assign y679 = (add_sel & s679) | (sub_sel & sub679) | (and_sel & and679) | (or_sel & or679);
  assign y680 = (add_sel & s680) | (sub_sel & sub680) | (and_sel & and680) | (or_sel & or680);
  assign y681 = (add_sel & s681) | (sub_sel & sub681) | (and_sel & and681) | (or_sel & or681);
  assign y682 = (add_sel & s682) | (sub_sel & sub682) | (and_sel & and682) | (or_sel & or682);
  assign y683 = (add_sel & s683) | (sub_sel & sub683) | (and_sel & and683) | (or_sel & or683);
  assign y684 = (add_sel & s684) | (sub_sel & sub684) | (and_sel & and684) | (or_sel & or684);
  assign y685 = (add_sel & s685) | (sub_sel & sub685) | (and_sel & and685) | (or_sel & or685);
  assign y686 = (add_sel & s686) | (sub_sel & sub686) | (and_sel & and686) | (or_sel & or686);
  assign y687 = (add_sel & s687) | (sub_sel & sub687) | (and_sel & and687) | (or_sel & or687);
  assign y688 = (add_sel & s688) | (sub_sel & sub688) | (and_sel & and688) | (or_sel & or688);
  assign y689 = (add_sel & s689) | (sub_sel & sub689) | (and_sel & and689) | (or_sel & or689);
  assign y690 = (add_sel & s690) | (sub_sel & sub690) | (and_sel & and690) | (or_sel & or690);
  assign y691 = (add_sel & s691) | (sub_sel & sub691) | (and_sel & and691) | (or_sel & or691);
  assign y692 = (add_sel & s692) | (sub_sel & sub692) | (and_sel & and692) | (or_sel & or692);
  assign y693 = (add_sel & s693) | (sub_sel & sub693) | (and_sel & and693) | (or_sel & or693);
  assign y694 = (add_sel & s694) | (sub_sel & sub694) | (and_sel & and694) | (or_sel & or694);
  assign y695 = (add_sel & s695) | (sub_sel & sub695) | (and_sel & and695) | (or_sel & or695);
  assign y696 = (add_sel & s696) | (sub_sel & sub696) | (and_sel & and696) | (or_sel & or696);
  assign y697 = (add_sel & s697) | (sub_sel & sub697) | (and_sel & and697) | (or_sel & or697);
  assign y698 = (add_sel & s698) | (sub_sel & sub698) | (and_sel & and698) | (or_sel & or698);
  assign y699 = (add_sel & s699) | (sub_sel & sub699) | (and_sel & and699) | (or_sel & or699);
  assign y700 = (add_sel & s700) | (sub_sel & sub700) | (and_sel & and700) | (or_sel & or700);
  assign y701 = (add_sel & s701) | (sub_sel & sub701) | (and_sel & and701) | (or_sel & or701);
  assign y702 = (add_sel & s702) | (sub_sel & sub702) | (and_sel & and702) | (or_sel & or702);
  assign y703 = (add_sel & s703) | (sub_sel & sub703) | (and_sel & and703) | (or_sel & or703);
  assign y704 = (add_sel & s704) | (sub_sel & sub704) | (and_sel & and704) | (or_sel & or704);
  assign y705 = (add_sel & s705) | (sub_sel & sub705) | (and_sel & and705) | (or_sel & or705);
  assign y706 = (add_sel & s706) | (sub_sel & sub706) | (and_sel & and706) | (or_sel & or706);
  assign y707 = (add_sel & s707) | (sub_sel & sub707) | (and_sel & and707) | (or_sel & or707);
  assign y708 = (add_sel & s708) | (sub_sel & sub708) | (and_sel & and708) | (or_sel & or708);
  assign y709 = (add_sel & s709) | (sub_sel & sub709) | (and_sel & and709) | (or_sel & or709);
  assign y710 = (add_sel & s710) | (sub_sel & sub710) | (and_sel & and710) | (or_sel & or710);
  assign y711 = (add_sel & s711) | (sub_sel & sub711) | (and_sel & and711) | (or_sel & or711);
  assign y712 = (add_sel & s712) | (sub_sel & sub712) | (and_sel & and712) | (or_sel & or712);
  assign y713 = (add_sel & s713) | (sub_sel & sub713) | (and_sel & and713) | (or_sel & or713);
  assign y714 = (add_sel & s714) | (sub_sel & sub714) | (and_sel & and714) | (or_sel & or714);
  assign y715 = (add_sel & s715) | (sub_sel & sub715) | (and_sel & and715) | (or_sel & or715);
  assign y716 = (add_sel & s716) | (sub_sel & sub716) | (and_sel & and716) | (or_sel & or716);
  assign y717 = (add_sel & s717) | (sub_sel & sub717) | (and_sel & and717) | (or_sel & or717);
  assign y718 = (add_sel & s718) | (sub_sel & sub718) | (and_sel & and718) | (or_sel & or718);
  assign y719 = (add_sel & s719) | (sub_sel & sub719) | (and_sel & and719) | (or_sel & or719);
  assign y720 = (add_sel & s720) | (sub_sel & sub720) | (and_sel & and720) | (or_sel & or720);
  assign y721 = (add_sel & s721) | (sub_sel & sub721) | (and_sel & and721) | (or_sel & or721);
  assign y722 = (add_sel & s722) | (sub_sel & sub722) | (and_sel & and722) | (or_sel & or722);
  assign y723 = (add_sel & s723) | (sub_sel & sub723) | (and_sel & and723) | (or_sel & or723);
  assign y724 = (add_sel & s724) | (sub_sel & sub724) | (and_sel & and724) | (or_sel & or724);
  assign y725 = (add_sel & s725) | (sub_sel & sub725) | (and_sel & and725) | (or_sel & or725);
  assign y726 = (add_sel & s726) | (sub_sel & sub726) | (and_sel & and726) | (or_sel & or726);
  assign y727 = (add_sel & s727) | (sub_sel & sub727) | (and_sel & and727) | (or_sel & or727);
  assign y728 = (add_sel & s728) | (sub_sel & sub728) | (and_sel & and728) | (or_sel & or728);
  assign y729 = (add_sel & s729) | (sub_sel & sub729) | (and_sel & and729) | (or_sel & or729);
  assign y730 = (add_sel & s730) | (sub_sel & sub730) | (and_sel & and730) | (or_sel & or730);
  assign y731 = (add_sel & s731) | (sub_sel & sub731) | (and_sel & and731) | (or_sel & or731);
  assign y732 = (add_sel & s732) | (sub_sel & sub732) | (and_sel & and732) | (or_sel & or732);
  assign y733 = (add_sel & s733) | (sub_sel & sub733) | (and_sel & and733) | (or_sel & or733);
  assign y734 = (add_sel & s734) | (sub_sel & sub734) | (and_sel & and734) | (or_sel & or734);
  assign y735 = (add_sel & s735) | (sub_sel & sub735) | (and_sel & and735) | (or_sel & or735);
  assign y736 = (add_sel & s736) | (sub_sel & sub736) | (and_sel & and736) | (or_sel & or736);
  assign y737 = (add_sel & s737) | (sub_sel & sub737) | (and_sel & and737) | (or_sel & or737);
  assign y738 = (add_sel & s738) | (sub_sel & sub738) | (and_sel & and738) | (or_sel & or738);
  assign y739 = (add_sel & s739) | (sub_sel & sub739) | (and_sel & and739) | (or_sel & or739);
  assign y740 = (add_sel & s740) | (sub_sel & sub740) | (and_sel & and740) | (or_sel & or740);
  assign y741 = (add_sel & s741) | (sub_sel & sub741) | (and_sel & and741) | (or_sel & or741);
  assign y742 = (add_sel & s742) | (sub_sel & sub742) | (and_sel & and742) | (or_sel & or742);
  assign y743 = (add_sel & s743) | (sub_sel & sub743) | (and_sel & and743) | (or_sel & or743);
  assign y744 = (add_sel & s744) | (sub_sel & sub744) | (and_sel & and744) | (or_sel & or744);
  assign y745 = (add_sel & s745) | (sub_sel & sub745) | (and_sel & and745) | (or_sel & or745);
  assign y746 = (add_sel & s746) | (sub_sel & sub746) | (and_sel & and746) | (or_sel & or746);
  assign y747 = (add_sel & s747) | (sub_sel & sub747) | (and_sel & and747) | (or_sel & or747);
  assign y748 = (add_sel & s748) | (sub_sel & sub748) | (and_sel & and748) | (or_sel & or748);
  assign y749 = (add_sel & s749) | (sub_sel & sub749) | (and_sel & and749) | (or_sel & or749);
  assign y750 = (add_sel & s750) | (sub_sel & sub750) | (and_sel & and750) | (or_sel & or750);
  assign y751 = (add_sel & s751) | (sub_sel & sub751) | (and_sel & and751) | (or_sel & or751);
  assign y752 = (add_sel & s752) | (sub_sel & sub752) | (and_sel & and752) | (or_sel & or752);
  assign y753 = (add_sel & s753) | (sub_sel & sub753) | (and_sel & and753) | (or_sel & or753);
  assign y754 = (add_sel & s754) | (sub_sel & sub754) | (and_sel & and754) | (or_sel & or754);
  assign y755 = (add_sel & s755) | (sub_sel & sub755) | (and_sel & and755) | (or_sel & or755);
  assign y756 = (add_sel & s756) | (sub_sel & sub756) | (and_sel & and756) | (or_sel & or756);
  assign y757 = (add_sel & s757) | (sub_sel & sub757) | (and_sel & and757) | (or_sel & or757);
  assign y758 = (add_sel & s758) | (sub_sel & sub758) | (and_sel & and758) | (or_sel & or758);
  assign y759 = (add_sel & s759) | (sub_sel & sub759) | (and_sel & and759) | (or_sel & or759);
  assign y760 = (add_sel & s760) | (sub_sel & sub760) | (and_sel & and760) | (or_sel & or760);
  assign y761 = (add_sel & s761) | (sub_sel & sub761) | (and_sel & and761) | (or_sel & or761);
  assign y762 = (add_sel & s762) | (sub_sel & sub762) | (and_sel & and762) | (or_sel & or762);
  assign y763 = (add_sel & s763) | (sub_sel & sub763) | (and_sel & and763) | (or_sel & or763);
  assign y764 = (add_sel & s764) | (sub_sel & sub764) | (and_sel & and764) | (or_sel & or764);
  assign y765 = (add_sel & s765) | (sub_sel & sub765) | (and_sel & and765) | (or_sel & or765);
  assign y766 = (add_sel & s766) | (sub_sel & sub766) | (and_sel & and766) | (or_sel & or766);
  assign y767 = (add_sel & s767) | (sub_sel & sub767) | (and_sel & and767) | (or_sel & or767);
  assign y768 = (add_sel & s768) | (sub_sel & sub768) | (and_sel & and768) | (or_sel & or768);
  assign y769 = (add_sel & s769) | (sub_sel & sub769) | (and_sel & and769) | (or_sel & or769);
  assign y770 = (add_sel & s770) | (sub_sel & sub770) | (and_sel & and770) | (or_sel & or770);
  assign y771 = (add_sel & s771) | (sub_sel & sub771) | (and_sel & and771) | (or_sel & or771);
  assign y772 = (add_sel & s772) | (sub_sel & sub772) | (and_sel & and772) | (or_sel & or772);
  assign y773 = (add_sel & s773) | (sub_sel & sub773) | (and_sel & and773) | (or_sel & or773);
  assign y774 = (add_sel & s774) | (sub_sel & sub774) | (and_sel & and774) | (or_sel & or774);
  assign y775 = (add_sel & s775) | (sub_sel & sub775) | (and_sel & and775) | (or_sel & or775);
  assign y776 = (add_sel & s776) | (sub_sel & sub776) | (and_sel & and776) | (or_sel & or776);
  assign y777 = (add_sel & s777) | (sub_sel & sub777) | (and_sel & and777) | (or_sel & or777);
  assign y778 = (add_sel & s778) | (sub_sel & sub778) | (and_sel & and778) | (or_sel & or778);
  assign y779 = (add_sel & s779) | (sub_sel & sub779) | (and_sel & and779) | (or_sel & or779);
  assign y780 = (add_sel & s780) | (sub_sel & sub780) | (and_sel & and780) | (or_sel & or780);
  assign y781 = (add_sel & s781) | (sub_sel & sub781) | (and_sel & and781) | (or_sel & or781);
  assign y782 = (add_sel & s782) | (sub_sel & sub782) | (and_sel & and782) | (or_sel & or782);
  assign y783 = (add_sel & s783) | (sub_sel & sub783) | (and_sel & and783) | (or_sel & or783);
  assign y784 = (add_sel & s784) | (sub_sel & sub784) | (and_sel & and784) | (or_sel & or784);
  assign y785 = (add_sel & s785) | (sub_sel & sub785) | (and_sel & and785) | (or_sel & or785);
  assign y786 = (add_sel & s786) | (sub_sel & sub786) | (and_sel & and786) | (or_sel & or786);
  assign y787 = (add_sel & s787) | (sub_sel & sub787) | (and_sel & and787) | (or_sel & or787);
  assign y788 = (add_sel & s788) | (sub_sel & sub788) | (and_sel & and788) | (or_sel & or788);
  assign y789 = (add_sel & s789) | (sub_sel & sub789) | (and_sel & and789) | (or_sel & or789);
  assign y790 = (add_sel & s790) | (sub_sel & sub790) | (and_sel & and790) | (or_sel & or790);
  assign y791 = (add_sel & s791) | (sub_sel & sub791) | (and_sel & and791) | (or_sel & or791);
  assign y792 = (add_sel & s792) | (sub_sel & sub792) | (and_sel & and792) | (or_sel & or792);
  assign y793 = (add_sel & s793) | (sub_sel & sub793) | (and_sel & and793) | (or_sel & or793);
  assign y794 = (add_sel & s794) | (sub_sel & sub794) | (and_sel & and794) | (or_sel & or794);
  assign y795 = (add_sel & s795) | (sub_sel & sub795) | (and_sel & and795) | (or_sel & or795);
  assign y796 = (add_sel & s796) | (sub_sel & sub796) | (and_sel & and796) | (or_sel & or796);
  assign y797 = (add_sel & s797) | (sub_sel & sub797) | (and_sel & and797) | (or_sel & or797);
  assign y798 = (add_sel & s798) | (sub_sel & sub798) | (and_sel & and798) | (or_sel & or798);
  assign y799 = (add_sel & s799) | (sub_sel & sub799) | (and_sel & and799) | (or_sel & or799);
  assign y800 = (add_sel & s800) | (sub_sel & sub800) | (and_sel & and800) | (or_sel & or800);
  assign y801 = (add_sel & s801) | (sub_sel & sub801) | (and_sel & and801) | (or_sel & or801);
  assign y802 = (add_sel & s802) | (sub_sel & sub802) | (and_sel & and802) | (or_sel & or802);
  assign y803 = (add_sel & s803) | (sub_sel & sub803) | (and_sel & and803) | (or_sel & or803);
  assign y804 = (add_sel & s804) | (sub_sel & sub804) | (and_sel & and804) | (or_sel & or804);
  assign y805 = (add_sel & s805) | (sub_sel & sub805) | (and_sel & and805) | (or_sel & or805);
  assign y806 = (add_sel & s806) | (sub_sel & sub806) | (and_sel & and806) | (or_sel & or806);
  assign y807 = (add_sel & s807) | (sub_sel & sub807) | (and_sel & and807) | (or_sel & or807);
  assign y808 = (add_sel & s808) | (sub_sel & sub808) | (and_sel & and808) | (or_sel & or808);
  assign y809 = (add_sel & s809) | (sub_sel & sub809) | (and_sel & and809) | (or_sel & or809);
  assign y810 = (add_sel & s810) | (sub_sel & sub810) | (and_sel & and810) | (or_sel & or810);
  assign y811 = (add_sel & s811) | (sub_sel & sub811) | (and_sel & and811) | (or_sel & or811);
  assign y812 = (add_sel & s812) | (sub_sel & sub812) | (and_sel & and812) | (or_sel & or812);
  assign y813 = (add_sel & s813) | (sub_sel & sub813) | (and_sel & and813) | (or_sel & or813);
  assign y814 = (add_sel & s814) | (sub_sel & sub814) | (and_sel & and814) | (or_sel & or814);
  assign y815 = (add_sel & s815) | (sub_sel & sub815) | (and_sel & and815) | (or_sel & or815);
  assign y816 = (add_sel & s816) | (sub_sel & sub816) | (and_sel & and816) | (or_sel & or816);
  assign y817 = (add_sel & s817) | (sub_sel & sub817) | (and_sel & and817) | (or_sel & or817);
  assign y818 = (add_sel & s818) | (sub_sel & sub818) | (and_sel & and818) | (or_sel & or818);
  assign y819 = (add_sel & s819) | (sub_sel & sub819) | (and_sel & and819) | (or_sel & or819);
  assign y820 = (add_sel & s820) | (sub_sel & sub820) | (and_sel & and820) | (or_sel & or820);
  assign y821 = (add_sel & s821) | (sub_sel & sub821) | (and_sel & and821) | (or_sel & or821);
  assign y822 = (add_sel & s822) | (sub_sel & sub822) | (and_sel & and822) | (or_sel & or822);
  assign y823 = (add_sel & s823) | (sub_sel & sub823) | (and_sel & and823) | (or_sel & or823);
  assign y824 = (add_sel & s824) | (sub_sel & sub824) | (and_sel & and824) | (or_sel & or824);
  assign y825 = (add_sel & s825) | (sub_sel & sub825) | (and_sel & and825) | (or_sel & or825);
  assign y826 = (add_sel & s826) | (sub_sel & sub826) | (and_sel & and826) | (or_sel & or826);
  assign y827 = (add_sel & s827) | (sub_sel & sub827) | (and_sel & and827) | (or_sel & or827);
  assign y828 = (add_sel & s828) | (sub_sel & sub828) | (and_sel & and828) | (or_sel & or828);
  assign y829 = (add_sel & s829) | (sub_sel & sub829) | (and_sel & and829) | (or_sel & or829);
  assign y830 = (add_sel & s830) | (sub_sel & sub830) | (and_sel & and830) | (or_sel & or830);
  assign y831 = (add_sel & s831) | (sub_sel & sub831) | (and_sel & and831) | (or_sel & or831);
  assign y832 = (add_sel & s832) | (sub_sel & sub832) | (and_sel & and832) | (or_sel & or832);
  assign y833 = (add_sel & s833) | (sub_sel & sub833) | (and_sel & and833) | (or_sel & or833);
  assign y834 = (add_sel & s834) | (sub_sel & sub834) | (and_sel & and834) | (or_sel & or834);
  assign y835 = (add_sel & s835) | (sub_sel & sub835) | (and_sel & and835) | (or_sel & or835);
  assign y836 = (add_sel & s836) | (sub_sel & sub836) | (and_sel & and836) | (or_sel & or836);
  assign y837 = (add_sel & s837) | (sub_sel & sub837) | (and_sel & and837) | (or_sel & or837);
  assign y838 = (add_sel & s838) | (sub_sel & sub838) | (and_sel & and838) | (or_sel & or838);
  assign y839 = (add_sel & s839) | (sub_sel & sub839) | (and_sel & and839) | (or_sel & or839);
  assign y840 = (add_sel & s840) | (sub_sel & sub840) | (and_sel & and840) | (or_sel & or840);
  assign y841 = (add_sel & s841) | (sub_sel & sub841) | (and_sel & and841) | (or_sel & or841);
  assign y842 = (add_sel & s842) | (sub_sel & sub842) | (and_sel & and842) | (or_sel & or842);
  assign y843 = (add_sel & s843) | (sub_sel & sub843) | (and_sel & and843) | (or_sel & or843);
  assign y844 = (add_sel & s844) | (sub_sel & sub844) | (and_sel & and844) | (or_sel & or844);
  assign y845 = (add_sel & s845) | (sub_sel & sub845) | (and_sel & and845) | (or_sel & or845);
  assign y846 = (add_sel & s846) | (sub_sel & sub846) | (and_sel & and846) | (or_sel & or846);
  assign y847 = (add_sel & s847) | (sub_sel & sub847) | (and_sel & and847) | (or_sel & or847);
  assign y848 = (add_sel & s848) | (sub_sel & sub848) | (and_sel & and848) | (or_sel & or848);
  assign y849 = (add_sel & s849) | (sub_sel & sub849) | (and_sel & and849) | (or_sel & or849);
  assign y850 = (add_sel & s850) | (sub_sel & sub850) | (and_sel & and850) | (or_sel & or850);
  assign y851 = (add_sel & s851) | (sub_sel & sub851) | (and_sel & and851) | (or_sel & or851);
  assign y852 = (add_sel & s852) | (sub_sel & sub852) | (and_sel & and852) | (or_sel & or852);
  assign y853 = (add_sel & s853) | (sub_sel & sub853) | (and_sel & and853) | (or_sel & or853);
  assign y854 = (add_sel & s854) | (sub_sel & sub854) | (and_sel & and854) | (or_sel & or854);
  assign y855 = (add_sel & s855) | (sub_sel & sub855) | (and_sel & and855) | (or_sel & or855);
  assign y856 = (add_sel & s856) | (sub_sel & sub856) | (and_sel & and856) | (or_sel & or856);
  assign y857 = (add_sel & s857) | (sub_sel & sub857) | (and_sel & and857) | (or_sel & or857);
  assign y858 = (add_sel & s858) | (sub_sel & sub858) | (and_sel & and858) | (or_sel & or858);
  assign y859 = (add_sel & s859) | (sub_sel & sub859) | (and_sel & and859) | (or_sel & or859);
  assign y860 = (add_sel & s860) | (sub_sel & sub860) | (and_sel & and860) | (or_sel & or860);
  assign y861 = (add_sel & s861) | (sub_sel & sub861) | (and_sel & and861) | (or_sel & or861);
  assign y862 = (add_sel & s862) | (sub_sel & sub862) | (and_sel & and862) | (or_sel & or862);
  assign y863 = (add_sel & s863) | (sub_sel & sub863) | (and_sel & and863) | (or_sel & or863);
  assign y864 = (add_sel & s864) | (sub_sel & sub864) | (and_sel & and864) | (or_sel & or864);
  assign y865 = (add_sel & s865) | (sub_sel & sub865) | (and_sel & and865) | (or_sel & or865);
  assign y866 = (add_sel & s866) | (sub_sel & sub866) | (and_sel & and866) | (or_sel & or866);
  assign y867 = (add_sel & s867) | (sub_sel & sub867) | (and_sel & and867) | (or_sel & or867);
  assign y868 = (add_sel & s868) | (sub_sel & sub868) | (and_sel & and868) | (or_sel & or868);
  assign y869 = (add_sel & s869) | (sub_sel & sub869) | (and_sel & and869) | (or_sel & or869);
  assign y870 = (add_sel & s870) | (sub_sel & sub870) | (and_sel & and870) | (or_sel & or870);
  assign y871 = (add_sel & s871) | (sub_sel & sub871) | (and_sel & and871) | (or_sel & or871);
  assign y872 = (add_sel & s872) | (sub_sel & sub872) | (and_sel & and872) | (or_sel & or872);
  assign y873 = (add_sel & s873) | (sub_sel & sub873) | (and_sel & and873) | (or_sel & or873);
  assign y874 = (add_sel & s874) | (sub_sel & sub874) | (and_sel & and874) | (or_sel & or874);
  assign y875 = (add_sel & s875) | (sub_sel & sub875) | (and_sel & and875) | (or_sel & or875);
  assign y876 = (add_sel & s876) | (sub_sel & sub876) | (and_sel & and876) | (or_sel & or876);
  assign y877 = (add_sel & s877) | (sub_sel & sub877) | (and_sel & and877) | (or_sel & or877);
  assign y878 = (add_sel & s878) | (sub_sel & sub878) | (and_sel & and878) | (or_sel & or878);
  assign y879 = (add_sel & s879) | (sub_sel & sub879) | (and_sel & and879) | (or_sel & or879);
  assign y880 = (add_sel & s880) | (sub_sel & sub880) | (and_sel & and880) | (or_sel & or880);
  assign y881 = (add_sel & s881) | (sub_sel & sub881) | (and_sel & and881) | (or_sel & or881);
  assign y882 = (add_sel & s882) | (sub_sel & sub882) | (and_sel & and882) | (or_sel & or882);
  assign y883 = (add_sel & s883) | (sub_sel & sub883) | (and_sel & and883) | (or_sel & or883);
  assign y884 = (add_sel & s884) | (sub_sel & sub884) | (and_sel & and884) | (or_sel & or884);
  assign y885 = (add_sel & s885) | (sub_sel & sub885) | (and_sel & and885) | (or_sel & or885);
  assign y886 = (add_sel & s886) | (sub_sel & sub886) | (and_sel & and886) | (or_sel & or886);
  assign y887 = (add_sel & s887) | (sub_sel & sub887) | (and_sel & and887) | (or_sel & or887);
  assign y888 = (add_sel & s888) | (sub_sel & sub888) | (and_sel & and888) | (or_sel & or888);
  assign y889 = (add_sel & s889) | (sub_sel & sub889) | (and_sel & and889) | (or_sel & or889);
  assign y890 = (add_sel & s890) | (sub_sel & sub890) | (and_sel & and890) | (or_sel & or890);
  assign y891 = (add_sel & s891) | (sub_sel & sub891) | (and_sel & and891) | (or_sel & or891);
  assign y892 = (add_sel & s892) | (sub_sel & sub892) | (and_sel & and892) | (or_sel & or892);
  assign y893 = (add_sel & s893) | (sub_sel & sub893) | (and_sel & and893) | (or_sel & or893);
  assign y894 = (add_sel & s894) | (sub_sel & sub894) | (and_sel & and894) | (or_sel & or894);
  assign y895 = (add_sel & s895) | (sub_sel & sub895) | (and_sel & and895) | (or_sel & or895);
  assign y896 = (add_sel & s896) | (sub_sel & sub896) | (and_sel & and896) | (or_sel & or896);
  assign y897 = (add_sel & s897) | (sub_sel & sub897) | (and_sel & and897) | (or_sel & or897);
  assign y898 = (add_sel & s898) | (sub_sel & sub898) | (and_sel & and898) | (or_sel & or898);
  assign y899 = (add_sel & s899) | (sub_sel & sub899) | (and_sel & and899) | (or_sel & or899);
  assign y900 = (add_sel & s900) | (sub_sel & sub900) | (and_sel & and900) | (or_sel & or900);
  assign y901 = (add_sel & s901) | (sub_sel & sub901) | (and_sel & and901) | (or_sel & or901);
  assign y902 = (add_sel & s902) | (sub_sel & sub902) | (and_sel & and902) | (or_sel & or902);
  assign y903 = (add_sel & s903) | (sub_sel & sub903) | (and_sel & and903) | (or_sel & or903);
  assign y904 = (add_sel & s904) | (sub_sel & sub904) | (and_sel & and904) | (or_sel & or904);
  assign y905 = (add_sel & s905) | (sub_sel & sub905) | (and_sel & and905) | (or_sel & or905);
  assign y906 = (add_sel & s906) | (sub_sel & sub906) | (and_sel & and906) | (or_sel & or906);
  assign y907 = (add_sel & s907) | (sub_sel & sub907) | (and_sel & and907) | (or_sel & or907);
  assign y908 = (add_sel & s908) | (sub_sel & sub908) | (and_sel & and908) | (or_sel & or908);
  assign y909 = (add_sel & s909) | (sub_sel & sub909) | (and_sel & and909) | (or_sel & or909);
  assign y910 = (add_sel & s910) | (sub_sel & sub910) | (and_sel & and910) | (or_sel & or910);
  assign y911 = (add_sel & s911) | (sub_sel & sub911) | (and_sel & and911) | (or_sel & or911);
  assign y912 = (add_sel & s912) | (sub_sel & sub912) | (and_sel & and912) | (or_sel & or912);
  assign y913 = (add_sel & s913) | (sub_sel & sub913) | (and_sel & and913) | (or_sel & or913);
  assign y914 = (add_sel & s914) | (sub_sel & sub914) | (and_sel & and914) | (or_sel & or914);
  assign y915 = (add_sel & s915) | (sub_sel & sub915) | (and_sel & and915) | (or_sel & or915);
  assign y916 = (add_sel & s916) | (sub_sel & sub916) | (and_sel & and916) | (or_sel & or916);
  assign y917 = (add_sel & s917) | (sub_sel & sub917) | (and_sel & and917) | (or_sel & or917);
  assign y918 = (add_sel & s918) | (sub_sel & sub918) | (and_sel & and918) | (or_sel & or918);
  assign y919 = (add_sel & s919) | (sub_sel & sub919) | (and_sel & and919) | (or_sel & or919);
  assign y920 = (add_sel & s920) | (sub_sel & sub920) | (and_sel & and920) | (or_sel & or920);
  assign y921 = (add_sel & s921) | (sub_sel & sub921) | (and_sel & and921) | (or_sel & or921);
  assign y922 = (add_sel & s922) | (sub_sel & sub922) | (and_sel & and922) | (or_sel & or922);
  assign y923 = (add_sel & s923) | (sub_sel & sub923) | (and_sel & and923) | (or_sel & or923);
  assign y924 = (add_sel & s924) | (sub_sel & sub924) | (and_sel & and924) | (or_sel & or924);
  assign y925 = (add_sel & s925) | (sub_sel & sub925) | (and_sel & and925) | (or_sel & or925);
  assign y926 = (add_sel & s926) | (sub_sel & sub926) | (and_sel & and926) | (or_sel & or926);
  assign y927 = (add_sel & s927) | (sub_sel & sub927) | (and_sel & and927) | (or_sel & or927);
  assign y928 = (add_sel & s928) | (sub_sel & sub928) | (and_sel & and928) | (or_sel & or928);
  assign y929 = (add_sel & s929) | (sub_sel & sub929) | (and_sel & and929) | (or_sel & or929);
  assign y930 = (add_sel & s930) | (sub_sel & sub930) | (and_sel & and930) | (or_sel & or930);
  assign y931 = (add_sel & s931) | (sub_sel & sub931) | (and_sel & and931) | (or_sel & or931);
  assign y932 = (add_sel & s932) | (sub_sel & sub932) | (and_sel & and932) | (or_sel & or932);
  assign y933 = (add_sel & s933) | (sub_sel & sub933) | (and_sel & and933) | (or_sel & or933);
  assign y934 = (add_sel & s934) | (sub_sel & sub934) | (and_sel & and934) | (or_sel & or934);
  assign y935 = (add_sel & s935) | (sub_sel & sub935) | (and_sel & and935) | (or_sel & or935);
  assign y936 = (add_sel & s936) | (sub_sel & sub936) | (and_sel & and936) | (or_sel & or936);
  assign y937 = (add_sel & s937) | (sub_sel & sub937) | (and_sel & and937) | (or_sel & or937);
  assign y938 = (add_sel & s938) | (sub_sel & sub938) | (and_sel & and938) | (or_sel & or938);
  assign y939 = (add_sel & s939) | (sub_sel & sub939) | (and_sel & and939) | (or_sel & or939);
  assign y940 = (add_sel & s940) | (sub_sel & sub940) | (and_sel & and940) | (or_sel & or940);
  assign y941 = (add_sel & s941) | (sub_sel & sub941) | (and_sel & and941) | (or_sel & or941);
  assign y942 = (add_sel & s942) | (sub_sel & sub942) | (and_sel & and942) | (or_sel & or942);
  assign y943 = (add_sel & s943) | (sub_sel & sub943) | (and_sel & and943) | (or_sel & or943);
  assign y944 = (add_sel & s944) | (sub_sel & sub944) | (and_sel & and944) | (or_sel & or944);
  assign y945 = (add_sel & s945) | (sub_sel & sub945) | (and_sel & and945) | (or_sel & or945);
  assign y946 = (add_sel & s946) | (sub_sel & sub946) | (and_sel & and946) | (or_sel & or946);
  assign y947 = (add_sel & s947) | (sub_sel & sub947) | (and_sel & and947) | (or_sel & or947);
  assign y948 = (add_sel & s948) | (sub_sel & sub948) | (and_sel & and948) | (or_sel & or948);
  assign y949 = (add_sel & s949) | (sub_sel & sub949) | (and_sel & and949) | (or_sel & or949);
  assign y950 = (add_sel & s950) | (sub_sel & sub950) | (and_sel & and950) | (or_sel & or950);
  assign y951 = (add_sel & s951) | (sub_sel & sub951) | (and_sel & and951) | (or_sel & or951);
  assign y952 = (add_sel & s952) | (sub_sel & sub952) | (and_sel & and952) | (or_sel & or952);
  assign y953 = (add_sel & s953) | (sub_sel & sub953) | (and_sel & and953) | (or_sel & or953);
  assign y954 = (add_sel & s954) | (sub_sel & sub954) | (and_sel & and954) | (or_sel & or954);
  assign y955 = (add_sel & s955) | (sub_sel & sub955) | (and_sel & and955) | (or_sel & or955);
  assign y956 = (add_sel & s956) | (sub_sel & sub956) | (and_sel & and956) | (or_sel & or956);
  assign y957 = (add_sel & s957) | (sub_sel & sub957) | (and_sel & and957) | (or_sel & or957);
  assign y958 = (add_sel & s958) | (sub_sel & sub958) | (and_sel & and958) | (or_sel & or958);
  assign y959 = (add_sel & s959) | (sub_sel & sub959) | (and_sel & and959) | (or_sel & or959);
  assign y960 = (add_sel & s960) | (sub_sel & sub960) | (and_sel & and960) | (or_sel & or960);
  assign y961 = (add_sel & s961) | (sub_sel & sub961) | (and_sel & and961) | (or_sel & or961);
  assign y962 = (add_sel & s962) | (sub_sel & sub962) | (and_sel & and962) | (or_sel & or962);
  assign y963 = (add_sel & s963) | (sub_sel & sub963) | (and_sel & and963) | (or_sel & or963);
  assign y964 = (add_sel & s964) | (sub_sel & sub964) | (and_sel & and964) | (or_sel & or964);
  assign y965 = (add_sel & s965) | (sub_sel & sub965) | (and_sel & and965) | (or_sel & or965);
  assign y966 = (add_sel & s966) | (sub_sel & sub966) | (and_sel & and966) | (or_sel & or966);
  assign y967 = (add_sel & s967) | (sub_sel & sub967) | (and_sel & and967) | (or_sel & or967);
  assign y968 = (add_sel & s968) | (sub_sel & sub968) | (and_sel & and968) | (or_sel & or968);
  assign y969 = (add_sel & s969) | (sub_sel & sub969) | (and_sel & and969) | (or_sel & or969);
  assign y970 = (add_sel & s970) | (sub_sel & sub970) | (and_sel & and970) | (or_sel & or970);
  assign y971 = (add_sel & s971) | (sub_sel & sub971) | (and_sel & and971) | (or_sel & or971);
  assign y972 = (add_sel & s972) | (sub_sel & sub972) | (and_sel & and972) | (or_sel & or972);
  assign y973 = (add_sel & s973) | (sub_sel & sub973) | (and_sel & and973) | (or_sel & or973);
  assign y974 = (add_sel & s974) | (sub_sel & sub974) | (and_sel & and974) | (or_sel & or974);
  assign y975 = (add_sel & s975) | (sub_sel & sub975) | (and_sel & and975) | (or_sel & or975);
  assign y976 = (add_sel & s976) | (sub_sel & sub976) | (and_sel & and976) | (or_sel & or976);
  assign y977 = (add_sel & s977) | (sub_sel & sub977) | (and_sel & and977) | (or_sel & or977);
  assign y978 = (add_sel & s978) | (sub_sel & sub978) | (and_sel & and978) | (or_sel & or978);
  assign y979 = (add_sel & s979) | (sub_sel & sub979) | (and_sel & and979) | (or_sel & or979);
  assign y980 = (add_sel & s980) | (sub_sel & sub980) | (and_sel & and980) | (or_sel & or980);
  assign y981 = (add_sel & s981) | (sub_sel & sub981) | (and_sel & and981) | (or_sel & or981);
  assign y982 = (add_sel & s982) | (sub_sel & sub982) | (and_sel & and982) | (or_sel & or982);
  assign y983 = (add_sel & s983) | (sub_sel & sub983) | (and_sel & and983) | (or_sel & or983);
  assign y984 = (add_sel & s984) | (sub_sel & sub984) | (and_sel & and984) | (or_sel & or984);
  assign y985 = (add_sel & s985) | (sub_sel & sub985) | (and_sel & and985) | (or_sel & or985);
  assign y986 = (add_sel & s986) | (sub_sel & sub986) | (and_sel & and986) | (or_sel & or986);
  assign y987 = (add_sel & s987) | (sub_sel & sub987) | (and_sel & and987) | (or_sel & or987);
  assign y988 = (add_sel & s988) | (sub_sel & sub988) | (and_sel & and988) | (or_sel & or988);
  assign y989 = (add_sel & s989) | (sub_sel & sub989) | (and_sel & and989) | (or_sel & or989);
  assign y990 = (add_sel & s990) | (sub_sel & sub990) | (and_sel & and990) | (or_sel & or990);
  assign y991 = (add_sel & s991) | (sub_sel & sub991) | (and_sel & and991) | (or_sel & or991);
  assign y992 = (add_sel & s992) | (sub_sel & sub992) | (and_sel & and992) | (or_sel & or992);
  assign y993 = (add_sel & s993) | (sub_sel & sub993) | (and_sel & and993) | (or_sel & or993);
  assign y994 = (add_sel & s994) | (sub_sel & sub994) | (and_sel & and994) | (or_sel & or994);
  assign y995 = (add_sel & s995) | (sub_sel & sub995) | (and_sel & and995) | (or_sel & or995);
  assign y996 = (add_sel & s996) | (sub_sel & sub996) | (and_sel & and996) | (or_sel & or996);
  assign y997 = (add_sel & s997) | (sub_sel & sub997) | (and_sel & and997) | (or_sel & or997);
  assign y998 = (add_sel & s998) | (sub_sel & sub998) | (and_sel & and998) | (or_sel & or998);
  assign y999 = (add_sel & s999) | (sub_sel & sub999) | (and_sel & and999) | (or_sel & or999);
  assign y1000 = (add_sel & s1000) | (sub_sel & sub1000) | (and_sel & and1000) | (or_sel & or1000);
  assign y1001 = (add_sel & s1001) | (sub_sel & sub1001) | (and_sel & and1001) | (or_sel & or1001);
  assign y1002 = (add_sel & s1002) | (sub_sel & sub1002) | (and_sel & and1002) | (or_sel & or1002);
  assign y1003 = (add_sel & s1003) | (sub_sel & sub1003) | (and_sel & and1003) | (or_sel & or1003);
  assign y1004 = (add_sel & s1004) | (sub_sel & sub1004) | (and_sel & and1004) | (or_sel & or1004);
  assign y1005 = (add_sel & s1005) | (sub_sel & sub1005) | (and_sel & and1005) | (or_sel & or1005);
  assign y1006 = (add_sel & s1006) | (sub_sel & sub1006) | (and_sel & and1006) | (or_sel & or1006);
  assign y1007 = (add_sel & s1007) | (sub_sel & sub1007) | (and_sel & and1007) | (or_sel & or1007);
  assign y1008 = (add_sel & s1008) | (sub_sel & sub1008) | (and_sel & and1008) | (or_sel & or1008);
  assign y1009 = (add_sel & s1009) | (sub_sel & sub1009) | (and_sel & and1009) | (or_sel & or1009);
  assign y1010 = (add_sel & s1010) | (sub_sel & sub1010) | (and_sel & and1010) | (or_sel & or1010);
  assign y1011 = (add_sel & s1011) | (sub_sel & sub1011) | (and_sel & and1011) | (or_sel & or1011);
  assign y1012 = (add_sel & s1012) | (sub_sel & sub1012) | (and_sel & and1012) | (or_sel & or1012);
  assign y1013 = (add_sel & s1013) | (sub_sel & sub1013) | (and_sel & and1013) | (or_sel & or1013);
  assign y1014 = (add_sel & s1014) | (sub_sel & sub1014) | (and_sel & and1014) | (or_sel & or1014);
  assign y1015 = (add_sel & s1015) | (sub_sel & sub1015) | (and_sel & and1015) | (or_sel & or1015);
  assign y1016 = (add_sel & s1016) | (sub_sel & sub1016) | (and_sel & and1016) | (or_sel & or1016);
  assign y1017 = (add_sel & s1017) | (sub_sel & sub1017) | (and_sel & and1017) | (or_sel & or1017);
  assign y1018 = (add_sel & s1018) | (sub_sel & sub1018) | (and_sel & and1018) | (or_sel & or1018);
  assign y1019 = (add_sel & s1019) | (sub_sel & sub1019) | (and_sel & and1019) | (or_sel & or1019);
  assign y1020 = (add_sel & s1020) | (sub_sel & sub1020) | (and_sel & and1020) | (or_sel & or1020);
  assign y1021 = (add_sel & s1021) | (sub_sel & sub1021) | (and_sel & and1021) | (or_sel & or1021);
  assign y1022 = (add_sel & s1022) | (sub_sel & sub1022) | (and_sel & and1022) | (or_sel & or1022);
  assign y1023 = (add_sel & s1023) | (sub_sel & sub1023) | (and_sel & and1023) | (or_sel & or1023);
endmodule