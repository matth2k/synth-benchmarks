// IWLS benchmark module "example2.blif" printed on Wed May 29 16:34:03 2002
module example2 (a, b, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, \xx , y, z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0, o0, p0, q0, r0, s0, t0, u0, v0, w0, x0, y0, z0, a1, b1, c1, d1, e1, f1, g1, h1, i1, j1, k1, l1, m1, n1, o1, p1, q1, r1, s1, t1, u1, v1, w1, x1, y1, z1, a2, b2, c2, d2, e2, f2, g2, h2, i2, j2, k2, l2, m2, n2, o2, p2, q2, r2, s2, t2, u2, v2, w2, x2, y2, z2, a3, b3, c3, d3, e3, f3, g3, h3, i3, j3, k3, l3, m3, n3, o3, p3, q3, r3, s3, t3, u3, v3, w3, x3, y3, z3, a4, b4, c4, d4, e4, f4, g4, h4, i4, j4, k4, l4, m4, n4, o4, p4, q4, r4, s4, t4, u4, v4);
input
  a,
  b,
  d,
  e,
  f,
  g,
  h,
  i,
  j,
  k,
  l,
  m,
  n,
  o,
  p,
  q,
  r,
  s,
  t,
  u,
  v,
  w,
  \xx ,
  y,
  z,
  a0,
  a1,
  a2,
  b0,
  b1,
  b2,
  c0,
  c1,
  c2,
  d0,
  d1,
  d2,
  e0,
  e1,
  e2,
  f0,
  f1,
  f2,
  g0,
  g1,
  g2,
  h0,
  h1,
  h2,
  i0,
  i1,
  j0,
  j1,
  k0,
  k1,
  l0,
  l1,
  m0,
  m1,
  n0,
  n1,
  o0,
  o1,
  p0,
  p1,
  q0,
  q1,
  r0,
  r1,
  s0,
  s1,
  t0,
  t1,
  u0,
  u1,
  v0,
  v1,
  w0,
  w1,
  x0,
  x1,
  y0,
  y1,
  z0,
  z1;
output
  a3,
  a4,
  b3,
  b4,
  c3,
  c4,
  d3,
  d4,
  e3,
  e4,
  f3,
  f4,
  g3,
  g4,
  h3,
  h4,
  i2,
  i3,
  i4,
  j2,
  j3,
  j4,
  k2,
  k3,
  k4,
  l2,
  l3,
  l4,
  m2,
  m3,
  m4,
  n2,
  n3,
  n4,
  o2,
  o3,
  o4,
  p2,
  p3,
  p4,
  q2,
  q3,
  q4,
  r2,
  r3,
  r4,
  s2,
  s3,
  s4,
  t2,
  t3,
  t4,
  u2,
  u3,
  u4,
  v2,
  v3,
  v4,
  w2,
  w3,
  x2,
  x3,
  y2,
  y3,
  z2,
  z3;
wire
  \[59] ,
  \[15] ,
  \[16] ,
  \[17] ,
  p10,
  \[18] ,
  \[19] ,
  l10,
  \[60] ,
  \[61] ,
  \[62] ,
  \[0] ,
  \[63] ,
  \[1] ,
  \[64] ,
  h10,
  \[20] ,
  \[2] ,
  \[65] ,
  \[21] ,
  \[3] ,
  \[22] ,
  \[4] ,
  \[23] ,
  \[5] ,
  u10,
  \[24] ,
  d10,
  \[6] ,
  \[25] ,
  \[7] ,
  \[26] ,
  \[8] ,
  \[27] ,
  \[9] ,
  q10,
  \[28] ,
  \[29] ,
  m10,
  i10,
  \[30] ,
  \[31] ,
  \[32] ,
  \[33] ,
  v10,
  \[34] ,
  e10,
  \[35] ,
  \[36] ,
  \[37] ,
  r10,
  \[38] ,
  a10,
  \[39] ,
  n10,
  j10,
  \[40] ,
  \[41] ,
  \[42] ,
  \[43] ,
  \[44] ,
  f10,
  \[45] ,
  \[46] ,
  \[47] ,
  s10,
  \[48] ,
  b10,
  \[49] ,
  o10,
  y9,
  z9,
  k10,
  \[50] ,
  \[51] ,
  \[52] ,
  \[53] ,
  \[54] ,
  g10,
  \[10] ,
  \[55] ,
  \[11] ,
  \[56] ,
  \[12] ,
  \[57] ,
  \[13] ,
  t10,
  \[58] ,
  \[14] ,
  c10;
assign
  \[59]  = (n10 & (p0 & (a2 & ~b))) | ((~c2 & (p0 & (a2 & ~b))) | ((l10 & (a2 & ~b)) | (m10 & ~b))),
  \[15]  = (z0 & p0) | (~p0 & i0),
  \[16]  = (y0 & p0) | (~p0 & j0),
  \[17]  = (x0 & p0) | (~p0 & k0),
  p10 = ~a2 & (f & (l10 & (~b & ~b1))),
  \[18]  = (w0 & p0) | (~p0 & l0),
  \[19]  = (v0 & p0) | (~p0 & m0),
  l10 = ~c2 & b2,
  \[60]  = (j10 & (c2 & (~d2 & (d10 & ~b)))) | ((j10 & (c2 & (~e10 & (d10 & ~b)))) | ((k10 & (~d2 & (d10 & ~b))) | ((k10 & (~e10 & (d10 & ~b))) | ((l10 & ~b) | (m10 & ~b))))),
  \[61]  = (k10 & (e10 & (d2 & h10))) | ((j10 & (e10 & (d2 & h10))) | (i10 & (d2 & h10))),
  \[62]  = (f10 & e2) | g10,
  \[0]  = (\[4]  & p0) | ((b1 & p0) | (~p0 & h)),
  \[63]  = f10 & f2,
  \[1]  = (~b2 & (~a2 & ~b)) | ((~c10 & ~b) | (~c2 & ~b)),
  \[64]  = (~a2 & (f & (l10 & ~b))) | (f10 & g2),
  h10 = c2 & ~b,
  \[20]  = (u0 & p0) | (~p0 & n0),
  \[2]  = (k10 & (y1 & h10)) | (j10 & (p1 & h10)),
  \[65]  = f10 & h2,
  \[21]  = (t0 & p0) | (~p0 & o0),
  \[3]  = l10 & (~b & b1),
  \[22]  = (~d10 & (\[2]  & ~q0)) | g10,
  \[4]  = (c10 & ~b) | h10,
  \[23]  = (~c2 & (~f & g)) | (b | ~a),
  \[5]  = (o1 & p0) | (~p0 & y),
  u10 = ~h2 | (g2 | (~f2 | (~e2 | (~d2 | (x1 | ~s0))))),
  \[24]  = (~c10 & (~s0 & (~f & (g & ~b)))) | (~c2 & (~s0 & (~f & (g & ~b)))),
  d10 = (~h2 & e2) | (h2 & ~e2),
  \[6]  = (n1 & p0) | (~p0 & z),
  \[25]  = z9 & g,
  \[7]  = (m1 & p0) | (~p0 & a0),
  \[26]  = z9 & t0,
  \[8]  = (l1 & p0) | (~p0 & b0),
  \[27]  = z9 & u0,
  \[9]  = (k1 & p0) | (~p0 & c0),
  q10 = j10 & (c2 & (~b & ~d10)),
  \[28]  = z9 & v0,
  \[29]  = z9 & w0,
  m10 = (~c2 & ~f) | (n10 & t10),
  i10 = (k10 & ~d10) | ((j10 & ~d10) | (~f & ~c10)),
  \[30]  = z9 & x0,
  \[31]  = z9 & y0,
  \[32]  = z9 & z0,
  \[33]  = (r0 & (b10 & (a10 & g))) | (z9 & a1),
  v10 = ~f2 & ~e2,
  \[34]  = y9 & b1,
  e10 = v10 & (~h2 & ~g2),
  a3 = \[18] ,
  a4 = \[44] ,
  \[35]  = y9 & c1,
  b3 = \[19] ,
  b4 = \[45] ,
  \[36]  = y9 & d1,
  c3 = \[20] ,
  c4 = \[46] ,
  \[37]  = y9 & e1,
  r10 = (f2 & e2) | v10,
  d3 = \[21] ,
  d4 = \[47] ,
  \[38]  = y9 & f1,
  a10 = ~c10 & (~f & h10),
  e3 = \[22] ,
  e4 = \[48] ,
  \[39]  = y9 & g1,
  f3 = \[23] ,
  f4 = \[49] ,
  g3 = \[24] ,
  g4 = \[50] ,
  h3 = \[25] ,
  h4 = \[51] ,
  n10 = b2 & f,
  i2 = \[0] ,
  i3 = \[26] ,
  i4 = \[52] ,
  j2 = \[1] ,
  j3 = \[27] ,
  j4 = \[53] ,
  k2 = \[2] ,
  k3 = \[28] ,
  k4 = \[54] ,
  l2 = \[3] ,
  l3 = \[29] ,
  l4 = \[55] ,
  j10 = ~b2 & a2,
  \[40]  = y9 & h1,
  m2 = \[4] ,
  m3 = \[30] ,
  m4 = \[56] ,
  \[41]  = y9 & i1,
  n2 = \[5] ,
  n3 = \[31] ,
  n4 = \[57] ,
  \[42]  = y9 & j1,
  o2 = \[6] ,
  o3 = \[32] ,
  o4 = \[58] ,
  \[43]  = y9 & k1,
  p2 = \[7] ,
  p3 = \[33] ,
  p4 = \[59] ,
  \[44]  = y9 & l1,
  f10 = h10 & i10,
  q2 = \[8] ,
  q3 = \[34] ,
  q4 = \[60] ,
  \[45]  = y9 & m1,
  r2 = \[9] ,
  r3 = \[35] ,
  r4 = \[61] ,
  \[46]  = y9 & n1,
  s2 = \[10] ,
  s3 = \[36] ,
  s4 = \[62] ,
  \[47]  = (~p1 & (~q0 & (d2 & (d10 & (e10 & (c2 & (~b & j10))))))) | ((p1 & (q0 & (d2 & (d10 & (e10 & (c2 & (~b & j10))))))) | ((y1 & (~d10 & (c2 & (~b & j10)))) | ((q1 & (~d10 & (c2 & (~b & j10)))) | ((q & o10) | (i & p10))))),
  t2 = \[11] ,
  s10 = (~r10 & ~g2) | (r10 & g2),
  t3 = \[37] ,
  t4 = \[63] ,
  \[48]  = (q10 & r1) | ((p10 & j) | (o10 & r)),
  b10 = (~s10 & h2) | (s10 & ~h2),
  u2 = \[12] ,
  u3 = \[38] ,
  u4 = \[64] ,
  \[49]  = (q10 & s1) | ((p10 & k) | (o10 & s)),
  v2 = \[13] ,
  v3 = \[39] ,
  v4 = \[65] ,
  w2 = \[14] ,
  w3 = \[40] ,
  x2 = \[15] ,
  x3 = \[41] ,
  o10 = ~a2 & (f & \[3] ),
  y2 = \[16] ,
  y3 = \[42] ,
  y9 = (r0 & (b10 & a10)) | z9,
  z2 = \[17] ,
  z3 = \[43] ,
  z9 = (~r10 & (~h2 & (~r0 & a10))) | (r10 & (h2 & (~r0 & a10))),
  k10 = b2 & ~a2,
  \[50]  = (q10 & t1) | ((p10 & l) | (o10 & t)),
  \[51]  = (q10 & u1) | ((p10 & m) | (o10 & u)),
  \[52]  = (q10 & v1) | ((p10 & n) | (o10 & v)),
  \[53]  = (q10 & w1) | ((p10 & o) | (o10 & w)),
  \[54]  = (p10 & p) | (o10 & \xx ),
  g10 = (t10 & (~b & n10)) | (~c2 & (~b & n10)),
  \[10]  = (j1 & p0) | (~p0 & d0),
  \[55]  = v10 & (a10 & (h2 & (g2 & ~d2))),
  \[11]  = (i1 & p0) | (~p0 & e0),
  \[56]  = (~y1 & (~q0 & (d10 & (c2 & ~a2)))) | ((y1 & (q0 & (d10 & (c2 & ~a2)))) | ((~e10 & (d10 & (c10 & c2))) | ((~d2 & (d10 & (c10 & c2))) | ((z1 & (~d10 & (c10 & c2))) | ((~b2 & ~a2) | (~a | b)))))),
  \[12]  = (h1 & p0) | (~p0 & f0),
  \[57]  = e & (~d & (~b & a)),
  \[13]  = (g1 & p0) | (~p0 & g0),
  t10 = u10 & (a2 & ~r0),
  \[58]  = (~u10 & (~r0 & (a2 & (h10 & n10)))) | ((j10 & (~r0 & (p0 & (~c2 & ~b)))) | ((r0 & (~p0 & (a2 & (h10 & n10)))) | ((k10 & (~c2 & ~b)) | (~f & (~c2 & ~b))))),
  \[14]  = (a1 & p0) | (~p0 & h0),
  c10 = ~b2 | ~a2;
endmodule

