// IWLS benchmark module "cu" printed on Wed May 29 16:31:30 2002
module cu(a, b, c, d, e, f, g, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, \xx , y, z);
input
  a,
  b,
  c,
  d,
  e,
  f,
  g,
  i,
  j,
  k,
  l,
  m,
  n,
  o;
output
  p,
  q,
  r,
  s,
  t,
  u,
  v,
  w,
  \xx ,
  y,
  z;
wire
  o0,
  p0,
  \[0] ,
  a1,
  t0,
  \[1] ,
  b1,
  \[2] ,
  \[3] ,
  \[4] ,
  x0,
  \[5] ,
  f1,
  y0,
  \[6] ,
  g1,
  z0,
  \[7] ,
  \[8] ,
  \[10] ,
  i1,
  \[9] ,
  j1;
assign
  o0 = (~f & ~e) | ((~f & ~c) | ((f & e) | ((f & c) | ((~e & c) | (e & ~c))))),
  p0 = ~o0 & ~d,
  p = \[0] ,
  q = \[1] ,
  r = \[2] ,
  s = \[3] ,
  t = \[4] ,
  u = \[5] ,
  v = \[6] ,
  w = \[7] ,
  \xx  = \[8] ,
  y = \[9] ,
  z = \[10] ,
  \[0]  = ~p0,
  a1 = (l & (b & ~a)) | ((m & (b & a)) | ((k & (~b & a)) | ~f1)),
  t0 = a | (b | (c | d)),
  \[1]  = ~o0 & ~d,
  b1 = (c & f) | ((c & o) | (d | ~e)),
  \[2]  = ~t0 & (~e & (f & ~o)),
  \[3]  = ~x0 & (~e & (f & ~o)),
  \[4]  = ~y0 & (~e & (f & ~o)),
  x0 = ~a | (b | (c | d)),
  \[5]  = ~z0 & (~e & (f & ~o)),
  f1 = ~g1 & ~i,
  y0 = a | (~b | (c | d)),
  \[6]  = (~b1 & ~a1) | (~b1 & c),
  g1 = (j & (~b & ~a)) | (~o | (~f | n)),
  z0 = ~a | (~b | (c | d)),
  \[7]  = ~i1 & ~o,
  \[8]  = (~b1 & ~j1) | (~b1 & c),
  \[10]  = (g & (~d & ~f)) | (g & (~d & ~c)),
  i1 = c | (d | (e | ~f)),
  \[9]  = g & o,
  j1 = ~f | (n | ~o);
endmodule

