module s9234 (
  CK,
  g102,
  g107,
  g22,
  g23,
  g301,
  g306,
  g310,
  g314,
  g319,
  g32,
  g36,
  g37,
  g38,
  g39,
  g40,
  g41,
  g42,
  g44,
  g45,
  g46,
  g47,
  g557,
  g558,
  g559,
  g560,
  g561,
  g562,
  g563,
  g564,
  g567,
  g639,
  g702,
  g705,
  g89,
  g94,
  g98,
  g4100,
  g2584,
  g4108,
  g6374,
  g5692,
  g6728,
  g6372,
  g4109,
  g4105,
  g4809,
  g3222,
  g3600,
  g5137,
  g1293,
  g1290,
  g4104,
  g6370,
  g4107,
  g4422,
  g4099,
  g6362,
  g4098,
  g6360,
  g6364,
  g4106,
  g4103,
  g4321,
  g5469,
  g6368,
  g6282,
  g6284,
  g4101,
  g6366,
  g4112,
  g4307,
  g5468,
  g4121,
  g4102,
  g4110
);
  input CK;
  wire CK;
  input g102;
  wire g102;
  input g107;
  wire g107;
  input g22;
  wire g22;
  input g23;
  wire g23;
  input g301;
  wire g301;
  input g306;
  wire g306;
  input g310;
  wire g310;
  input g314;
  wire g314;
  input g319;
  wire g319;
  input g32;
  wire g32;
  input g36;
  wire g36;
  input g37;
  wire g37;
  input g38;
  wire g38;
  input g39;
  wire g39;
  input g40;
  wire g40;
  input g41;
  wire g41;
  input g42;
  wire g42;
  input g44;
  wire g44;
  input g45;
  wire g45;
  input g46;
  wire g46;
  input g47;
  wire g47;
  input g557;
  wire g557;
  input g558;
  wire g558;
  input g559;
  wire g559;
  input g560;
  wire g560;
  input g561;
  wire g561;
  input g562;
  wire g562;
  input g563;
  wire g563;
  input g564;
  wire g564;
  input g567;
  wire g567;
  input g639;
  wire g639;
  input g702;
  wire g702;
  input g705;
  wire g705;
  input g89;
  wire g89;
  input g94;
  wire g94;
  input g98;
  wire g98;
  output g4100;
  wire g4100;
  output g2584;
  wire g2584;
  output g4108;
  wire g4108;
  output g6374;
  wire g6374;
  output g5692;
  wire g5692;
  output g6728;
  wire g6728;
  output g6372;
  wire g6372;
  output g4109;
  wire g4109;
  output g4105;
  wire g4105;
  output g4809;
  wire g4809;
  output g3222;
  wire g3222;
  output g3600;
  wire g3600;
  output g5137;
  wire g5137;
  output g1293;
  wire g1293;
  output g1290;
  wire g1290;
  output g4104;
  wire g4104;
  output g6370;
  wire g6370;
  output g4107;
  wire g4107;
  output g4422;
  wire g4422;
  output g4099;
  wire g4099;
  output g6362;
  wire g6362;
  output g4098;
  wire g4098;
  output g6360;
  wire g6360;
  output g6364;
  wire g6364;
  output g4106;
  wire g4106;
  output g4103;
  wire g4103;
  output g4321;
  wire g4321;
  output g5469;
  wire g5469;
  output g6368;
  wire g6368;
  output g6282;
  wire g6282;
  output g6284;
  wire g6284;
  output g4101;
  wire g4101;
  output g6366;
  wire g6366;
  output g4112;
  wire g4112;
  output g4307;
  wire g4307;
  output g5468;
  wire g5468;
  output g4121;
  wire g4121;
  output g4102;
  wire g4102;
  output g4110;
  wire g4110;
  wire __0__;
  wire __1__;
  wire __2__;
  wire __3__;
  wire __4__;
  wire __5__;
  wire __6__;
  wire __7__;
  wire __8__;
  wire __9__;
  wire __10__;
  wire __11__;
  wire __12__;
  wire __13__;
  wire __14__;
  wire __15__;
  wire __16__;
  wire __17__;
  wire __18__;
  wire __19__;
  wire __20__;
  wire __21__;
  wire __22__;
  wire __23__;
  wire __24__;
  wire __25__;
  wire __26__;
  wire __27__;
  wire __28__;
  wire __29__;
  wire __30__;
  wire __31__;
  wire __32__;
  wire __33__;
  wire __34__;
  wire __35__;
  wire __36__;
  wire __37__;
  wire __38__;
  wire __39__;
  wire __40__;
  wire __41__;
  wire __42__;
  wire __43__;
  wire __44__;
  wire __45__;
  wire __46__;
  wire __47__;
  wire __48__;
  wire __49__;
  wire __50__;
  wire __51__;
  wire __52__;
  wire __53__;
  wire __54__;
  wire __55__;
  wire __56__;
  wire __57__;
  wire __58__;
  wire __59__;
  wire __60__;
  wire __61__;
  wire __62__;
  wire __63__;
  wire __64__;
  wire __65__;
  wire __66__;
  wire __67__;
  wire __68__;
  wire __69__;
  wire __70__;
  wire __71__;
  wire __72__;
  wire __73__;
  wire __74__;
  wire __75__;
  wire __76__;
  wire __77__;
  wire __78__;
  wire __79__;
  wire __80__;
  wire __81__;
  wire __82__;
  wire __83__;
  wire __84__;
  wire __85__;
  wire __86__;
  wire __87__;
  wire __88__;
  wire __89__;
  wire __90__;
  wire __91__;
  wire __92__;
  wire __93__;
  wire __94__;
  wire __95__;
  wire __96__;
  wire __97__;
  wire __98__;
  wire __99__;
  wire __100__;
  wire __101__;
  wire __102__;
  wire __103__;
  wire __104__;
  wire __105__;
  wire __106__;
  wire __107__;
  wire __108__;
  wire __109__;
  wire __110__;
  wire __111__;
  wire __112__;
  wire __113__;
  wire __114__;
  wire __115__;
  wire __116__;
  wire __117__;
  wire __118__;
  wire __119__;
  wire __120__;
  wire __121__;
  wire __122__;
  wire __123__;
  wire __124__;
  wire __125__;
  wire __126__;
  wire __127__;
  wire __128__;
  wire __129__;
  wire __130__;
  wire __131__;
  wire __132__;
  wire __133__;
  wire __134__;
  wire __135__;
  wire __136__;
  wire __137__;
  wire __138__;
  wire __139__;
  wire __140__;
  wire __142__;
  wire __143__;
  wire __144__;
  wire __145__;
  wire __146__;
  wire __147__;
  wire __148__;
  wire __149__;
  wire __151__;
  wire __152__;
  wire __153__;
  wire __154__;
  wire __155__;
  wire __156__;
  wire __157__;
  wire __158__;
  wire __159__;
  wire __160__;
  wire __161__;
  wire __162__;
  wire __163__;
  wire __164__;
  wire __165__;
  wire __166__;
  wire __167__;
  wire __168__;
  wire __169__;
  wire __170__;
  wire __171__;
  wire __172__;
  wire __173__;
  wire __174__;
  wire __175__;
  wire __176__;
  wire __177__;
  wire __178__;
  wire __179__;
  wire __180__;
  wire __181__;
  wire __182__;
  wire __183__;
  wire __184__;
  wire __185__;
  wire __186__;
  wire __187__;
  wire __188__;
  wire __189__;
  wire __190__;
  wire __191__;
  wire __192__;
  wire __193__;
  wire __194__;
  wire __195__;
  wire __196__;
  wire __197__;
  wire __198__;
  wire __199__;
  wire __200__;
  wire __201__;
  wire __202__;
  wire __203__;
  wire __204__;
  wire __205__;
  wire __206__;
  wire __207__;
  wire __208__;
  wire __209__;
  wire __210__;
  wire __211__;
  wire __212__;
  wire __213__;
  wire __214__;
  wire __215__;
  wire __216__;
  wire __217__;
  wire __218__;
  wire __219__;
  wire __220__;
  wire __221__;
  wire __222__;
  wire __223__;
  wire __224__;
  wire __225__;
  wire __226__;
  wire __227__;
  wire __228__;
  wire __229__;
  wire __230__;
  wire __231__;
  wire __232__;
  wire __233__;
  wire __234__;
  wire __235__;
  wire __236__;
  wire __237__;
  wire __238__;
  wire __239__;
  wire __240__;
  wire __241__;
  wire __242__;
  wire __243__;
  wire __244__;
  wire __245__;
  wire __246__;
  wire __247__;
  wire __248__;
  wire __249__;
  wire __250__;
  wire __251__;
  wire __252__;
  wire __253__;
  wire __254__;
  wire __255__;
  wire __256__;
  wire __257__;
  wire __258__;
  wire __259__;
  wire __260__;
  wire __261__;
  wire __262__;
  wire __263__;
  wire __264__;
  wire __265__;
  wire __266__;
  wire __267__;
  wire __268__;
  wire __269__;
  wire __270__;
  wire __271__;
  wire __272__;
  wire __273__;
  wire __274__;
  wire __275__;
  wire __276__;
  wire __277__;
  wire __278__;
  wire __279__;
  wire __280__;
  wire __281__;
  wire __282__;
  wire __283__;
  wire __284__;
  wire __285__;
  wire __286__;
  wire __287__;
  wire __288__;
  wire __289__;
  wire __290__;
  wire __291__;
  wire __292__;
  wire __293__;
  wire __294__;
  wire __295__;
  wire __296__;
  wire __297__;
  wire __298__;
  wire __299__;
  wire __300__;
  wire __301__;
  wire __302__;
  wire __303__;
  wire __304__;
  wire __305__;
  wire __306__;
  wire __307__;
  wire __308__;
  wire __309__;
  wire __310__;
  wire __311__;
  wire __312__;
  wire __313__;
  wire __314__;
  wire __315__;
  wire __316__;
  wire __317__;
  wire __318__;
  wire __319__;
  wire __320__;
  wire __321__;
  wire __322__;
  wire __323__;
  wire __324__;
  wire __325__;
  wire __326__;
  wire __327__;
  wire __328__;
  wire __329__;
  wire __330__;
  wire __331__;
  wire __332__;
  wire __333__;
  wire __334__;
  wire __335__;
  wire __336__;
  wire __337__;
  wire __338__;
  wire __339__;
  wire __340__;
  wire __341__;
  wire __342__;
  wire __343__;
  wire __344__;
  wire __345__;
  wire __346__;
  wire __347__;
  wire __348__;
  wire __349__;
  wire __350__;
  wire __351__;
  wire __352__;
  wire __353__;
  wire __354__;
  wire __355__;
  wire __356__;
  wire __357__;
  wire __358__;
  wire __359__;
  wire __360__;
  wire __361__;
  wire __362__;
  wire __363__;
  wire __364__;
  wire __365__;
  wire __366__;
  wire __367__;
  wire __368__;
  wire __369__;
  wire __370__;
  wire __371__;
  INV __372__ (
    .I(__1__),
    .O(__0__)
  );
  LUT4 #(
    .INIT(16'he0ff)
  ) __373__ (
    .I3(__120__),
    .I2(__16__),
    .I1(__60__),
    .I0(__139__),
    .O(__1__)
  );
  INV __374__ (
    .I(__115__),
    .O(__2__)
  );
  INV __375__ (
    .I(__135__),
    .O(__3__)
  );
  INV __376__ (
    .I(g47),
    .O(__4__)
  );
  INV __377__ (
    .I(__109__),
    .O(__5__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __378__ (
    .D(__15__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__6__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __379__ (
    .D(__228__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__7__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __380__ (
    .D(__275__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__8__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __381__ (
    .D(__117__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__9__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __382__ (
    .D(__63__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__10__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __383__ (
    .D(__293__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__11__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __384__ (
    .D(g37),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__12__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __385__ (
    .D(__284__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__13__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __386__ (
    .D(__321__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__14__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __387__ (
    .D(__292__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__15__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __388__ (
    .D(g40),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__16__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __389__ (
    .D(__130__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__17__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __390__ (
    .D(__3__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__18__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __391__ (
    .D(__347__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__19__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __392__ (
    .D(__336__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__20__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __393__ (
    .D(__137__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__21__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __394__ (
    .D(__371__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__22__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __395__ (
    .D(__327__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__23__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __396__ (
    .D(__270__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__24__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __397__ (
    .D(__369__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__25__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __398__ (
    .D(__265__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__26__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __399__ (
    .D(__309__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__27__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __400__ (
    .D(__255__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__28__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __401__ (
    .D(__349__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__29__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __402__ (
    .D(__264__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__30__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __403__ (
    .D(__43__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__31__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __404__ (
    .D(__224__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__32__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __405__ (
    .D(g702),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__33__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __406__ (
    .D(__5__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__34__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __407__ (
    .D(__208__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__35__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __408__ (
    .D(__258__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__36__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __409__ (
    .D(__279__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__37__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __410__ (
    .D(__276__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__38__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __411__ (
    .D(__236__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__39__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __412__ (
    .D(__85__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__40__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __413__ (
    .D(g46),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__41__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __414__ (
    .D(__335__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__42__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __415__ (
    .D(__110__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__43__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __416__ (
    .D(__199__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__44__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __417__ (
    .D(__339__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__45__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __418__ (
    .D(__325__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__46__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __419__ (
    .D(__92__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__47__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __420__ (
    .D(__2__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__48__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __421__ (
    .D(__290__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__49__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __422__ (
    .D(__307__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__50__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __423__ (
    .D(__239__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__51__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __424__ (
    .D(__334__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__52__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __425__ (
    .D(__149__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__53__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __426__ (
    .D(__338__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__54__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __427__ (
    .D(__345__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__55__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __428__ (
    .D(__17__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__56__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __429__ (
    .D(__319__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__57__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __430__ (
    .D(__207__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__58__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __431__ (
    .D(__252__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__59__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __432__ (
    .D(g32),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__60__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __433__ (
    .D(__44__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__61__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __434__ (
    .D(__201__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__62__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __435__ (
    .D(__303__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__63__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __436__ (
    .D(__253__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__64__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __437__ (
    .D(__333__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__65__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __438__ (
    .D(__329__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__66__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __439__ (
    .D(__360__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__67__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __440__ (
    .D(__32__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__68__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __441__ (
    .D(__285__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__69__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __442__ (
    .D(__316__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__70__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __443__ (
    .D(__230__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__71__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __444__ (
    .D(__242__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__72__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __445__ (
    .D(__121__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__73__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __446__ (
    .D(__164__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__74__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __447__ (
    .D(__259__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__75__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __448__ (
    .D(__361__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__76__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __449__ (
    .D(__323__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__77__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __450__ (
    .D(__337__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__78__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __451__ (
    .D(__288__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__79__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __452__ (
    .D(__134__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__80__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __453__ (
    .D(__344__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__81__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __454__ (
    .D(__314__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__82__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __455__ (
    .D(__328__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__83__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __456__ (
    .D(__322__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__84__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __457__ (
    .D(__94__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__85__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __458__ (
    .D(__128__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__86__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __459__ (
    .D(__286__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__87__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __460__ (
    .D(__266__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__88__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __461__ (
    .D(__257__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__89__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __462__ (
    .D(__312__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__90__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __463__ (
    .D(__268__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__91__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __464__ (
    .D(__267__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__92__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __465__ (
    .D(__244__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__93__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __466__ (
    .D(__198__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__94__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __467__ (
    .D(__125__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__95__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __468__ (
    .D(__269__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__96__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __469__ (
    .D(__232__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__97__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __470__ (
    .D(__320__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__98__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __471__ (
    .D(__282__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__99__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __472__ (
    .D(__249__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__100__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __473__ (
    .D(__332__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__101__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __474__ (
    .D(__211__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__102__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __475__ (
    .D(__326__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__103__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __476__ (
    .D(__203__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__104__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __477__ (
    .D(__126__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__105__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __478__ (
    .D(__263__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__106__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __479__ (
    .D(__313__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__107__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __480__ (
    .D(__206__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__108__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __481__ (
    .D(__10__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__109__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __482__ (
    .D(g42),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__110__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __483__ (
    .D(__346__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__111__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __484__ (
    .D(__273__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__112__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __485__ (
    .D(g567),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__113__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __486__ (
    .D(__304__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__114__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __487__ (
    .D(__289__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__115__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __488__ (
    .D(__89__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__116__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __489__ (
    .D(__107__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__117__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __490__ (
    .D(__65__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__118__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __491__ (
    .D(__283__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__119__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __492__ (
    .D(g39),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__120__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __493__ (
    .D(__370__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__121__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __494__ (
    .D(__62__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__122__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __495__ (
    .D(__234__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__123__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __496__ (
    .D(__260__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__124__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __497__ (
    .D(__72__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__125__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __498__ (
    .D(__356__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__126__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __499__ (
    .D(__363__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__127__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __500__ (
    .D(__261__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__128__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __501__ (
    .D(__318__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__129__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __502__ (
    .D(__343__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__130__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __503__ (
    .D(__324__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__131__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __504__ (
    .D(__200__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__132__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __505__ (
    .D(__4__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__133__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __506__ (
    .D(__25__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__134__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __507__ (
    .D(__68__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__135__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __508__ (
    .D(__105__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__136__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __509__ (
    .D(g45),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__137__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __510__ (
    .D(__308__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__138__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __511__ (
    .D(g38),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__139__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __512__ (
    .D(__350__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__140__)
  );
  LUT6 #(
    .INIT(64'h00007fffffff0000)
  ) __514__ (
    .I5(__39__),
    .I4(__104__),
    .I3(__54__),
    .I2(__64__),
    .I1(__93__),
    .I0(__103__),
    .O(__142__)
  );
  LUT6 #(
    .INIT(64'hccccaaaaff00f0f0)
  ) __515__ (
    .I5(__54__),
    .I4(__64__),
    .I3(__40__),
    .I2(__136__),
    .I1(__109__),
    .I0(__135__),
    .O(__143__)
  );
  LUT6 #(
    .INIT(64'hccccaaaaff00f0f0)
  ) __516__ (
    .I5(__54__),
    .I4(__64__),
    .I3(__9__),
    .I2(__80__),
    .I1(__56__),
    .I0(__95__),
    .O(__144__)
  );
  LUT2 #(
    .INIT(4'h9)
  ) __517__ (
    .I1(__39__),
    .I0(__104__),
    .O(__145__)
  );
  LUT6 #(
    .INIT(64'h33cc0ff055aa55aa)
  ) __518__ (
    .I5(__145__),
    .I4(__103__),
    .I3(__43__),
    .I2(__144__),
    .I1(__143__),
    .I0(__142__),
    .O(__146__)
  );
  LUT6 #(
    .INIT(64'h8000000000000000)
  ) __519__ (
    .I5(__39__),
    .I4(__104__),
    .I3(__54__),
    .I2(__64__),
    .I1(__93__),
    .I0(__103__),
    .O(__147__)
  );
  LUT5 #(
    .INIT(32'h00ff0efe)
  ) __520__ (
    .I4(__69__),
    .I3(__147__),
    .I2(__53__),
    .I1(__43__),
    .I0(__142__),
    .O(__148__)
  );
  LUT5 #(
    .INIT(32'h44fff0f0)
  ) __521__ (
    .I4(__23__),
    .I3(__148__),
    .I2(__9__),
    .I1(__53__),
    .I0(__146__),
    .O(__149__)
  );
  LUT6 #(
    .INIT(64'h8000000000000000)
  ) __523__ (
    .I5(__51__),
    .I4(__77__),
    .I3(__87__),
    .I2(__129__),
    .I1(__49__),
    .I0(__131__),
    .O(__151__)
  );
  LUT6 #(
    .INIT(64'hb00b00000000b00b)
  ) __524__ (
    .I5(__86__),
    .I4(__11__),
    .I3(__118__),
    .I2(__96__),
    .I1(__14__),
    .I0(__73__),
    .O(__152__)
  );
  LUT2 #(
    .INIT(4'h9)
  ) __525__ (
    .I1(__61__),
    .I0(__132__),
    .O(__153__)
  );
  LUT4 #(
    .INIT(16'h9009)
  ) __526__ (
    .I3(__47__),
    .I2(__124__),
    .I1(__113__),
    .I0(__50__),
    .O(__154__)
  );
  LUT6 #(
    .INIT(64'h9009000000000000)
  ) __527__ (
    .I5(__154__),
    .I4(__153__),
    .I3(__116__),
    .I2(__76__),
    .I1(__122__),
    .I0(__91__),
    .O(__155__)
  );
  LUT6 #(
    .INIT(64'hb00b000000000000)
  ) __528__ (
    .I5(__155__),
    .I4(__152__),
    .I3(__46__),
    .I2(__6__),
    .I1(__73__),
    .I0(__14__),
    .O(__156__)
  );
  LUT6 #(
    .INIT(64'h0f050f030f0f0f0f)
  ) __529__ (
    .I5(__156__),
    .I4(__111__),
    .I3(__7__),
    .I2(__74__),
    .I1(__151__),
    .I0(__147__),
    .O(__157__)
  );
  LUT5 #(
    .INIT(32'h00004000)
  ) __530__ (
    .I4(__95__),
    .I3(__60__),
    .I2(__120__),
    .I1(__16__),
    .I0(__139__),
    .O(__158__)
  );
  LUT4 #(
    .INIT(16'h4000)
  ) __531__ (
    .I3(__9__),
    .I2(__80__),
    .I1(__158__),
    .I0(__56__),
    .O(__159__)
  );
  LUT4 #(
    .INIT(16'h9669)
  ) __532__ (
    .I3(__105__),
    .I2(__85__),
    .I1(__10__),
    .I0(__68__),
    .O(__160__)
  );
  LUT4 #(
    .INIT(16'h9669)
  ) __533__ (
    .I3(__17__),
    .I2(__125__),
    .I1(__134__),
    .I0(__117__),
    .O(__161__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __534__ (
    .I1(g702),
    .I0(__133__),
    .O(__162__)
  );
  LUT6 #(
    .INIT(64'hebbe000000000000)
  ) __535__ (
    .I5(__108__),
    .I4(__162__),
    .I3(__99__),
    .I2(__161__),
    .I1(__160__),
    .I0(g41),
    .O(__163__)
  );
  LUT6 #(
    .INIT(64'h555555555555d515)
  ) __536__ (
    .I5(__109__),
    .I4(g41),
    .I3(__136__),
    .I2(__163__),
    .I1(__159__),
    .I0(__157__),
    .O(__164__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __537__ (
    .I1(__87__),
    .I0(__131__),
    .O(__165__)
  );
  LUT4 #(
    .INIT(16'h8000)
  ) __538__ (
    .I3(__87__),
    .I2(__129__),
    .I1(__49__),
    .I0(__131__),
    .O(__166__)
  );
  LUT6 #(
    .INIT(64'h5555fffefffcffff)
  ) __539__ (
    .I5(__51__),
    .I4(__77__),
    .I3(__90__),
    .I2(__114__),
    .I1(__31__),
    .I0(__166__),
    .O(__167__)
  );
  LUT6 #(
    .INIT(64'h00007fffffff0000)
  ) __540__ (
    .I5(__51__),
    .I4(__77__),
    .I3(__87__),
    .I2(__129__),
    .I1(__49__),
    .I0(__131__),
    .O(__168__)
  );
  LUT5 #(
    .INIT(32'haaaaaaa8)
  ) __541__ (
    .I4(__90__),
    .I3(__114__),
    .I2(__31__),
    .I1(__168__),
    .I0(__167__),
    .O(__169__)
  );
  LUT4 #(
    .INIT(16'h0001)
  ) __542__ (
    .I3(__120__),
    .I2(__16__),
    .I1(__139__),
    .I0(__12__),
    .O(__170__)
  );
  LUT6 #(
    .INIT(64'h3c00aaaa00000000)
  ) __543__ (
    .I5(__170__),
    .I4(__55__),
    .I3(__169__),
    .I2(__49__),
    .I1(__165__),
    .I0(__40__),
    .O(__171__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __544__ (
    .I1(__54__),
    .I0(__64__),
    .O(__172__)
  );
  LUT4 #(
    .INIT(16'h8000)
  ) __545__ (
    .I3(__54__),
    .I2(__64__),
    .I1(__93__),
    .I0(__103__),
    .O(__173__)
  );
  LUT6 #(
    .INIT(64'h5555fffefffcffff)
  ) __546__ (
    .I5(__39__),
    .I4(__104__),
    .I3(__69__),
    .I2(__53__),
    .I1(__43__),
    .I0(__173__),
    .O(__174__)
  );
  LUT5 #(
    .INIT(32'haaaaaaa8)
  ) __547__ (
    .I4(__69__),
    .I3(__53__),
    .I2(__43__),
    .I1(__142__),
    .I0(__174__),
    .O(__175__)
  );
  LUT3 #(
    .INIT(8'h08)
  ) __548__ (
    .I2(__88__),
    .I1(g41),
    .I0(__48__),
    .O(__176__)
  );
  LUT5 #(
    .INIT(32'h00000008)
  ) __549__ (
    .I4(__120__),
    .I3(__16__),
    .I2(__139__),
    .I1(__12__),
    .I0(__176__),
    .O(__177__)
  );
  LUT6 #(
    .INIT(64'h3c00aaaa00000000)
  ) __550__ (
    .I5(__177__),
    .I4(__23__),
    .I3(__175__),
    .I2(__103__),
    .I1(__172__),
    .I0(__40__),
    .O(__178__)
  );
  LUT3 #(
    .INIT(8'h01)
  ) __551__ (
    .I2(__120__),
    .I1(__16__),
    .I0(__139__),
    .O(__179__)
  );
  LUT4 #(
    .INIT(16'he0ff)
  ) __552__ (
    .I3(__120__),
    .I2(__16__),
    .I1(__60__),
    .I0(__139__),
    .O(__180__)
  );
  LUT6 #(
    .INIT(64'h0e00000000000000)
  ) __553__ (
    .I5(g702),
    .I4(__133__),
    .I3(g41),
    .I2(__88__),
    .I1(__115__),
    .I0(__48__),
    .O(__181__)
  );
  LUT6 #(
    .INIT(64'hbfffffffffffffff)
  ) __554__ (
    .I5(__80__),
    .I4(__181__),
    .I3(__60__),
    .I2(__120__),
    .I1(__16__),
    .I0(__139__),
    .O(__182__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __555__ (
    .I2(__120__),
    .I1(__16__),
    .I0(__139__),
    .O(__183__)
  );
  LUT5 #(
    .INIT(32'hcaffffff)
  ) __556__ (
    .I4(__181__),
    .I3(__183__),
    .I2(__135__),
    .I1(__136__),
    .I0(__40__),
    .O(__184__)
  );
  LUT6 #(
    .INIT(64'h4fff000000000000)
  ) __557__ (
    .I5(__184__),
    .I4(__182__),
    .I3(__163__),
    .I2(__176__),
    .I1(__180__),
    .I0(__179__),
    .O(__185__)
  );
  LUT4 #(
    .INIT(16'h4000)
  ) __558__ (
    .I3(__60__),
    .I2(__120__),
    .I1(__16__),
    .I0(__139__),
    .O(__186__)
  );
  LUT6 #(
    .INIT(64'h0000000080000000)
  ) __559__ (
    .I5(__109__),
    .I4(__95__),
    .I3(__9__),
    .I2(__80__),
    .I1(__181__),
    .I0(__186__),
    .O(__187__)
  );
  LUT6 #(
    .INIT(64'h8000000000000000)
  ) __560__ (
    .I5(__109__),
    .I4(__95__),
    .I3(__9__),
    .I2(__80__),
    .I1(__181__),
    .I0(__186__),
    .O(__188__)
  );
  LUT5 #(
    .INIT(32'h80000000)
  ) __561__ (
    .I4(__9__),
    .I3(__80__),
    .I2(__181__),
    .I1(__158__),
    .I0(__56__),
    .O(__189__)
  );
  LUT6 #(
    .INIT(64'h0000000000008000)
  ) __562__ (
    .I5(__9__),
    .I4(__139__),
    .I3(__80__),
    .I2(__60__),
    .I1(__120__),
    .I0(__16__),
    .O(__190__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __563__ (
    .I1(__181__),
    .I0(__190__),
    .O(__191__)
  );
  LUT5 #(
    .INIT(32'h00008000)
  ) __564__ (
    .I4(__136__),
    .I3(__181__),
    .I2(__40__),
    .I1(__135__),
    .I0(__183__),
    .O(__192__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __565__ (
    .I5(__192__),
    .I4(g562),
    .I3(__191__),
    .I2(__123__),
    .I1(__189__),
    .I0(__97__),
    .O(__193__)
  );
  LUT6 #(
    .INIT(64'h0000000000008000)
  ) __566__ (
    .I5(__109__),
    .I4(__56__),
    .I3(__9__),
    .I2(__80__),
    .I1(__181__),
    .I0(__158__),
    .O(__194__)
  );
  LUT6 #(
    .INIT(64'h0000000080000000)
  ) __567__ (
    .I5(__56__),
    .I4(__109__),
    .I3(__9__),
    .I2(__80__),
    .I1(__181__),
    .I0(__158__),
    .O(__195__)
  );
  LUT4 #(
    .INIT(16'h0777)
  ) __568__ (
    .I3(__195__),
    .I2(__132__),
    .I1(__7__),
    .I0(__194__),
    .O(__196__)
  );
  LUT6 #(
    .INIT(64'h153f000000000000)
  ) __569__ (
    .I5(__196__),
    .I4(__193__),
    .I3(__188__),
    .I2(__187__),
    .I1(__24__),
    .I0(__78__),
    .O(__197__)
  );
  LUT6 #(
    .INIT(64'hfffffff8ffffffff)
  ) __570__ (
    .I5(__197__),
    .I4(__185__),
    .I3(__178__),
    .I2(__171__),
    .I1(__40__),
    .I0(__0__),
    .O(__198__)
  );
  LUT4 #(
    .INIT(16'h7800)
  ) __571__ (
    .I3(__21__),
    .I2(__44__),
    .I1(__128__),
    .I0(g567),
    .O(__199__)
  );
  LUT6 #(
    .INIT(64'hccccec4ccccccccc)
  ) __572__ (
    .I5(__109__),
    .I4(g41),
    .I3(__40__),
    .I2(__163__),
    .I1(__132__),
    .I0(__159__),
    .O(__200__)
  );
  LUT5 #(
    .INIT(32'h6ccc0000)
  ) __573__ (
    .I4(__21__),
    .I3(__44__),
    .I2(__128__),
    .I1(__62__),
    .I0(g567),
    .O(__201__)
  );
  LUT4 #(
    .INIT(16'h0001)
  ) __574__ (
    .I3(__69__),
    .I2(__53__),
    .I1(__43__),
    .I0(__142__),
    .O(__202__)
  );
  LUT6 #(
    .INIT(64'hdffdffffdffd0000)
  ) __575__ (
    .I5(__56__),
    .I4(__23__),
    .I3(__104__),
    .I2(__173__),
    .I1(__202__),
    .I0(__174__),
    .O(__203__)
  );
  LUT6 #(
    .INIT(64'h9669699669969669)
  ) __576__ (
    .I5(g40),
    .I4(g38),
    .I3(g37),
    .I2(g39),
    .I1(g32),
    .I0(g36),
    .O(__204__)
  );
  LUT6 #(
    .INIT(64'h9669699669969669)
  ) __577__ (
    .I5(__99__),
    .I4(__161__),
    .I3(__105__),
    .I2(__85__),
    .I1(__10__),
    .I0(__68__),
    .O(__205__)
  );
  LUT2 #(
    .INIT(4'h9)
  ) __578__ (
    .I1(__205__),
    .I0(__204__),
    .O(__206__)
  );
  LUT5 #(
    .INIT(32'haaacaaaa)
  ) __579__ (
    .I4(__156__),
    .I3(__7__),
    .I2(__74__),
    .I1(__66__),
    .I0(__58__),
    .O(__207__)
  );
  LUT5 #(
    .INIT(32'haaacaaaa)
  ) __580__ (
    .I4(__156__),
    .I3(__7__),
    .I2(__74__),
    .I1(__127__),
    .I0(__35__),
    .O(__208__)
  );
  LUT6 #(
    .INIT(64'hfaffffffffffffff)
  ) __581__ (
    .I5(g41),
    .I4(__108__),
    .I3(__33__),
    .I2(g22),
    .I1(__205__),
    .I0(__126__),
    .O(__209__)
  );
  LUT6 #(
    .INIT(64'hfaffffffffffffff)
  ) __582__ (
    .I5(g41),
    .I4(__108__),
    .I3(__33__),
    .I2(g22),
    .I1(__205__),
    .I0(__72__),
    .O(__210__)
  );
  LUT5 #(
    .INIT(32'haaaaea2a)
  ) __583__ (
    .I4(g41),
    .I3(__136__),
    .I2(__163__),
    .I1(__190__),
    .I0(__102__),
    .O(__211__)
  );
  LUT6 #(
    .INIT(64'h3c00aaaa00000000)
  ) __584__ (
    .I5(__177__),
    .I4(__23__),
    .I3(__175__),
    .I2(__54__),
    .I1(__64__),
    .I0(__135__),
    .O(__212__)
  );
  LUT6 #(
    .INIT(64'h3c00aaaa00000000)
  ) __585__ (
    .I5(__170__),
    .I4(__55__),
    .I3(__169__),
    .I2(__87__),
    .I1(__131__),
    .I0(__135__),
    .O(__213__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __586__ (
    .I1(__9__),
    .I0(__80__),
    .O(__214__)
  );
  LUT6 #(
    .INIT(64'h0000000000008000)
  ) __587__ (
    .I5(__109__),
    .I4(__56__),
    .I3(__214__),
    .I2(__181__),
    .I1(__158__),
    .I0(__111__),
    .O(__215__)
  );
  LUT5 #(
    .INIT(32'h80000000)
  ) __588__ (
    .I4(__120__),
    .I3(__16__),
    .I2(__139__),
    .I1(__136__),
    .I0(__8__),
    .O(__216__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __589__ (
    .I1(__23__),
    .I0(__190__),
    .O(__217__)
  );
  LUT6 #(
    .INIT(64'h0000000000000777)
  ) __590__ (
    .I5(__217__),
    .I4(__216__),
    .I3(__192__),
    .I2(g563),
    .I1(__195__),
    .I0(__11__),
    .O(__218__)
  );
  LUT5 #(
    .INIT(32'h00004000)
  ) __591__ (
    .I4(__40__),
    .I3(__120__),
    .I2(__16__),
    .I1(__139__),
    .I0(__136__),
    .O(__219__)
  );
  LUT4 #(
    .INIT(16'ha3ff)
  ) __592__ (
    .I3(__219__),
    .I2(__135__),
    .I1(__82__),
    .I0(__18__),
    .O(__220__)
  );
  LUT6 #(
    .INIT(64'h0000000080000000)
  ) __593__ (
    .I5(__109__),
    .I4(__95__),
    .I3(__9__),
    .I2(__80__),
    .I1(__186__),
    .I0(__35__),
    .O(__221__)
  );
  LUT6 #(
    .INIT(64'h0000000007770000)
  ) __594__ (
    .I5(__221__),
    .I4(__220__),
    .I3(__188__),
    .I2(__26__),
    .I1(__189__),
    .I0(__100__),
    .O(__222__)
  );
  LUT6 #(
    .INIT(64'h0007000000000000)
  ) __595__ (
    .I5(__222__),
    .I4(__218__),
    .I3(__185__),
    .I2(__215__),
    .I1(__135__),
    .I0(__0__),
    .O(__223__)
  );
  LUT3 #(
    .INIT(8'hef)
  ) __596__ (
    .I2(__223__),
    .I1(__213__),
    .I0(__212__),
    .O(__224__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __597__ (
    .I1(__39__),
    .I0(__104__),
    .O(__225__)
  );
  LUT6 #(
    .INIT(64'hff00000040404040)
  ) __598__ (
    .I5(__111__),
    .I4(__173__),
    .I3(__225__),
    .I2(__51__),
    .I1(__166__),
    .I0(__77__),
    .O(__226__)
  );
  LUT4 #(
    .INIT(16'h0008)
  ) __599__ (
    .I3(__109__),
    .I2(g41),
    .I1(__163__),
    .I0(__159__),
    .O(__227__)
  );
  LUT5 #(
    .INIT(32'hf0f07700)
  ) __600__ (
    .I4(__227__),
    .I3(__7__),
    .I2(__40__),
    .I1(__156__),
    .I0(__226__),
    .O(__228__)
  );
  LUT6 #(
    .INIT(64'h8000000000000000)
  ) __601__ (
    .I5(__79__),
    .I4(__20__),
    .I3(__75__),
    .I2(__106__),
    .I1(__138__),
    .I0(__83__),
    .O(__229__)
  );
  LUT3 #(
    .INIT(8'h60)
  ) __602__ (
    .I2(g639),
    .I1(__71__),
    .I0(__229__),
    .O(__230__)
  );
  LUT6 #(
    .INIT(64'h0000aaff00fcaafc)
  ) __603__ (
    .I5(__69__),
    .I4(__147__),
    .I3(__53__),
    .I2(__43__),
    .I1(__142__),
    .I0(__146__),
    .O(__231__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __604__ (
    .I2(__156__),
    .I1(__231__),
    .I0(__97__),
    .O(__232__)
  );
  LUT5 #(
    .INIT(32'hf1ffffff)
  ) __605__ (
    .I4(__108__),
    .I3(__33__),
    .I2(g22),
    .I1(g41),
    .I0(__205__),
    .O(__233__)
  );
  LUT5 #(
    .INIT(32'haaaaea2a)
  ) __606__ (
    .I4(g41),
    .I3(__40__),
    .I2(__163__),
    .I1(__190__),
    .I0(__123__),
    .O(__234__)
  );
  LUT5 #(
    .INIT(32'h80000000)
  ) __607__ (
    .I4(__104__),
    .I3(__54__),
    .I2(__64__),
    .I1(__93__),
    .I0(__103__),
    .O(__235__)
  );
  LUT6 #(
    .INIT(64'hfefe0000ff00ff00)
  ) __608__ (
    .I5(__23__),
    .I4(__174__),
    .I3(__95__),
    .I2(__39__),
    .I1(__202__),
    .I0(__235__),
    .O(__236__)
  );
  LUT5 #(
    .INIT(32'h80000000)
  ) __609__ (
    .I4(__77__),
    .I3(__87__),
    .I2(__129__),
    .I1(__49__),
    .I0(__131__),
    .O(__237__)
  );
  LUT4 #(
    .INIT(16'h0001)
  ) __610__ (
    .I3(__90__),
    .I2(__114__),
    .I1(__31__),
    .I0(__168__),
    .O(__238__)
  );
  LUT6 #(
    .INIT(64'hfefe0000ff00ff00)
  ) __611__ (
    .I5(__55__),
    .I4(__167__),
    .I3(__95__),
    .I2(__51__),
    .I1(__238__),
    .I0(__237__),
    .O(__239__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __612__ (
    .I5(__188__),
    .I4(__52__),
    .I3(__187__),
    .I2(__28__),
    .I1(__192__),
    .I0(g559),
    .O(__240__)
  );
  LUT5 #(
    .INIT(32'h07770000)
  ) __613__ (
    .I4(__240__),
    .I3(__95__),
    .I2(__0__),
    .I1(__195__),
    .I0(__76__),
    .O(__241__)
  );
  LUT6 #(
    .INIT(64'hfffff888ffffffff)
  ) __614__ (
    .I5(__241__),
    .I4(__185__),
    .I3(__170__),
    .I2(__239__),
    .I1(__177__),
    .I0(__236__),
    .O(__242__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __615__ (
    .I2(__54__),
    .I1(__64__),
    .I0(__103__),
    .O(__243__)
  );
  LUT6 #(
    .INIT(64'h00005ff5cccccccc)
  ) __616__ (
    .I5(__23__),
    .I4(__202__),
    .I3(__93__),
    .I2(__243__),
    .I1(__136__),
    .I0(__174__),
    .O(__244__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __617__ (
    .I1(g89),
    .I0(g102),
    .O(__245__)
  );
  LUT6 #(
    .INIT(64'h0f0f333300ff5555)
  ) __618__ (
    .I5(__87__),
    .I4(__131__),
    .I3(__40__),
    .I2(__109__),
    .I1(__135__),
    .I0(__136__),
    .O(__246__)
  );
  LUT6 #(
    .INIT(64'h0f0f333300ff5555)
  ) __619__ (
    .I5(__87__),
    .I4(__131__),
    .I3(__9__),
    .I2(__56__),
    .I1(__95__),
    .I0(__80__),
    .O(__247__)
  );
  LUT6 #(
    .INIT(64'ha5c300000000a5c3)
  ) __620__ (
    .I5(__51__),
    .I4(__77__),
    .I3(__49__),
    .I2(__31__),
    .I1(__247__),
    .I0(__246__),
    .O(__248__)
  );
  LUT6 #(
    .INIT(64'h7630ffff76300000)
  ) __621__ (
    .I5(__100__),
    .I4(__156__),
    .I3(__90__),
    .I2(__114__),
    .I1(__151__),
    .I0(__248__),
    .O(__249__)
  );
  LUT4 #(
    .INIT(16'h0660)
  ) __622__ (
    .I3(__51__),
    .I2(__77__),
    .I1(__31__),
    .I0(__168__),
    .O(__250__)
  );
  LUT6 #(
    .INIT(64'h000f020a030f030f)
  ) __623__ (
    .I5(__90__),
    .I4(__248__),
    .I3(__151__),
    .I2(__238__),
    .I1(__114__),
    .I0(__250__),
    .O(__251__)
  );
  LUT5 #(
    .INIT(32'heaebfaff)
  ) __624__ (
    .I4(__90__),
    .I3(__114__),
    .I2(__151__),
    .I1(__248__),
    .I0(__251__),
    .O(__252__)
  );
  LUT5 #(
    .INIT(32'h02ff0200)
  ) __625__ (
    .I4(__109__),
    .I3(__23__),
    .I2(__64__),
    .I1(__202__),
    .I0(__174__),
    .O(__253__)
  );
  LUT6 #(
    .INIT(64'hfaffffffffffffff)
  ) __626__ (
    .I5(g41),
    .I4(__108__),
    .I3(__33__),
    .I2(g22),
    .I1(__205__),
    .I0(__63__),
    .O(__254__)
  );
  LUT5 #(
    .INIT(32'haaacaaaa)
  ) __627__ (
    .I4(__156__),
    .I3(__7__),
    .I2(__74__),
    .I1(__13__),
    .I0(__28__),
    .O(__255__)
  );
  LUT5 #(
    .INIT(32'h80000000)
  ) __628__ (
    .I4(__62__),
    .I3(__92__),
    .I2(__44__),
    .I1(__128__),
    .I0(g567),
    .O(__256__)
  );
  LUT3 #(
    .INIT(8'h60)
  ) __629__ (
    .I2(__21__),
    .I1(__89__),
    .I0(__256__),
    .O(__257__)
  );
  LUT5 #(
    .INIT(32'h6ccc0000)
  ) __630__ (
    .I4(g639),
    .I3(__140__),
    .I2(__71__),
    .I1(__36__),
    .I0(__229__),
    .O(__258__)
  );
  LUT3 #(
    .INIT(8'h60)
  ) __631__ (
    .I2(g639),
    .I1(__75__),
    .I0(__83__),
    .O(__259__)
  );
  LUT5 #(
    .INIT(32'hcc4ccccc)
  ) __632__ (
    .I4(__109__),
    .I3(g41),
    .I2(__163__),
    .I1(__124__),
    .I0(__159__),
    .O(__260__)
  );
  LUT3 #(
    .INIT(8'h60)
  ) __633__ (
    .I2(__21__),
    .I1(__128__),
    .I0(g567),
    .O(__261__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __634__ (
    .I1(__75__),
    .I0(__83__),
    .O(__262__)
  );
  LUT6 #(
    .INIT(64'h7fff800000000000)
  ) __635__ (
    .I5(g639),
    .I4(__106__),
    .I3(__79__),
    .I2(__20__),
    .I1(__138__),
    .I0(__262__),
    .O(__263__)
  );
  LUT5 #(
    .INIT(32'haaacaaaa)
  ) __636__ (
    .I4(__156__),
    .I3(__7__),
    .I2(__74__),
    .I1(__81__),
    .I0(__30__),
    .O(__264__)
  );
  LUT5 #(
    .INIT(32'haaacaaaa)
  ) __637__ (
    .I4(__156__),
    .I3(__7__),
    .I2(__74__),
    .I1(__29__),
    .I0(__26__),
    .O(__265__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __638__ (
    .I1(g45),
    .I0(__88__),
    .O(__266__)
  );
  LUT6 #(
    .INIT(64'h7fff800000000000)
  ) __639__ (
    .I5(__21__),
    .I4(__92__),
    .I3(__62__),
    .I2(__44__),
    .I1(__128__),
    .I0(g567),
    .O(__267__)
  );
  LUT6 #(
    .INIT(64'hccccec4ccccccccc)
  ) __640__ (
    .I5(__109__),
    .I4(g41),
    .I3(__136__),
    .I2(__163__),
    .I1(__91__),
    .I0(__159__),
    .O(__268__)
  );
  LUT5 #(
    .INIT(32'hcccccc4c)
  ) __641__ (
    .I4(__109__),
    .I3(g41),
    .I2(__163__),
    .I1(__96__),
    .I0(__159__),
    .O(__269__)
  );
  LUT5 #(
    .INIT(32'haaacaaaa)
  ) __642__ (
    .I4(__156__),
    .I3(__7__),
    .I2(__74__),
    .I1(__35__),
    .I0(__24__),
    .O(__270__)
  );
  LUT6 #(
    .INIT(64'hccf0330faaaa5555)
  ) __643__ (
    .I5(__145__),
    .I4(__43__),
    .I3(__103__),
    .I2(__144__),
    .I1(__143__),
    .I0(__142__),
    .O(__271__)
  );
  LUT6 #(
    .INIT(64'h707b00ff00ff00bb)
  ) __644__ (
    .I5(__39__),
    .I4(__104__),
    .I3(__69__),
    .I2(__173__),
    .I1(__53__),
    .I0(__271__),
    .O(__272__)
  );
  LUT2 #(
    .INIT(4'he)
  ) __645__ (
    .I1(__272__),
    .I0(__231__),
    .O(__273__)
  );
  LUT6 #(
    .INIT(64'hfaffffffffffffff)
  ) __646__ (
    .I5(g41),
    .I4(__108__),
    .I3(__33__),
    .I2(g22),
    .I1(__205__),
    .I0(__94__),
    .O(__274__)
  );
  LUT4 #(
    .INIT(16'hff01)
  ) __647__ (
    .I3(__8__),
    .I2(g41),
    .I1(g22),
    .I0(__205__),
    .O(__275__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __648__ (
    .I2(__156__),
    .I1(__251__),
    .I0(__38__),
    .O(__276__)
  );
  LUT6 #(
    .INIT(64'h8000000000000000)
  ) __649__ (
    .I5(__70__),
    .I4(__140__),
    .I3(__71__),
    .I2(__36__),
    .I1(__37__),
    .I0(__229__),
    .O(__277__)
  );
  LUT5 #(
    .INIT(32'h7fff0000)
  ) __650__ (
    .I4(g639),
    .I3(__84__),
    .I2(__277__),
    .I1(__98__),
    .I0(__19__),
    .O(__278__)
  );
  LUT6 #(
    .INIT(64'h7fff800000000000)
  ) __651__ (
    .I5(__278__),
    .I4(__37__),
    .I3(__140__),
    .I2(__71__),
    .I1(__36__),
    .I0(__229__),
    .O(__279__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __652__ (
    .I1(__63__),
    .I0(__126__),
    .O(__280__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __653__ (
    .I1(__32__),
    .I0(__94__),
    .O(__281__)
  );
  LUT6 #(
    .INIT(64'h9669699669969669)
  ) __654__ (
    .I5(__107__),
    .I4(__130__),
    .I3(__25__),
    .I2(__72__),
    .I1(__281__),
    .I0(__280__),
    .O(__282__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __655__ (
    .I2(__156__),
    .I1(__272__),
    .I0(__119__),
    .O(__283__)
  );
  LUT5 #(
    .INIT(32'haaacaaaa)
  ) __656__ (
    .I4(__156__),
    .I3(__7__),
    .I2(__74__),
    .I1(__57__),
    .I0(__13__),
    .O(__284__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __657__ (
    .I2(__23__),
    .I1(__272__),
    .I0(__80__),
    .O(__285__)
  );
  LUT5 #(
    .INIT(32'h3c00aaaa)
  ) __658__ (
    .I4(__55__),
    .I3(__169__),
    .I2(__87__),
    .I1(__131__),
    .I0(__135__),
    .O(__286__)
  );
  LUT4 #(
    .INIT(16'hb0bb)
  ) __659__ (
    .I3(__101__),
    .I2(__34__),
    .I1(__82__),
    .I0(__18__),
    .O(__287__)
  );
  LUT6 #(
    .INIT(64'h7fff800000000000)
  ) __660__ (
    .I5(g639),
    .I4(__79__),
    .I3(__20__),
    .I2(__75__),
    .I1(__138__),
    .I0(__83__),
    .O(__288__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __661__ (
    .I1(g45),
    .I0(__115__),
    .O(__289__)
  );
  LUT6 #(
    .INIT(64'h2888ffff28880000)
  ) __662__ (
    .I5(__40__),
    .I4(__55__),
    .I3(__87__),
    .I2(__131__),
    .I1(__49__),
    .I0(__169__),
    .O(__290__)
  );
  LUT6 #(
    .INIT(64'h8000000000000000)
  ) __663__ (
    .I5(__89__),
    .I4(__62__),
    .I3(__92__),
    .I2(__44__),
    .I1(__128__),
    .I0(g567),
    .O(__291__)
  );
  LUT4 #(
    .INIT(16'h7800)
  ) __664__ (
    .I3(__21__),
    .I2(__15__),
    .I1(__121__),
    .I0(__291__),
    .O(__292__)
  );
  LUT6 #(
    .INIT(64'hccccec4ccccccccc)
  ) __665__ (
    .I5(__109__),
    .I4(g41),
    .I3(__135__),
    .I2(__163__),
    .I1(__11__),
    .I0(__159__),
    .O(__293__)
  );
  LUT6 #(
    .INIT(64'h02ff000002000000)
  ) __666__ (
    .I5(__109__),
    .I4(__170__),
    .I3(__55__),
    .I2(__131__),
    .I1(__238__),
    .I0(__167__),
    .O(__294__)
  );
  LUT6 #(
    .INIT(64'h02ff000002000000)
  ) __667__ (
    .I5(__109__),
    .I4(__177__),
    .I3(__23__),
    .I2(__64__),
    .I1(__202__),
    .I0(__174__),
    .O(__295__)
  );
  LUT4 #(
    .INIT(16'h4000)
  ) __668__ (
    .I3(__181__),
    .I2(__101__),
    .I1(__219__),
    .I0(__135__),
    .O(__296__)
  );
  LUT6 #(
    .INIT(64'h0000000000008000)
  ) __669__ (
    .I5(__40__),
    .I4(__135__),
    .I3(__181__),
    .I2(__183__),
    .I1(__136__),
    .I0(__42__),
    .O(__297__)
  );
  LUT6 #(
    .INIT(64'h0000000000000777)
  ) __670__ (
    .I5(__297__),
    .I4(__296__),
    .I3(__192__),
    .I2(g564),
    .I1(__96__),
    .I0(__194__),
    .O(__298__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __671__ (
    .I2(__181__),
    .I1(__135__),
    .I0(__219__),
    .O(__299__)
  );
  LUT6 #(
    .INIT(64'h0000707770777077)
  ) __672__ (
    .I5(__187__),
    .I4(__127__),
    .I3(__299__),
    .I2(__34__),
    .I1(__55__),
    .I0(__191__),
    .O(__300__)
  );
  LUT4 #(
    .INIT(16'h1d3f)
  ) __673__ (
    .I3(__189__),
    .I2(__29__),
    .I1(__188__),
    .I0(__38__),
    .O(__301__)
  );
  LUT5 #(
    .INIT(32'h70000000)
  ) __674__ (
    .I4(__301__),
    .I3(__300__),
    .I2(__298__),
    .I1(__195__),
    .I0(__50__),
    .O(__302__)
  );
  LUT6 #(
    .INIT(64'hfffffff8ffffffff)
  ) __675__ (
    .I5(__302__),
    .I4(__185__),
    .I3(__295__),
    .I2(__294__),
    .I1(__109__),
    .I0(__0__),
    .O(__303__)
  );
  LUT6 #(
    .INIT(64'h7630ffff76300000)
  ) __676__ (
    .I5(__80__),
    .I4(__55__),
    .I3(__90__),
    .I2(__114__),
    .I1(__151__),
    .I0(__248__),
    .O(__304__)
  );
  LUT6 #(
    .INIT(64'hfaffffffffffffff)
  ) __677__ (
    .I5(g41),
    .I4(__108__),
    .I3(__33__),
    .I2(g22),
    .I1(__205__),
    .I0(__282__),
    .O(__305__)
  );
  LUT6 #(
    .INIT(64'hfaffffffffffffff)
  ) __678__ (
    .I5(g41),
    .I4(__108__),
    .I3(__33__),
    .I2(g22),
    .I1(__205__),
    .I0(__25__),
    .O(__306__)
  );
  LUT5 #(
    .INIT(32'hcceccccc)
  ) __679__ (
    .I4(__109__),
    .I3(g41),
    .I2(__163__),
    .I1(__50__),
    .I0(__159__),
    .O(__307__)
  );
  LUT4 #(
    .INIT(16'h78ff)
  ) __680__ (
    .I3(g639),
    .I2(__138__),
    .I1(__75__),
    .I0(__83__),
    .O(__308__)
  );
  LUT5 #(
    .INIT(32'haaacaaaa)
  ) __681__ (
    .I4(__156__),
    .I3(__7__),
    .I2(__74__),
    .I1(__45__),
    .I0(__27__),
    .O(__309__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __682__ (
    .I5(__188__),
    .I4(__45__),
    .I3(__187__),
    .I2(__66__),
    .I1(__192__),
    .I0(g558),
    .O(__310__)
  );
  LUT6 #(
    .INIT(64'h0000000007770000)
  ) __683__ (
    .I5(__185__),
    .I4(__310__),
    .I3(__9__),
    .I2(__0__),
    .I1(__195__),
    .I0(__14__),
    .O(__311__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __684__ (
    .I2(__55__),
    .I1(__251__),
    .I0(__9__),
    .O(__312__)
  );
  LUT6 #(
    .INIT(64'hbb33f3f333333333)
  ) __685__ (
    .I5(__179__),
    .I4(__12__),
    .I3(__176__),
    .I2(__312__),
    .I1(__311__),
    .I0(__149__),
    .O(__313__)
  );
  LUT4 #(
    .INIT(16'hff40)
  ) __686__ (
    .I3(__82__),
    .I2(__69__),
    .I1(__53__),
    .I0(__271__),
    .O(__314__)
  );
  LUT5 #(
    .INIT(32'h80000000)
  ) __687__ (
    .I4(__140__),
    .I3(__71__),
    .I2(__36__),
    .I1(__37__),
    .I0(__229__),
    .O(__315__)
  );
  LUT3 #(
    .INIT(8'h60)
  ) __688__ (
    .I2(__278__),
    .I1(__70__),
    .I0(__315__),
    .O(__316__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __689__ (
    .I2(__87__),
    .I1(__49__),
    .I0(__131__),
    .O(__317__)
  );
  LUT6 #(
    .INIT(64'h00005ff5cccccccc)
  ) __690__ (
    .I5(__55__),
    .I4(__238__),
    .I3(__129__),
    .I2(__317__),
    .I1(__136__),
    .I0(__167__),
    .O(__318__)
  );
  LUT5 #(
    .INIT(32'haaacaaaa)
  ) __691__ (
    .I4(__156__),
    .I3(__7__),
    .I2(__74__),
    .I1(__24__),
    .I0(__57__),
    .O(__319__)
  );
  LUT6 #(
    .INIT(64'hf8f078f0ffffffff)
  ) __692__ (
    .I5(g639),
    .I4(__84__),
    .I3(__277__),
    .I2(__98__),
    .I1(__19__),
    .I0(__22__),
    .O(__320__)
  );
  LUT5 #(
    .INIT(32'hcceccccc)
  ) __693__ (
    .I4(__109__),
    .I3(g41),
    .I2(__163__),
    .I1(__14__),
    .I0(__159__),
    .O(__321__)
  );
  LUT6 #(
    .INIT(64'h7fff800000000000)
  ) __694__ (
    .I5(g639),
    .I4(__84__),
    .I3(__277__),
    .I2(__98__),
    .I1(__19__),
    .I0(__22__),
    .O(__322__)
  );
  LUT6 #(
    .INIT(64'hdffdffffdffd0000)
  ) __695__ (
    .I5(__56__),
    .I4(__55__),
    .I3(__77__),
    .I2(__166__),
    .I1(__238__),
    .I0(__167__),
    .O(__323__)
  );
  LUT5 #(
    .INIT(32'h02ff0200)
  ) __696__ (
    .I4(__109__),
    .I3(__55__),
    .I2(__131__),
    .I1(__238__),
    .I0(__167__),
    .O(__324__)
  );
  LUT5 #(
    .INIT(32'hcceccccc)
  ) __697__ (
    .I4(__109__),
    .I3(g41),
    .I2(__163__),
    .I1(__46__),
    .I0(__159__),
    .O(__325__)
  );
  LUT6 #(
    .INIT(64'h2888ffff28880000)
  ) __698__ (
    .I5(__40__),
    .I4(__23__),
    .I3(__54__),
    .I2(__64__),
    .I1(__103__),
    .I0(__175__),
    .O(__326__)
  );
  LUT5 #(
    .INIT(32'haaaaea2a)
  ) __699__ (
    .I4(g41),
    .I3(__135__),
    .I2(__163__),
    .I1(__190__),
    .I0(__23__),
    .O(__327__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __700__ (
    .I1(g639),
    .I0(__83__),
    .O(__328__)
  );
  LUT5 #(
    .INIT(32'haaacaaaa)
  ) __701__ (
    .I4(__156__),
    .I3(__7__),
    .I2(__74__),
    .I1(__28__),
    .I0(__66__),
    .O(__329__)
  );
  LUT2 #(
    .INIT(4'h7)
  ) __702__ (
    .I1(__21__),
    .I0(g567),
    .O(__330__)
  );
  LUT6 #(
    .INIT(64'hfaffffffffffffff)
  ) __703__ (
    .I5(g41),
    .I4(__108__),
    .I3(__33__),
    .I2(g22),
    .I1(__205__),
    .I0(__32__),
    .O(__331__)
  );
  LUT5 #(
    .INIT(32'hfef0f0f0)
  ) __704__ (
    .I4(__90__),
    .I3(__114__),
    .I2(__101__),
    .I1(__248__),
    .I0(__250__),
    .O(__332__)
  );
  LUT5 #(
    .INIT(32'h6ccc0000)
  ) __705__ (
    .I4(__21__),
    .I3(__121__),
    .I2(__291__),
    .I1(__65__),
    .I0(__15__),
    .O(__333__)
  );
  LUT5 #(
    .INIT(32'haaacaaaa)
  ) __706__ (
    .I4(__156__),
    .I3(__7__),
    .I2(__74__),
    .I1(__30__),
    .I0(__52__),
    .O(__334__)
  );
  LUT4 #(
    .INIT(16'haabe)
  ) __707__ (
    .I3(g22),
    .I2(__205__),
    .I1(__204__),
    .I0(__42__),
    .O(__335__)
  );
  LUT5 #(
    .INIT(32'h6ccc0000)
  ) __708__ (
    .I4(g639),
    .I3(__75__),
    .I2(__138__),
    .I1(__20__),
    .I0(__83__),
    .O(__336__)
  );
  LUT5 #(
    .INIT(32'haaacaaaa)
  ) __709__ (
    .I4(__156__),
    .I3(__7__),
    .I2(__74__),
    .I1(__26__),
    .I0(__78__),
    .O(__337__)
  );
  LUT6 #(
    .INIT(64'h0220ffff02200000)
  ) __710__ (
    .I5(__135__),
    .I4(__23__),
    .I3(__54__),
    .I2(__64__),
    .I1(__202__),
    .I0(__174__),
    .O(__338__)
  );
  LUT5 #(
    .INIT(32'haaacaaaa)
  ) __711__ (
    .I4(__156__),
    .I3(__7__),
    .I2(__74__),
    .I1(__52__),
    .I0(__45__),
    .O(__339__)
  );
  LUT6 #(
    .INIT(64'hfaffffffffffffff)
  ) __712__ (
    .I5(g41),
    .I4(__108__),
    .I3(__33__),
    .I2(g22),
    .I1(__205__),
    .I0(__130__),
    .O(__340__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __713__ (
    .I5(__188__),
    .I4(__30__),
    .I3(__187__),
    .I2(__13__),
    .I1(__192__),
    .I0(g560),
    .O(__341__)
  );
  LUT5 #(
    .INIT(32'h07770000)
  ) __714__ (
    .I4(__341__),
    .I3(__56__),
    .I2(__0__),
    .I1(__195__),
    .I0(__124__),
    .O(__342__)
  );
  LUT6 #(
    .INIT(64'hfffff888ffffffff)
  ) __715__ (
    .I5(__342__),
    .I4(__185__),
    .I3(__170__),
    .I2(__323__),
    .I1(__177__),
    .I0(__203__),
    .O(__343__)
  );
  LUT5 #(
    .INIT(32'haaacaaaa)
  ) __716__ (
    .I4(__156__),
    .I3(__7__),
    .I2(__74__),
    .I1(__78__),
    .I0(__81__),
    .O(__344__)
  );
  LUT5 #(
    .INIT(32'haaaaea2a)
  ) __717__ (
    .I4(g41),
    .I3(__109__),
    .I2(__163__),
    .I1(__190__),
    .I0(__55__),
    .O(__345__)
  );
  LUT6 #(
    .INIT(64'haaaaaaaaaaaaea2a)
  ) __718__ (
    .I5(__109__),
    .I4(g41),
    .I3(__135__),
    .I2(__163__),
    .I1(__159__),
    .I0(__111__),
    .O(__346__)
  );
  LUT5 #(
    .INIT(32'h5a5a0000)
  ) __719__ (
    .I4(g639),
    .I3(__84__),
    .I2(__277__),
    .I1(__98__),
    .I0(__19__),
    .O(__347__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __720__ (
    .I1(__156__),
    .I0(__7__),
    .O(__348__)
  );
  LUT6 #(
    .INIT(64'hf0f0ccaaf0f0f0f0)
  ) __721__ (
    .I5(__348__),
    .I4(__74__),
    .I3(__111__),
    .I2(__29__),
    .I1(__43__),
    .I0(__31__),
    .O(__349__)
  );
  LUT4 #(
    .INIT(16'h7800)
  ) __722__ (
    .I3(g639),
    .I2(__140__),
    .I1(__71__),
    .I0(__229__),
    .O(__350__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __723__ (
    .I1(__187__),
    .I0(__57__),
    .O(__351__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __724__ (
    .I1(__188__),
    .I0(__81__),
    .O(__352__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __725__ (
    .I5(__192__),
    .I4(g561),
    .I3(__191__),
    .I2(__102__),
    .I1(__119__),
    .I0(__189__),
    .O(__353__)
  );
  LUT4 #(
    .INIT(16'h0777)
  ) __726__ (
    .I3(__195__),
    .I2(__91__),
    .I1(__74__),
    .I0(__194__),
    .O(__354__)
  );
  LUT6 #(
    .INIT(64'h0007000000000000)
  ) __727__ (
    .I5(__354__),
    .I4(__353__),
    .I3(__352__),
    .I2(__351__),
    .I1(__136__),
    .I0(__0__),
    .O(__355__)
  );
  LUT6 #(
    .INIT(64'hfffff888ffffffff)
  ) __728__ (
    .I5(__355__),
    .I4(__185__),
    .I3(__170__),
    .I2(__318__),
    .I1(__177__),
    .I0(__244__),
    .O(__356__)
  );
  LUT4 #(
    .INIT(16'h8000)
  ) __729__ (
    .I3(__70__),
    .I2(__37__),
    .I1(__19__),
    .I0(__22__),
    .O(__357__)
  );
  LUT6 #(
    .INIT(64'hccccaaaaff00f0f0)
  ) __730__ (
    .I5(__70__),
    .I4(__37__),
    .I3(__9__),
    .I2(__80__),
    .I1(__56__),
    .I0(__95__),
    .O(__358__)
  );
  LUT6 #(
    .INIT(64'hccccaaaaff00f0f0)
  ) __731__ (
    .I5(__70__),
    .I4(__37__),
    .I3(__40__),
    .I2(__136__),
    .I1(__109__),
    .I0(__135__),
    .O(__359__)
  );
  LUT6 #(
    .INIT(64'hf0cc5555fffff0cc)
  ) __732__ (
    .I5(__84__),
    .I4(__98__),
    .I3(__19__),
    .I2(__359__),
    .I1(__358__),
    .I0(__357__),
    .O(__360__)
  );
  LUT5 #(
    .INIT(32'hcc4ccccc)
  ) __733__ (
    .I4(__109__),
    .I3(g41),
    .I2(__163__),
    .I1(__76__),
    .I0(__159__),
    .O(__361__)
  );
  LUT6 #(
    .INIT(64'hfaffffffffffffff)
  ) __734__ (
    .I5(g41),
    .I4(__108__),
    .I3(__33__),
    .I2(g22),
    .I1(__205__),
    .I0(__107__),
    .O(__362__)
  );
  LUT5 #(
    .INIT(32'haaacaaaa)
  ) __735__ (
    .I4(__156__),
    .I3(__7__),
    .I2(__74__),
    .I1(__27__),
    .I0(__127__),
    .O(__363__)
  );
  LUT4 #(
    .INIT(16'h3a00)
  ) __736__ (
    .I3(__177__),
    .I2(__23__),
    .I1(__272__),
    .I0(__80__),
    .O(__364__)
  );
  LUT4 #(
    .INIT(16'h89cf)
  ) __737__ (
    .I3(__90__),
    .I2(__114__),
    .I1(__151__),
    .I0(__248__),
    .O(__365__)
  );
  LUT5 #(
    .INIT(32'h00003a00)
  ) __738__ (
    .I4(__12__),
    .I3(__179__),
    .I2(__55__),
    .I1(__365__),
    .I0(__80__),
    .O(__366__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __739__ (
    .I5(__27__),
    .I4(__188__),
    .I3(__187__),
    .I2(__58__),
    .I1(g557),
    .I0(__192__),
    .O(__367__)
  );
  LUT3 #(
    .INIT(8'h70)
  ) __740__ (
    .I2(__367__),
    .I1(__195__),
    .I0(__46__),
    .O(__368__)
  );
  LUT6 #(
    .INIT(64'hfffffff8ffffffff)
  ) __741__ (
    .I5(__368__),
    .I4(__366__),
    .I3(__185__),
    .I2(__364__),
    .I1(__80__),
    .I0(__0__),
    .O(__369__)
  );
  LUT3 #(
    .INIT(8'h60)
  ) __742__ (
    .I2(__21__),
    .I1(__121__),
    .I0(__291__),
    .O(__370__)
  );
  LUT6 #(
    .INIT(64'he6aa66aaffffffff)
  ) __743__ (
    .I5(g639),
    .I4(__84__),
    .I3(__277__),
    .I2(__98__),
    .I1(__19__),
    .I0(__22__),
    .O(__371__)
  );
  assign g4100 = g36;
  assign g2584 = __245__;
  assign g4108 = g45;
  assign g6374 = __340__;
  assign g5692 = 1'b0;
  assign g6728 = 1'b0;
  assign g6372 = __209__;
  assign g4109 = g46;
  assign g4105 = g40;
  assign g4809 = __287__;
  assign g3222 = g705;
  assign g3600 = __67__;
  assign g5137 = __67__;
  assign g1293 = __133__;
  assign g1290 = __41__;
  assign g4104 = g22;
  assign g6370 = __274__;
  assign g4107 = g44;
  assign g4422 = g564;
  assign g4099 = g32;
  assign g6362 = __362__;
  assign g4098 = g23;
  assign g6360 = __210__;
  assign g6364 = __254__;
  assign g4106 = g42;
  assign g4103 = g39;
  assign g4321 = __59__;
  assign g5469 = __59__;
  assign g6368 = __331__;
  assign g6282 = __233__;
  assign g6284 = __305__;
  assign g4101 = g37;
  assign g6366 = __306__;
  assign g4112 = g47;
  assign g4307 = __112__;
  assign g5468 = __112__;
  assign g4121 = __330__;
  assign g4102 = g38;
  assign g4110 = g41;
endmodule
