module s13207 (
  CK,
  g1,
  g10,
  g1000,
  g1008,
  g1016,
  g1080,
  g11,
  g1194,
  g1196,
  g1198,
  g1202,
  g1203,
  g1206,
  g1234,
  g1553,
  g1554,
  g21,
  g22,
  g23,
  g24,
  g25,
  g26,
  g27,
  g28,
  g29,
  g30,
  g31,
  g32,
  g37,
  g41,
  g42,
  g43,
  g44,
  g45,
  g49,
  g633,
  g634,
  g635,
  g645,
  g647,
  g648,
  g690,
  g694,
  g698,
  g702,
  g722,
  g723,
  g751,
  g752,
  g753,
  g754,
  g755,
  g756,
  g757,
  g781,
  g786,
  g795,
  g9,
  g929,
  g941,
  g955,
  g962,
  g4657,
  g3191,
  g785,
  g6308,
  g4664,
  g1195,
  g7048,
  g7763,
  g6909,
  g6289,
  g9378,
  g6212,
  g7730,
  g1817,
  g206,
  g291,
  g372,
  g453,
  g534,
  g594,
  g7294,
  g7295,
  g7283,
  g4663,
  g8872,
  g6298,
  g6303,
  g6293,
  g6305,
  g3856,
  g8661,
  g6269,
  g8958,
  g8234,
  g9132,
  g3857,
  g6425,
  g8218,
  g6236,
  g7731,
  g4372,
  g4371,
  g1894,
  g4660,
  g5669,
  g7504,
  g1201,
  g6302,
  g3130,
  g7424,
  g6300,
  g9128,
  g9204,
  g6295,
  g6376,
  g9310,
  g7063,
  g8663,
  g5571,
  g6849,
  g6288,
  g9312,
  g1824,
  g9297,
  g6290,
  g4316,
  g1205,
  g9299,
  g5678,
  g7505,
  g3854,
  g1911,
  g5687,
  g7508,
  g3096,
  g7290,
  g6207,
  g7729,
  g1724,
  g1944,
  g7289,
  g5729,
  g1804,
  g7474,
  g2662,
  g6304,
  g1015,
  g6648,
  g8216,
  g1783,
  g7425,
  g2844,
  g3159,
  g7292,
  g7288,
  g6292,
  g7284,
  g5143,
  g7514,
  g1810,
  g9305,
  g6306,
  g1870,
  g6297,
  g1197,
  g3829,
  g3859,
  g3860,
  g6850,
  g7293,
  g6895,
  g7103,
  g9280,
  g4373,
  g6223,
  g7732,
  g1006,
  g6307,
  g9314,
  g4267,
  g1871,
  g7298,
  g1829,
  g6675,
  g8219,
  g7423,
  g6299,
  g6291,
  g7285,
  g7286,
  g4661,
  g5682,
  g7506,
  g9308,
  g7287,
  g1017,
  g3077,
  g6294,
  g5164,
  g7291,
  g6301,
  g1246,
  g2888,
  g1193,
  g1798,
  g6653,
  g8217,
  g4655,
  g5684,
  g7507,
  g6296,
  g4370
);
  input CK;
  wire CK;
  input g1;
  wire g1;
  input g10;
  wire g10;
  input g1000;
  wire g1000;
  input g1008;
  wire g1008;
  input g1016;
  wire g1016;
  input g1080;
  wire g1080;
  input g11;
  wire g11;
  input g1194;
  wire g1194;
  input g1196;
  wire g1196;
  input g1198;
  wire g1198;
  input g1202;
  wire g1202;
  input g1203;
  wire g1203;
  input g1206;
  wire g1206;
  input g1234;
  wire g1234;
  input g1553;
  wire g1553;
  input g1554;
  wire g1554;
  input g21;
  wire g21;
  input g22;
  wire g22;
  input g23;
  wire g23;
  input g24;
  wire g24;
  input g25;
  wire g25;
  input g26;
  wire g26;
  input g27;
  wire g27;
  input g28;
  wire g28;
  input g29;
  wire g29;
  input g30;
  wire g30;
  input g31;
  wire g31;
  input g32;
  wire g32;
  input g37;
  wire g37;
  input g41;
  wire g41;
  input g42;
  wire g42;
  input g43;
  wire g43;
  input g44;
  wire g44;
  input g45;
  wire g45;
  input g49;
  wire g49;
  input g633;
  wire g633;
  input g634;
  wire g634;
  input g635;
  wire g635;
  input g645;
  wire g645;
  input g647;
  wire g647;
  input g648;
  wire g648;
  input g690;
  wire g690;
  input g694;
  wire g694;
  input g698;
  wire g698;
  input g702;
  wire g702;
  input g722;
  wire g722;
  input g723;
  wire g723;
  input g751;
  wire g751;
  input g752;
  wire g752;
  input g753;
  wire g753;
  input g754;
  wire g754;
  input g755;
  wire g755;
  input g756;
  wire g756;
  input g757;
  wire g757;
  input g781;
  wire g781;
  input g786;
  wire g786;
  input g795;
  wire g795;
  input g9;
  wire g9;
  input g929;
  wire g929;
  input g941;
  wire g941;
  input g955;
  wire g955;
  input g962;
  wire g962;
  output g4657;
  wire g4657;
  output g3191;
  wire g3191;
  output g785;
  wire g785;
  output g6308;
  wire g6308;
  output g4664;
  wire g4664;
  output g1195;
  wire g1195;
  output g7048;
  wire g7048;
  output g7763;
  wire g7763;
  output g6909;
  wire g6909;
  output g6289;
  wire g6289;
  output g9378;
  wire g9378;
  output g6212;
  wire g6212;
  output g7730;
  wire g7730;
  output g1817;
  wire g1817;
  output g206;
  wire g206;
  output g291;
  wire g291;
  output g372;
  wire g372;
  output g453;
  wire g453;
  output g534;
  wire g534;
  output g594;
  wire g594;
  output g7294;
  wire g7294;
  output g7295;
  wire g7295;
  output g7283;
  wire g7283;
  output g4663;
  wire g4663;
  output g8872;
  wire g8872;
  output g6298;
  wire g6298;
  output g6303;
  wire g6303;
  output g6293;
  wire g6293;
  output g6305;
  wire g6305;
  output g3856;
  wire g3856;
  output g8661;
  wire g8661;
  output g6269;
  wire g6269;
  output g8958;
  wire g8958;
  output g8234;
  wire g8234;
  output g9132;
  wire g9132;
  output g3857;
  wire g3857;
  output g6425;
  wire g6425;
  output g8218;
  wire g8218;
  output g6236;
  wire g6236;
  output g7731;
  wire g7731;
  output g4372;
  wire g4372;
  output g4371;
  wire g4371;
  output g1894;
  wire g1894;
  output g4660;
  wire g4660;
  output g5669;
  wire g5669;
  output g7504;
  wire g7504;
  output g1201;
  wire g1201;
  output g6302;
  wire g6302;
  output g3130;
  wire g3130;
  output g7424;
  wire g7424;
  output g6300;
  wire g6300;
  output g9128;
  wire g9128;
  output g9204;
  wire g9204;
  output g6295;
  wire g6295;
  output g6376;
  wire g6376;
  output g9310;
  wire g9310;
  output g7063;
  wire g7063;
  output g8663;
  wire g8663;
  output g5571;
  wire g5571;
  output g6849;
  wire g6849;
  output g6288;
  wire g6288;
  output g9312;
  wire g9312;
  output g1824;
  wire g1824;
  output g9297;
  wire g9297;
  output g6290;
  wire g6290;
  output g4316;
  wire g4316;
  output g1205;
  wire g1205;
  output g9299;
  wire g9299;
  output g5678;
  wire g5678;
  output g7505;
  wire g7505;
  output g3854;
  wire g3854;
  output g1911;
  wire g1911;
  output g5687;
  wire g5687;
  output g7508;
  wire g7508;
  output g3096;
  wire g3096;
  output g7290;
  wire g7290;
  output g6207;
  wire g6207;
  output g7729;
  wire g7729;
  output g1724;
  wire g1724;
  output g1944;
  wire g1944;
  output g7289;
  wire g7289;
  output g5729;
  wire g5729;
  output g1804;
  wire g1804;
  output g7474;
  wire g7474;
  output g2662;
  wire g2662;
  output g6304;
  wire g6304;
  output g1015;
  wire g1015;
  output g6648;
  wire g6648;
  output g8216;
  wire g8216;
  output g1783;
  wire g1783;
  output g7425;
  wire g7425;
  output g2844;
  wire g2844;
  output g3159;
  wire g3159;
  output g7292;
  wire g7292;
  output g7288;
  wire g7288;
  output g6292;
  wire g6292;
  output g7284;
  wire g7284;
  output g5143;
  wire g5143;
  output g7514;
  wire g7514;
  output g1810;
  wire g1810;
  output g9305;
  wire g9305;
  output g6306;
  wire g6306;
  output g1870;
  wire g1870;
  output g6297;
  wire g6297;
  output g1197;
  wire g1197;
  output g3829;
  wire g3829;
  output g3859;
  wire g3859;
  output g3860;
  wire g3860;
  output g6850;
  wire g6850;
  output g7293;
  wire g7293;
  output g6895;
  wire g6895;
  output g7103;
  wire g7103;
  output g9280;
  wire g9280;
  output g4373;
  wire g4373;
  output g6223;
  wire g6223;
  output g7732;
  wire g7732;
  output g1006;
  wire g1006;
  output g6307;
  wire g6307;
  output g9314;
  wire g9314;
  output g4267;
  wire g4267;
  output g1871;
  wire g1871;
  output g7298;
  wire g7298;
  output g1829;
  wire g1829;
  output g6675;
  wire g6675;
  output g8219;
  wire g8219;
  output g7423;
  wire g7423;
  output g6299;
  wire g6299;
  output g6291;
  wire g6291;
  output g7285;
  wire g7285;
  output g7286;
  wire g7286;
  output g4661;
  wire g4661;
  output g5682;
  wire g5682;
  output g7506;
  wire g7506;
  output g9308;
  wire g9308;
  output g7287;
  wire g7287;
  output g1017;
  wire g1017;
  output g3077;
  wire g3077;
  output g6294;
  wire g6294;
  output g5164;
  wire g5164;
  output g7291;
  wire g7291;
  output g6301;
  wire g6301;
  output g1246;
  wire g1246;
  output g2888;
  wire g2888;
  output g1193;
  wire g1193;
  output g1798;
  wire g1798;
  output g6653;
  wire g6653;
  output g8217;
  wire g8217;
  output g4655;
  wire g4655;
  output g5684;
  wire g5684;
  output g7507;
  wire g7507;
  output g6296;
  wire g6296;
  output g4370;
  wire g4370;
  wire __0__;
  wire __1__;
  wire __2__;
  wire __3__;
  wire __4__;
  wire __5__;
  wire __6__;
  wire __7__;
  wire __8__;
  wire __9__;
  wire __10__;
  wire __11__;
  wire __12__;
  wire __13__;
  wire __14__;
  wire __15__;
  wire __16__;
  wire __17__;
  wire __18__;
  wire __19__;
  wire __20__;
  wire __21__;
  wire __22__;
  wire __23__;
  wire __24__;
  wire __25__;
  wire __26__;
  wire __27__;
  wire __28__;
  wire __29__;
  wire __30__;
  wire __31__;
  wire __32__;
  wire __33__;
  wire __34__;
  wire __35__;
  wire __36__;
  wire __37__;
  wire __38__;
  wire __39__;
  wire __40__;
  wire __41__;
  wire __42__;
  wire __43__;
  wire __44__;
  wire __45__;
  wire __46__;
  wire __47__;
  wire __48__;
  wire __49__;
  wire __50__;
  wire __51__;
  wire __52__;
  wire __53__;
  wire __54__;
  wire __55__;
  wire __56__;
  wire __57__;
  wire __58__;
  wire __59__;
  wire __60__;
  wire __61__;
  wire __62__;
  wire __63__;
  wire __64__;
  wire __65__;
  wire __66__;
  wire __67__;
  wire __68__;
  wire __69__;
  wire __70__;
  wire __71__;
  wire __72__;
  wire __73__;
  wire __74__;
  wire __75__;
  wire __76__;
  wire __77__;
  wire __78__;
  wire __79__;
  wire __80__;
  wire __81__;
  wire __82__;
  wire __83__;
  wire __84__;
  wire __85__;
  wire __86__;
  wire __87__;
  wire __88__;
  wire __89__;
  wire __90__;
  wire __91__;
  wire __92__;
  wire __93__;
  wire __94__;
  wire __95__;
  wire __96__;
  wire __97__;
  wire __98__;
  wire __99__;
  wire __100__;
  wire __101__;
  wire __102__;
  wire __103__;
  wire __104__;
  wire __105__;
  wire __106__;
  wire __107__;
  wire __108__;
  wire __109__;
  wire __110__;
  wire __111__;
  wire __112__;
  wire __113__;
  wire __114__;
  wire __115__;
  wire __116__;
  wire __117__;
  wire __118__;
  wire __119__;
  wire __120__;
  wire __121__;
  wire __122__;
  wire __123__;
  wire __124__;
  wire __125__;
  wire __126__;
  wire __127__;
  wire __128__;
  wire __129__;
  wire __130__;
  wire __131__;
  wire __132__;
  wire __133__;
  wire __134__;
  wire __135__;
  wire __136__;
  wire __137__;
  wire __138__;
  wire __139__;
  wire __140__;
  wire __141__;
  wire __142__;
  wire __143__;
  wire __144__;
  wire __145__;
  wire __146__;
  wire __147__;
  wire __148__;
  wire __149__;
  wire __150__;
  wire __151__;
  wire __152__;
  wire __153__;
  wire __154__;
  wire __155__;
  wire __156__;
  wire __157__;
  wire __158__;
  wire __159__;
  wire __160__;
  wire __161__;
  wire __162__;
  wire __163__;
  wire __164__;
  wire __165__;
  wire __166__;
  wire __167__;
  wire __168__;
  wire __169__;
  wire __170__;
  wire __171__;
  wire __172__;
  wire __173__;
  wire __174__;
  wire __175__;
  wire __176__;
  wire __177__;
  wire __178__;
  wire __179__;
  wire __180__;
  wire __181__;
  wire __182__;
  wire __183__;
  wire __184__;
  wire __185__;
  wire __186__;
  wire __187__;
  wire __188__;
  wire __189__;
  wire __190__;
  wire __191__;
  wire __192__;
  wire __193__;
  wire __194__;
  wire __195__;
  wire __196__;
  wire __197__;
  wire __198__;
  wire __199__;
  wire __200__;
  wire __201__;
  wire __202__;
  wire __203__;
  wire __204__;
  wire __205__;
  wire __206__;
  wire __207__;
  wire __208__;
  wire __209__;
  wire __210__;
  wire __211__;
  wire __212__;
  wire __213__;
  wire __214__;
  wire __215__;
  wire __216__;
  wire __217__;
  wire __218__;
  wire __219__;
  wire __220__;
  wire __221__;
  wire __222__;
  wire __223__;
  wire __224__;
  wire __225__;
  wire __226__;
  wire __227__;
  wire __228__;
  wire __229__;
  wire __230__;
  wire __231__;
  wire __232__;
  wire __233__;
  wire __234__;
  wire __235__;
  wire __236__;
  wire __237__;
  wire __238__;
  wire __239__;
  wire __240__;
  wire __241__;
  wire __242__;
  wire __243__;
  wire __244__;
  wire __245__;
  wire __246__;
  wire __247__;
  wire __248__;
  wire __249__;
  wire __250__;
  wire __251__;
  wire __252__;
  wire __253__;
  wire __254__;
  wire __255__;
  wire __256__;
  wire __257__;
  wire __258__;
  wire __259__;
  wire __260__;
  wire __261__;
  wire __262__;
  wire __263__;
  wire __264__;
  wire __265__;
  wire __266__;
  wire __267__;
  wire __268__;
  wire __269__;
  wire __270__;
  wire __271__;
  wire __272__;
  wire __273__;
  wire __274__;
  wire __275__;
  wire __276__;
  wire __277__;
  wire __278__;
  wire __279__;
  wire __280__;
  wire __281__;
  wire __282__;
  wire __283__;
  wire __284__;
  wire __285__;
  wire __286__;
  wire __287__;
  wire __288__;
  wire __289__;
  wire __290__;
  wire __291__;
  wire __292__;
  wire __293__;
  wire __294__;
  wire __295__;
  wire __296__;
  wire __297__;
  wire __298__;
  wire __299__;
  wire __300__;
  wire __301__;
  wire __302__;
  wire __303__;
  wire __304__;
  wire __305__;
  wire __306__;
  wire __307__;
  wire __308__;
  wire __309__;
  wire __310__;
  wire __311__;
  wire __312__;
  wire __313__;
  wire __314__;
  wire __315__;
  wire __316__;
  wire __317__;
  wire __318__;
  wire __319__;
  wire __320__;
  wire __321__;
  wire __322__;
  wire __323__;
  wire __324__;
  wire __325__;
  wire __326__;
  wire __327__;
  wire __328__;
  wire __329__;
  wire __330__;
  wire __331__;
  wire __332__;
  wire __333__;
  wire __334__;
  wire __335__;
  wire __336__;
  wire __337__;
  wire __338__;
  wire __339__;
  wire __340__;
  wire __341__;
  wire __342__;
  wire __343__;
  wire __344__;
  wire __345__;
  wire __346__;
  wire __347__;
  wire __348__;
  wire __349__;
  wire __350__;
  wire __351__;
  wire __352__;
  wire __353__;
  wire __354__;
  wire __355__;
  wire __356__;
  wire __357__;
  wire __358__;
  wire __359__;
  wire __360__;
  wire __361__;
  wire __362__;
  wire __363__;
  wire __364__;
  wire __365__;
  wire __366__;
  wire __367__;
  wire __368__;
  wire __369__;
  wire __370__;
  wire __371__;
  wire __372__;
  wire __373__;
  wire __374__;
  wire __375__;
  wire __376__;
  wire __377__;
  wire __378__;
  wire __379__;
  wire __380__;
  wire __381__;
  wire __382__;
  wire __383__;
  wire __384__;
  wire __385__;
  wire __386__;
  wire __387__;
  wire __388__;
  wire __389__;
  wire __390__;
  wire __391__;
  wire __392__;
  wire __393__;
  wire __394__;
  wire __395__;
  wire __396__;
  wire __397__;
  wire __398__;
  wire __399__;
  wire __400__;
  wire __401__;
  wire __402__;
  wire __403__;
  wire __404__;
  wire __405__;
  wire __406__;
  wire __407__;
  wire __408__;
  wire __409__;
  wire __410__;
  wire __411__;
  wire __412__;
  wire __413__;
  wire __414__;
  wire __415__;
  wire __416__;
  wire __417__;
  wire __418__;
  wire __419__;
  wire __420__;
  wire __421__;
  wire __422__;
  wire __423__;
  wire __424__;
  wire __425__;
  wire __426__;
  wire __427__;
  wire __428__;
  wire __429__;
  wire __430__;
  wire __431__;
  wire __432__;
  wire __433__;
  wire __434__;
  wire __435__;
  wire __436__;
  wire __437__;
  wire __438__;
  wire __439__;
  wire __440__;
  wire __441__;
  wire __442__;
  wire __443__;
  wire __444__;
  wire __445__;
  wire __446__;
  wire __447__;
  wire __448__;
  wire __449__;
  wire __450__;
  wire __451__;
  wire __452__;
  wire __453__;
  wire __454__;
  wire __455__;
  wire __456__;
  wire __457__;
  wire __458__;
  wire __459__;
  wire __460__;
  wire __461__;
  wire __462__;
  wire __463__;
  wire __464__;
  wire __465__;
  wire __466__;
  wire __467__;
  wire __468__;
  wire __469__;
  wire __470__;
  wire __471__;
  wire __472__;
  wire __473__;
  wire __474__;
  wire __475__;
  wire __476__;
  wire __477__;
  wire __478__;
  wire __479__;
  wire __480__;
  wire __481__;
  wire __482__;
  wire __483__;
  wire __484__;
  wire __485__;
  wire __486__;
  wire __487__;
  wire __488__;
  wire __489__;
  wire __490__;
  wire __491__;
  wire __492__;
  wire __493__;
  wire __494__;
  wire __495__;
  wire __496__;
  wire __498__;
  wire __500__;
  wire __501__;
  wire __502__;
  wire __503__;
  wire __504__;
  wire __505__;
  wire __506__;
  wire __507__;
  wire __508__;
  wire __509__;
  wire __510__;
  wire __511__;
  wire __512__;
  wire __513__;
  wire __514__;
  wire __515__;
  wire __516__;
  wire __517__;
  wire __518__;
  wire __519__;
  wire __520__;
  wire __521__;
  wire __522__;
  wire __523__;
  wire __524__;
  wire __525__;
  wire __526__;
  wire __527__;
  wire __528__;
  wire __529__;
  wire __530__;
  wire __531__;
  wire __532__;
  wire __533__;
  wire __534__;
  wire __535__;
  wire __536__;
  wire __537__;
  wire __538__;
  wire __539__;
  wire __540__;
  wire __541__;
  wire __542__;
  wire __543__;
  wire __544__;
  wire __545__;
  wire __546__;
  wire __547__;
  wire __548__;
  wire __549__;
  wire __550__;
  wire __551__;
  wire __552__;
  wire __553__;
  wire __554__;
  wire __555__;
  wire __556__;
  wire __557__;
  wire __558__;
  wire __559__;
  wire __560__;
  wire __561__;
  wire __562__;
  wire __563__;
  wire __564__;
  wire __565__;
  wire __566__;
  wire __567__;
  wire __568__;
  wire __569__;
  wire __570__;
  wire __571__;
  wire __572__;
  wire __573__;
  wire __574__;
  wire __575__;
  wire __576__;
  wire __577__;
  wire __578__;
  wire __579__;
  wire __580__;
  wire __581__;
  wire __582__;
  wire __583__;
  wire __584__;
  wire __585__;
  wire __586__;
  wire __587__;
  wire __588__;
  wire __589__;
  wire __590__;
  wire __591__;
  wire __592__;
  wire __593__;
  wire __594__;
  wire __595__;
  wire __596__;
  wire __597__;
  wire __598__;
  wire __599__;
  wire __600__;
  wire __601__;
  wire __602__;
  wire __603__;
  wire __604__;
  wire __605__;
  wire __606__;
  wire __607__;
  wire __608__;
  wire __609__;
  wire __610__;
  wire __611__;
  wire __612__;
  wire __613__;
  wire __614__;
  wire __615__;
  wire __616__;
  wire __617__;
  wire __618__;
  wire __619__;
  wire __620__;
  wire __621__;
  wire __622__;
  wire __623__;
  wire __624__;
  wire __625__;
  wire __626__;
  wire __627__;
  wire __628__;
  wire __629__;
  wire __630__;
  wire __631__;
  wire __632__;
  wire __633__;
  wire __634__;
  wire __635__;
  wire __636__;
  wire __637__;
  wire __638__;
  wire __639__;
  wire __640__;
  wire __641__;
  wire __642__;
  wire __643__;
  wire __644__;
  wire __645__;
  wire __646__;
  wire __647__;
  wire __648__;
  wire __649__;
  wire __650__;
  wire __651__;
  wire __652__;
  wire __653__;
  wire __654__;
  wire __655__;
  wire __656__;
  wire __657__;
  wire __658__;
  wire __659__;
  wire __660__;
  wire __661__;
  wire __662__;
  wire __663__;
  wire __664__;
  wire __665__;
  wire __666__;
  wire __667__;
  wire __668__;
  wire __669__;
  wire __670__;
  wire __671__;
  wire __672__;
  wire __673__;
  wire __674__;
  wire __675__;
  wire __676__;
  wire __677__;
  wire __678__;
  wire __679__;
  wire __680__;
  wire __681__;
  wire __682__;
  wire __683__;
  wire __684__;
  wire __685__;
  wire __686__;
  wire __687__;
  wire __688__;
  wire __689__;
  wire __690__;
  wire __691__;
  wire __692__;
  wire __693__;
  wire __694__;
  wire __695__;
  wire __696__;
  wire __697__;
  wire __698__;
  wire __699__;
  wire __700__;
  wire __701__;
  wire __702__;
  wire __703__;
  wire __704__;
  wire __705__;
  wire __706__;
  wire __707__;
  wire __708__;
  wire __709__;
  wire __710__;
  wire __711__;
  wire __712__;
  wire __713__;
  wire __714__;
  wire __715__;
  wire __716__;
  wire __717__;
  wire __718__;
  wire __719__;
  wire __720__;
  wire __721__;
  wire __722__;
  wire __723__;
  wire __724__;
  wire __725__;
  wire __726__;
  wire __727__;
  wire __728__;
  wire __729__;
  wire __730__;
  wire __731__;
  wire __732__;
  wire __733__;
  wire __734__;
  wire __735__;
  wire __736__;
  wire __737__;
  wire __738__;
  wire __739__;
  wire __740__;
  wire __741__;
  wire __742__;
  wire __743__;
  wire __744__;
  wire __745__;
  wire __746__;
  wire __747__;
  wire __748__;
  wire __749__;
  wire __750__;
  wire __751__;
  wire __752__;
  wire __753__;
  wire __754__;
  wire __755__;
  wire __756__;
  wire __757__;
  wire __758__;
  wire __759__;
  wire __760__;
  wire __761__;
  wire __762__;
  wire __763__;
  wire __764__;
  wire __765__;
  wire __766__;
  wire __767__;
  wire __768__;
  wire __769__;
  wire __770__;
  wire __771__;
  wire __772__;
  wire __773__;
  wire __774__;
  wire __775__;
  wire __776__;
  wire __777__;
  wire __778__;
  wire __779__;
  wire __780__;
  wire __781__;
  wire __782__;
  wire __783__;
  wire __784__;
  wire __785__;
  wire __786__;
  wire __787__;
  wire __788__;
  wire __789__;
  wire __790__;
  wire __791__;
  wire __792__;
  wire __793__;
  wire __794__;
  wire __795__;
  wire __796__;
  wire __797__;
  wire __798__;
  wire __799__;
  wire __800__;
  wire __801__;
  wire __802__;
  wire __803__;
  wire __804__;
  wire __805__;
  wire __806__;
  wire __807__;
  wire __808__;
  wire __809__;
  wire __810__;
  wire __811__;
  wire __812__;
  wire __813__;
  wire __814__;
  wire __815__;
  wire __816__;
  wire __817__;
  wire __818__;
  wire __819__;
  wire __820__;
  wire __821__;
  wire __822__;
  wire __823__;
  wire __824__;
  wire __825__;
  wire __826__;
  wire __827__;
  wire __828__;
  wire __829__;
  wire __830__;
  wire __831__;
  wire __832__;
  wire __833__;
  wire __834__;
  wire __835__;
  wire __836__;
  wire __837__;
  wire __838__;
  wire __839__;
  wire __840__;
  wire __841__;
  wire __842__;
  wire __843__;
  wire __844__;
  wire __845__;
  wire __846__;
  wire __847__;
  wire __848__;
  wire __849__;
  wire __850__;
  wire __851__;
  wire __852__;
  wire __853__;
  wire __854__;
  wire __855__;
  wire __856__;
  wire __857__;
  wire __858__;
  wire __859__;
  wire __860__;
  wire __861__;
  wire __862__;
  wire __863__;
  wire __864__;
  wire __865__;
  wire __866__;
  wire __867__;
  wire __868__;
  wire __869__;
  wire __870__;
  wire __871__;
  wire __872__;
  wire __873__;
  wire __874__;
  wire __875__;
  wire __876__;
  wire __877__;
  wire __878__;
  wire __879__;
  wire __880__;
  wire __881__;
  wire __882__;
  wire __883__;
  wire __884__;
  wire __885__;
  wire __886__;
  wire __887__;
  wire __888__;
  wire __889__;
  wire __890__;
  wire __891__;
  wire __892__;
  wire __893__;
  wire __894__;
  wire __895__;
  wire __896__;
  wire __897__;
  wire __898__;
  wire __899__;
  wire __900__;
  wire __901__;
  wire __902__;
  wire __903__;
  wire __904__;
  wire __905__;
  wire __906__;
  wire __907__;
  wire __908__;
  wire __909__;
  wire __910__;
  wire __911__;
  wire __912__;
  wire __913__;
  wire __914__;
  wire __915__;
  wire __916__;
  wire __917__;
  wire __918__;
  wire __919__;
  wire __920__;
  wire __921__;
  wire __922__;
  wire __923__;
  wire __924__;
  wire __925__;
  wire __926__;
  wire __927__;
  wire __928__;
  wire __929__;
  wire __930__;
  wire __931__;
  wire __932__;
  wire __933__;
  wire __934__;
  wire __935__;
  wire __936__;
  wire __937__;
  wire __938__;
  wire __939__;
  wire __940__;
  wire __941__;
  wire __942__;
  wire __943__;
  wire __944__;
  wire __945__;
  wire __946__;
  wire __947__;
  wire __948__;
  wire __949__;
  wire __950__;
  wire __951__;
  wire __952__;
  wire __953__;
  wire __954__;
  wire __955__;
  wire __956__;
  wire __957__;
  wire __958__;
  wire __959__;
  wire __960__;
  wire __961__;
  wire __962__;
  wire __963__;
  wire __964__;
  wire __965__;
  wire __966__;
  wire __967__;
  wire __968__;
  wire __969__;
  wire __970__;
  wire __971__;
  wire __972__;
  wire __973__;
  wire __974__;
  wire __975__;
  wire __976__;
  wire __977__;
  wire __978__;
  wire __979__;
  wire __980__;
  wire __981__;
  wire __982__;
  wire __983__;
  wire __984__;
  wire __985__;
  wire __986__;
  wire __987__;
  wire __988__;
  wire __989__;
  wire __990__;
  wire __991__;
  wire __992__;
  wire __993__;
  wire __994__;
  wire __995__;
  wire __996__;
  wire __997__;
  wire __998__;
  wire __999__;
  wire __1000__;
  wire __1001__;
  wire __1002__;
  wire __1003__;
  wire __1004__;
  wire __1005__;
  wire __1006__;
  wire __1007__;
  wire __1008__;
  wire __1009__;
  wire __1010__;
  wire __1011__;
  wire __1012__;
  wire __1013__;
  wire __1014__;
  wire __1015__;
  wire __1016__;
  wire __1017__;
  wire __1018__;
  wire __1019__;
  wire __1020__;
  wire __1021__;
  wire __1022__;
  wire __1023__;
  wire __1024__;
  wire __1025__;
  wire __1026__;
  wire __1027__;
  wire __1028__;
  wire __1029__;
  wire __1030__;
  wire __1031__;
  wire __1032__;
  wire __1033__;
  wire __1034__;
  wire __1035__;
  wire __1036__;
  wire __1037__;
  wire __1038__;
  wire __1039__;
  wire __1040__;
  wire __1041__;
  wire __1042__;
  wire __1043__;
  wire __1044__;
  wire __1045__;
  wire __1046__;
  wire __1047__;
  wire __1048__;
  wire __1049__;
  wire __1050__;
  wire __1051__;
  wire __1052__;
  wire __1053__;
  wire __1054__;
  wire __1055__;
  wire __1056__;
  wire __1057__;
  wire __1058__;
  wire __1059__;
  wire __1060__;
  wire __1061__;
  wire __1062__;
  wire __1063__;
  wire __1064__;
  wire __1065__;
  wire __1066__;
  wire __1067__;
  wire __1068__;
  wire __1069__;
  wire __1070__;
  wire __1071__;
  wire __1072__;
  wire __1073__;
  wire __1074__;
  wire __1075__;
  wire __1076__;
  wire __1077__;
  wire __1078__;
  wire __1079__;
  wire __1080__;
  wire __1081__;
  wire __1082__;
  wire __1083__;
  wire __1084__;
  wire __1085__;
  wire __1086__;
  INV __1087__ (
    .I(__503__),
    .O(__0__)
  );
  INV __1088__ (
    .I(__430__),
    .O(__1__)
  );
  INV __1089__ (
    .I(__330__),
    .O(__2__)
  );
  INV __1090__ (
    .I(__416__),
    .O(__3__)
  );
  INV __1091__ (
    .I(__62__),
    .O(__4__)
  );
  INV __1092__ (
    .I(__87__),
    .O(__5__)
  );
  INV __1093__ (
    .I(__212__),
    .O(__6__)
  );
  INV __1094__ (
    .I(__70__),
    .O(__7__)
  );
  INV __1095__ (
    .I(g43),
    .O(__8__)
  );
  INV __1096__ (
    .I(__180__),
    .O(__9__)
  );
  INV __1097__ (
    .I(g929),
    .O(__10__)
  );
  INV __1098__ (
    .I(g955),
    .O(__11__)
  );
  INV __1099__ (
    .I(g795),
    .O(__12__)
  );
  INV __1100__ (
    .I(__261__),
    .O(__13__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1101__ (
    .D(__579__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__14__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1102__ (
    .D(__1021__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__15__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1103__ (
    .D(__921__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__16__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1104__ (
    .D(__875__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__17__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1105__ (
    .D(__808__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__18__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1106__ (
    .D(__1003__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__19__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1107__ (
    .D(__132__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__20__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1108__ (
    .D(__975__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__21__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1109__ (
    .D(g26),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__22__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1110__ (
    .D(__135__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__23__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1111__ (
    .D(__779__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__24__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1112__ (
    .D(__996__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__25__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1113__ (
    .D(__682__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__26__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1114__ (
    .D(__195__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__27__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1115__ (
    .D(__5__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__28__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1116__ (
    .D(__853__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__29__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1117__ (
    .D(g27),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__30__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1118__ (
    .D(g23),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__31__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1119__ (
    .D(__243__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__32__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1120__ (
    .D(__508__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__33__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1121__ (
    .D(__780__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__34__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1122__ (
    .D(__724__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__35__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1123__ (
    .D(__584__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__36__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1124__ (
    .D(__258__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__37__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1125__ (
    .D(__577__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__38__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1126__ (
    .D(__922__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__39__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1127__ (
    .D(__998__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__40__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1128__ (
    .D(__993__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__41__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1129__ (
    .D(__1073__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__42__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1130__ (
    .D(__986__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__43__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1131__ (
    .D(__400__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__44__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1132__ (
    .D(__797__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__45__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1133__ (
    .D(__781__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__46__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1134__ (
    .D(__896__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__47__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1135__ (
    .D(__880__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__48__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1136__ (
    .D(__772__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__49__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1137__ (
    .D(__952__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__50__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1138__ (
    .D(__545__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__51__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1139__ (
    .D(__447__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__52__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1140__ (
    .D(__701__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__53__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1141__ (
    .D(__1036__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__54__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1142__ (
    .D(__846__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__55__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1143__ (
    .D(__773__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__56__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1144__ (
    .D(__1046__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__57__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1145__ (
    .D(__891__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__58__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1146__ (
    .D(__1010__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__59__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1147__ (
    .D(__946__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__60__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1148__ (
    .D(__860__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__61__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1149__ (
    .D(__699__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__62__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1150__ (
    .D(g1),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__63__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1151__ (
    .D(__1000__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__64__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1152__ (
    .D(__472__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__65__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1153__ (
    .D(__120__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__66__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1154__ (
    .D(__983__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__67__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1155__ (
    .D(__255__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__68__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1156__ (
    .D(__743__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__69__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1157__ (
    .D(__7__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__70__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1158__ (
    .D(__279__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__71__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1159__ (
    .D(__1020__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__72__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1160__ (
    .D(__618__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__73__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1161__ (
    .D(__489__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__74__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1162__ (
    .D(__897__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__75__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1163__ (
    .D(__802__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__76__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1164__ (
    .D(__706__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__77__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1165__ (
    .D(__798__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__78__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1166__ (
    .D(__626__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__79__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1167__ (
    .D(__473__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__80__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1168__ (
    .D(__342__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__81__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1169__ (
    .D(g1202),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__82__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1170__ (
    .D(__1011__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__83__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1171__ (
    .D(__929__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__84__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1172__ (
    .D(__439__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__85__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1173__ (
    .D(__1080__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__86__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1174__ (
    .D(__980__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__87__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1175__ (
    .D(__770__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__88__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1176__ (
    .D(__813__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__89__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1177__ (
    .D(__1053__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__90__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1178__ (
    .D(__938__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__91__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1179__ (
    .D(__979__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__92__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1180__ (
    .D(__928__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__93__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1181__ (
    .D(__959__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__94__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1182__ (
    .D(__222__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__95__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1183__ (
    .D(__1018__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__96__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1184__ (
    .D(__1032__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__97__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1185__ (
    .D(__992__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__98__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1186__ (
    .D(__106__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__99__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1187__ (
    .D(__1004__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__100__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1188__ (
    .D(g29),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__101__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1189__ (
    .D(__1014__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__102__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1190__ (
    .D(__769__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__103__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1191__ (
    .D(__1075__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__104__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1192__ (
    .D(__61__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__105__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1193__ (
    .D(__228__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__106__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1194__ (
    .D(__824__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__107__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1195__ (
    .D(__1071__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__108__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1196__ (
    .D(__145__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__109__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1197__ (
    .D(__818__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__110__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1198__ (
    .D(__567__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__111__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1199__ (
    .D(__568__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__112__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1200__ (
    .D(__95__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__113__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1201__ (
    .D(__994__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__114__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1202__ (
    .D(__898__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__115__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1203__ (
    .D(__886__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__116__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1204__ (
    .D(__1044__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__117__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1205__ (
    .D(__1033__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__118__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1206__ (
    .D(__845__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__119__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1207__ (
    .D(__474__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__120__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1208__ (
    .D(__914__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__121__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1209__ (
    .D(__835__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__122__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1210__ (
    .D(__696__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__123__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1211__ (
    .D(__1043__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__124__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1212__ (
    .D(__832__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__125__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1213__ (
    .D(__757__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__126__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1214__ (
    .D(__732__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__127__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1215__ (
    .D(__988__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__128__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1216__ (
    .D(__812__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__129__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1217__ (
    .D(__570__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__130__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1218__ (
    .D(__746__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__131__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1219__ (
    .D(__308__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__132__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1220__ (
    .D(__848__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__133__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1221__ (
    .D(__587__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__134__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1222__ (
    .D(__286__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__135__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1223__ (
    .D(__810__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__136__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1224__ (
    .D(__32__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__137__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1225__ (
    .D(__956__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__138__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1226__ (
    .D(__736__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__139__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1227__ (
    .D(__868__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__140__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1228__ (
    .D(__733__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__141__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1229__ (
    .D(__269__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__142__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1230__ (
    .D(__720__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__143__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1231__ (
    .D(__985__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__144__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1232__ (
    .D(__506__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__145__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1233__ (
    .D(__2__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__146__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1234__ (
    .D(g1194),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__147__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1235__ (
    .D(__1060__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__148__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1236__ (
    .D(__185__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__149__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1237__ (
    .D(__566__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__150__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1238__ (
    .D(__200__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__151__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1239__ (
    .D(__987__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__152__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1240__ (
    .D(__1061__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__153__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1241__ (
    .D(__837__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__154__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1242__ (
    .D(__1079__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__155__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1243__ (
    .D(__79__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__156__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1244__ (
    .D(__795__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__157__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1245__ (
    .D(__1002__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__158__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1246__ (
    .D(__1057__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__159__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1247__ (
    .D(__320__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__160__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1248__ (
    .D(__1045__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__161__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1249__ (
    .D(__1084__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__162__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1250__ (
    .D(__221__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__163__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1251__ (
    .D(__173__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__164__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1252__ (
    .D(__965__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__165__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1253__ (
    .D(__588__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__166__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1254__ (
    .D(__1052__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__167__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1255__ (
    .D(__931__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__168__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1256__ (
    .D(__1026__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__169__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1257__ (
    .D(__1009__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__170__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1258__ (
    .D(__903__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__171__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1259__ (
    .D(__739__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__172__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1260__ (
    .D(__216__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__173__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1261__ (
    .D(__1051__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__174__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1262__ (
    .D(__229__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__175__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1263__ (
    .D(__792__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__176__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1264__ (
    .D(__9__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__177__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1265__ (
    .D(__972__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__178__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1266__ (
    .D(__1086__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__179__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1267__ (
    .D(__912__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__180__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1268__ (
    .D(__704__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__181__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1269__ (
    .D(__1040__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__182__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1270__ (
    .D(__1025__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__183__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1271__ (
    .D(__1019__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__184__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1272__ (
    .D(__791__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__185__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1273__ (
    .D(__796__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__186__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1274__ (
    .D(__698__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__187__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1275__ (
    .D(__501__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__188__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1276__ (
    .D(__709__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__189__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1277__ (
    .D(__885__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__190__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1278__ (
    .D(__220__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__191__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1279__ (
    .D(__457__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__192__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1280__ (
    .D(__788__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__193__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1281__ (
    .D(__1034__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__194__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1282__ (
    .D(__348__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__195__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1283__ (
    .D(__1068__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__196__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1284__ (
    .D(__73__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__197__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1285__ (
    .D(__55__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__198__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1286__ (
    .D(__1005__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__199__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1287__ (
    .D(__213__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__200__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1288__ (
    .D(__156__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__201__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1289__ (
    .D(__963__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__202__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1290__ (
    .D(__319__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__203__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1291__ (
    .D(__735__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__204__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1292__ (
    .D(__713__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__205__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1293__ (
    .D(__1059__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__206__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1294__ (
    .D(g941),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__207__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1295__ (
    .D(__801__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__208__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1296__ (
    .D(__1055__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__209__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1297__ (
    .D(__977__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__210__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1298__ (
    .D(__3__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__211__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1299__ (
    .D(__867__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__212__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1300__ (
    .D(__23__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__213__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1301__ (
    .D(__951__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__214__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1302__ (
    .D(1'b0),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__215__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1303__ (
    .D(__607__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__216__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1304__ (
    .D(__1063__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__217__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1305__ (
    .D(__582__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__218__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1306__ (
    .D(__953__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__219__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1307__ (
    .D(__995__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__220__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1308__ (
    .D(__251__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__221__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1309__ (
    .D(__355__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__222__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1310__ (
    .D(__1008__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__223__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1311__ (
    .D(g22),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__224__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1312__ (
    .D(__906__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__225__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1313__ (
    .D(__847__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__226__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1314__ (
    .D(__785__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__227__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1315__ (
    .D(__211__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__228__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1316__ (
    .D(g24),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__229__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1317__ (
    .D(__539__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__230__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1318__ (
    .D(__923__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__231__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1319__ (
    .D(__807__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__232__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1320__ (
    .D(__312__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__233__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1321__ (
    .D(__175__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__234__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1322__ (
    .D(__65__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__235__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1323__ (
    .D(__680__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__236__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1324__ (
    .D(__940__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__237__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1325__ (
    .D(__432__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__238__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1326__ (
    .D(g1234),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__239__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1327__ (
    .D(__1028__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__240__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1328__ (
    .D(__1022__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__241__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1329__ (
    .D(__919__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__242__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1330__ (
    .D(__139__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__243__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1331__ (
    .D(__982__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__244__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1332__ (
    .D(__870__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__245__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1333__ (
    .D(__863__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__246__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1334__ (
    .D(__415__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__247__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1335__ (
    .D(__686__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__248__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1336__ (
    .D(__481__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__249__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1337__ (
    .D(__794__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__250__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1338__ (
    .D(__864__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__251__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1339__ (
    .D(__800__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__252__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1340__ (
    .D(__205__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__253__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1341__ (
    .D(__833__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__254__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1342__ (
    .D(__830__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__255__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1343__ (
    .D(__300__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__256__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1344__ (
    .D(__1015__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__257__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1345__ (
    .D(__389__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__258__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1346__ (
    .D(__505__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__259__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1347__ (
    .D(__877__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__260__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1348__ (
    .D(__363__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__261__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1349__ (
    .D(__1039__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__262__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1350__ (
    .D(__718__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__263__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1351__ (
    .D(__970__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__264__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1352__ (
    .D(__465__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__265__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1353__ (
    .D(g1203),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__266__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1354__ (
    .D(__538__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__267__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1355__ (
    .D(__740__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__268__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1356__ (
    .D(__13__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__269__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1357__ (
    .D(__87__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__270__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1358__ (
    .D(__937__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__271__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1359__ (
    .D(__285__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__272__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1360__ (
    .D(__823__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__273__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1361__ (
    .D(__188__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__274__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1362__ (
    .D(__727__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__275__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1363__ (
    .D(__1056__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__276__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1364__ (
    .D(__190__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__277__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1365__ (
    .D(__742__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__278__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1366__ (
    .D(__1062__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__279__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1367__ (
    .D(__945__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__280__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1368__ (
    .D(__1030__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__281__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1369__ (
    .D(__990__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__282__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1370__ (
    .D(__790__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__283__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1371__ (
    .D(__1058__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__284__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1372__ (
    .D(__534__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__285__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1373__ (
    .D(__344__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__286__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1374__ (
    .D(__729__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__287__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1375__ (
    .D(__45__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__288__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1376__ (
    .D(__137__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__289__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1377__ (
    .D(__883__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__290__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1378__ (
    .D(__542__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__291__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1379__ (
    .D(__683__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__292__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1380__ (
    .D(__586__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__293__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1381__ (
    .D(__786__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__294__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1382__ (
    .D(__609__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__295__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1383__ (
    .D(__678__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__296__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1384__ (
    .D(__838__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__297__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1385__ (
    .D(__787__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__298__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1386__ (
    .D(__971__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__299__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1387__ (
    .D(__1006__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__300__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1388__ (
    .D(__822__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__301__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1389__ (
    .D(__908__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__302__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1390__ (
    .D(__738__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__303__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1391__ (
    .D(__969__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__304__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1392__ (
    .D(__803__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__305__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1393__ (
    .D(__1013__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__306__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1394__ (
    .D(__907__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__307__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1395__ (
    .D(__849__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__308__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1396__ (
    .D(__973__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__309__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1397__ (
    .D(__1083__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__310__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1398__ (
    .D(__723__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__311__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1399__ (
    .D(__968__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__312__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1400__ (
    .D(__503__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__313__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1401__ (
    .D(__679__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__314__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1402__ (
    .D(__446__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__315__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1403__ (
    .D(__140__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__316__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1404__ (
    .D(__543__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__317__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1405__ (
    .D(__1038__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__318__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1406__ (
    .D(__978__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__319__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1407__ (
    .D(__235__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__320__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1408__ (
    .D(__238__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__321__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1409__ (
    .D(__305__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__322__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1410__ (
    .D(__576__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__323__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1411__ (
    .D(__15__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__324__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1412__ (
    .D(__537__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__325__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1413__ (
    .D(__475__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__326__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1414__ (
    .D(__762__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__327__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1415__ (
    .D(__1065__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__328__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1416__ (
    .D(__950__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__329__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1417__ (
    .D(__180__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__330__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1418__ (
    .D(__163__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__331__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1419__ (
    .D(__336__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__332__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1420__ (
    .D(__967__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__333__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1421__ (
    .D(__1016__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__334__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1422__ (
    .D(__783__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__335__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1423__ (
    .D(__369__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__336__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1424__ (
    .D(__491__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__337__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1425__ (
    .D(__1001__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__338__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1426__ (
    .D(__272__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__339__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1427__ (
    .D(__881__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__340__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1428__ (
    .D(__728__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__341__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1429__ (
    .D(__397__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__342__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1430__ (
    .D(__68__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__343__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1431__ (
    .D(__192__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__344__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1432__ (
    .D(__1067__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__345__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1433__ (
    .D(__1042__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__346__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1434__ (
    .D(__224__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__347__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1435__ (
    .D(__387__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__348__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1436__ (
    .D(__1007__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__349__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1437__ (
    .D(g1196),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__350__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1438__ (
    .D(__834__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__351__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1439__ (
    .D(__708__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__352__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1440__ (
    .D(__851__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__353__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1441__ (
    .D(__841__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__354__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1442__ (
    .D(__641__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__355__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1443__ (
    .D(__815__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__356__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1444__ (
    .D(__1082__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__357__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1445__ (
    .D(__844__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__358__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1446__ (
    .D(__961__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__359__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1447__ (
    .D(__164__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__360__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1448__ (
    .D(__764__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__361__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1449__ (
    .D(__702__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__362__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1450__ (
    .D(__436__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__363__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1451__ (
    .D(__260__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__364__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1452__ (
    .D(__763__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__365__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1453__ (
    .D(__989__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__366__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1454__ (
    .D(__843__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__367__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1455__ (
    .D(__765__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__368__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1456__ (
    .D(__265__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__369__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1457__ (
    .D(__805__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__370__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1458__ (
    .D(__782__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__371__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1459__ (
    .D(__884__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__372__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1460__ (
    .D(__1037__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__373__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1461__ (
    .D(__871__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__374__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1462__ (
    .D(__960__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__375__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1463__ (
    .D(__821__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__376__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1464__ (
    .D(__498__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__377__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1465__ (
    .D(__949__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__378__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1466__ (
    .D(__948__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__379__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1467__ (
    .D(__289__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__380__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1468__ (
    .D(__1029__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__381__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1469__ (
    .D(__744__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__382__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1470__ (
    .D(__737__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__383__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1471__ (
    .D(__999__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__384__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1472__ (
    .D(__866__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__385__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1473__ (
    .D(__147__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__386__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1474__ (
    .D(__564__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__387__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1475__ (
    .D(__997__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__388__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1476__ (
    .D(__239__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__389__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1477__ (
    .D(__820__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__390__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1478__ (
    .D(__958__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__391__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1479__ (
    .D(__894__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__392__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1480__ (
    .D(__944__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__393__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1481__ (
    .D(__904__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__394__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1482__ (
    .D(__266__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__395__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1483__ (
    .D(__1012__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__396__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1484__ (
    .D(g43),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__397__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1485__ (
    .D(__422__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__398__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1486__ (
    .D(__24__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__399__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1487__ (
    .D(__174__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__400__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1488__ (
    .D(g28),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__401__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1489__ (
    .D(__1041__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__402__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1490__ (
    .D(__731__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__403__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1491__ (
    .D(__882__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__404__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1492__ (
    .D(__657__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__405__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1493__ (
    .D(__695__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__406__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1494__ (
    .D(__347__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__407__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1495__ (
    .D(__873__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__408__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1496__ (
    .D(__890__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__409__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1497__ (
    .D(__35__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__410__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1498__ (
    .D(__865__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__411__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1499__ (
    .D(__1027__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__412__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1500__ (
    .D(__905__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__413__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1501__ (
    .D(__902__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__414__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1502__ (
    .D(__809__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__415__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1503__ (
    .D(__911__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__416__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1504__ (
    .D(__862__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__417__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1505__ (
    .D(__574__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__418__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1506__ (
    .D(__82__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__419__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1507__ (
    .D(__859__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__420__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1508__ (
    .D(__858__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__421__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1509__ (
    .D(__268__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__422__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1510__ (
    .D(__829__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__423__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1511__ (
    .D(__957__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__424__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1512__ (
    .D(__304__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__425__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1513__ (
    .D(__774__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__426__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1514__ (
    .D(__879__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__427__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1515__ (
    .D(g10),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__428__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1516__ (
    .D(__1078__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__429__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1517__ (
    .D(__755__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__430__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1518__ (
    .D(__715__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__431__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1519__ (
    .D(__44__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__432__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1520__ (
    .D(__1023__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__433__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1521__ (
    .D(__826__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__434__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1522__ (
    .D(__684__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__435__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1523__ (
    .D(__448__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__436__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1524__ (
    .D(__160__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__437__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1525__ (
    .D(__341__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__438__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1526__ (
    .D(__454__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__439__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1527__ (
    .D(__1054__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__440__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1528__ (
    .D(__712__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__441__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1529__ (
    .D(__842__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__442__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1530__ (
    .D(g1206),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__443__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1531__ (
    .D(__955__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__444__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1532__ (
    .D(__852__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__445__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1533__ (
    .D(__893__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__446__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1534__ (
    .D(__151__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__447__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1535__ (
    .D(__162__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__448__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1536__ (
    .D(__687__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__449__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1537__ (
    .D(__130__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__450__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1538__ (
    .D(__1076__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__451__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1539__ (
    .D(__267__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__452__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1540__ (
    .D(__814__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__453__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1541__ (
    .D(__405__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__454__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1542__ (
    .D(__444__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__455__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1543__ (
    .D(__1024__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__456__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1544__ (
    .D(__196__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__457__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1545__ (
    .D(__876__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__458__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1546__ (
    .D(__872__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__459__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1547__ (
    .D(__745__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__460__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1548__ (
    .D(__804__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__461__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1549__ (
    .D(__878__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__462__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1550__ (
    .D(__776__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__463__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1551__ (
    .D(__910__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__464__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1552__ (
    .D(__703__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__465__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1553__ (
    .D(__337__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__466__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1554__ (
    .D(__741__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__467__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1555__ (
    .D(__177__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__468__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1556__ (
    .D(__197__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__469__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1557__ (
    .D(__784__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__470__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1558__ (
    .D(__37__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__471__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1559__ (
    .D(__947__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__472__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1560__ (
    .D(__901__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__473__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1561__ (
    .D(__91__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__474__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1562__ (
    .D(g37),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__475__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1563__ (
    .D(__900__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__476__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1564__ (
    .D(__1069__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__477__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1565__ (
    .D(__167__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__478__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1566__ (
    .D(__345__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__479__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1567__ (
    .D(__889__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__480__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1568__ (
    .D(__233__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__481__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1569__ (
    .D(__930__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__482__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1570__ (
    .D(__761__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__483__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1571__ (
    .D(__443__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__484__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1572__ (
    .D(__77__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__485__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1573__ (
    .D(__730__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__486__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1574__ (
    .D(__817__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__487__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1575__ (
    .D(__580__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__488__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1576__ (
    .D(g1198),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__489__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1577__ (
    .D(__248__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__490__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1578__ (
    .D(__991__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__491__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1579__ (
    .D(__1031__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__492__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1580__ (
    .D(__759__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__493__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1581__ (
    .D(__134__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__494__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1582__ (
    .D(__544__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__495__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1583__ (
    .D(__581__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__496__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __1585__ (
    .I3(__74__),
    .I2(__489__),
    .I1(__377__),
    .I0(__253__),
    .O(__498__)
  );
  LUT6 #(
    .INIT(64'h8000000000000000)
  ) __1587__ (
    .I5(__444__),
    .I4(__134__),
    .I3(__35__),
    .I2(__260__),
    .I1(__220__),
    .I0(__205__),
    .O(__500__)
  );
  LUT5 #(
    .INIT(32'hff7fff80)
  ) __1588__ (
    .I4(__188__),
    .I3(__258__),
    .I2(__248__),
    .I1(__145__),
    .I0(__500__),
    .O(__501__)
  );
  LUT4 #(
    .INIT(16'h0100)
  ) __1589__ (
    .I3(__348__),
    .I2(__454__),
    .I1(__173__),
    .I0(__233__),
    .O(__502__)
  );
  LUT5 #(
    .INIT(32'h00000100)
  ) __1590__ (
    .I4(g42),
    .I3(g44),
    .I2(g41),
    .I1(__296__),
    .I0(g45),
    .O(__503__)
  );
  LUT4 #(
    .INIT(16'h0001)
  ) __1591__ (
    .I3(__156__),
    .I2(__197__),
    .I1(__272__),
    .I0(__222__),
    .O(__504__)
  );
  LUT5 #(
    .INIT(32'hcaaaaaaa)
  ) __1592__ (
    .I4(__504__),
    .I3(__503__),
    .I2(__502__),
    .I1(__72__),
    .I0(__259__),
    .O(__505__)
  );
  LUT3 #(
    .INIT(8'hbe)
  ) __1593__ (
    .I2(__145__),
    .I1(__500__),
    .I0(__258__),
    .O(__506__)
  );
  LUT4 #(
    .INIT(16'h8000)
  ) __1594__ (
    .I3(__230__),
    .I2(__293__),
    .I1(__335__),
    .I0(__383__),
    .O(__507__)
  );
  LUT4 #(
    .INIT(16'hf7f8)
  ) __1595__ (
    .I3(__33__),
    .I2(__332__),
    .I1(__507__),
    .I0(__66__),
    .O(__508__)
  );
  LUT4 #(
    .INIT(16'h0100)
  ) __1596__ (
    .I3(__233__),
    .I2(__348__),
    .I1(__454__),
    .I0(__173__),
    .O(__509__)
  );
  LUT6 #(
    .INIT(64'h8000000000000000)
  ) __1597__ (
    .I5(__156__),
    .I4(__197__),
    .I3(__272__),
    .I2(__222__),
    .I1(__509__),
    .I0(__215__),
    .O(__510__)
  );
  LUT2 #(
    .INIT(4'h7)
  ) __1598__ (
    .I1(__285__),
    .I0(__510__),
    .O(__511__)
  );
  LUT4 #(
    .INIT(16'h4000)
  ) __1599__ (
    .I3(__348__),
    .I2(__173__),
    .I1(__233__),
    .I0(__454__),
    .O(__512__)
  );
  LUT4 #(
    .INIT(16'h4000)
  ) __1600__ (
    .I3(__454__),
    .I2(__173__),
    .I1(__233__),
    .I0(__348__),
    .O(__513__)
  );
  LUT4 #(
    .INIT(16'h0040)
  ) __1601__ (
    .I3(__454__),
    .I2(__348__),
    .I1(__233__),
    .I0(__173__),
    .O(__514__)
  );
  LUT4 #(
    .INIT(16'h0040)
  ) __1602__ (
    .I3(__348__),
    .I2(__454__),
    .I1(__233__),
    .I0(__173__),
    .O(__515__)
  );
  LUT4 #(
    .INIT(16'h2777)
  ) __1603__ (
    .I3(__515__),
    .I2(__325__),
    .I1(__54__),
    .I0(__514__),
    .O(__516__)
  );
  LUT4 #(
    .INIT(16'h0001)
  ) __1604__ (
    .I3(__348__),
    .I2(__454__),
    .I1(__173__),
    .I0(__233__),
    .O(__517__)
  );
  LUT6 #(
    .INIT(64'h0000000000000040)
  ) __1605__ (
    .I5(__156__),
    .I4(__197__),
    .I3(__272__),
    .I2(__517__),
    .I1(__338__),
    .I0(__222__),
    .O(__518__)
  );
  LUT6 #(
    .INIT(64'h0000000007770000)
  ) __1606__ (
    .I5(__518__),
    .I4(__516__),
    .I3(__513__),
    .I2(__84__),
    .I1(__512__),
    .I0(__43__),
    .O(__519__)
  );
  LUT4 #(
    .INIT(16'h0100)
  ) __1607__ (
    .I3(__222__),
    .I2(__156__),
    .I1(__197__),
    .I0(__272__),
    .O(__520__)
  );
  LUT6 #(
    .INIT(64'h0000000080000000)
  ) __1608__ (
    .I5(__173__),
    .I4(__520__),
    .I3(__348__),
    .I2(__454__),
    .I1(__233__),
    .I0(__503__),
    .O(__521__)
  );
  LUT4 #(
    .INIT(16'h8000)
  ) __1609__ (
    .I3(__156__),
    .I2(__197__),
    .I1(__272__),
    .I0(__222__),
    .O(__522__)
  );
  LUT6 #(
    .INIT(64'h0000000000008000)
  ) __1610__ (
    .I5(__454__),
    .I4(__233__),
    .I3(__348__),
    .I2(__173__),
    .I1(__503__),
    .I0(__522__),
    .O(__523__)
  );
  LUT5 #(
    .INIT(32'h00004000)
  ) __1611__ (
    .I4(__348__),
    .I3(__173__),
    .I2(__233__),
    .I1(__297__),
    .I0(__454__),
    .O(__524__)
  );
  LUT5 #(
    .INIT(32'h00000040)
  ) __1612__ (
    .I4(__348__),
    .I3(__454__),
    .I2(__233__),
    .I1(g690),
    .I0(__173__),
    .O(__525__)
  );
  LUT6 #(
    .INIT(64'h0000000000000777)
  ) __1613__ (
    .I5(__525__),
    .I4(__524__),
    .I3(__523__),
    .I2(g751),
    .I1(__521__),
    .I0(__458__),
    .O(__526__)
  );
  LUT6 #(
    .INIT(64'h0000000000008000)
  ) __1614__ (
    .I5(__173__),
    .I4(__233__),
    .I3(__520__),
    .I2(__348__),
    .I1(__454__),
    .I0(__503__),
    .O(__527__)
  );
  LUT4 #(
    .INIT(16'hefff)
  ) __1615__ (
    .I3(__503__),
    .I2(__522__),
    .I1(__348__),
    .I0(__454__),
    .O(__528__)
  );
  LUT6 #(
    .INIT(64'hfffff7ffff77ffff)
  ) __1616__ (
    .I5(__348__),
    .I4(__454__),
    .I3(__173__),
    .I2(__233__),
    .I1(__503__),
    .I0(__522__),
    .O(__529__)
  );
  LUT4 #(
    .INIT(16'h0040)
  ) __1617__ (
    .I3(__521__),
    .I2(__529__),
    .I1(__528__),
    .I0(__527__),
    .O(__530__)
  );
  LUT5 #(
    .INIT(32'hc1ffffff)
  ) __1618__ (
    .I4(__520__),
    .I3(__503__),
    .I2(__348__),
    .I1(__454__),
    .I0(__173__),
    .O(__531__)
  );
  LUT5 #(
    .INIT(32'h00000777)
  ) __1619__ (
    .I4(__531__),
    .I3(__513__),
    .I2(__286__),
    .I1(__515__),
    .I0(__285__),
    .O(__532__)
  );
  LUT5 #(
    .INIT(32'h0000feff)
  ) __1620__ (
    .I4(__504__),
    .I3(__520__),
    .I2(__348__),
    .I1(__454__),
    .I0(__173__),
    .O(__533__)
  );
  LUT6 #(
    .INIT(64'h0000ff0fbbbbbbbb)
  ) __1621__ (
    .I5(__533__),
    .I4(__532__),
    .I3(__530__),
    .I2(__526__),
    .I1(__519__),
    .I0(__0__),
    .O(__534__)
  );
  LUT2 #(
    .INIT(4'hb)
  ) __1622__ (
    .I1(__313__),
    .I0(__534__),
    .O(__535__)
  );
  LUT4 #(
    .INIT(16'h0100)
  ) __1623__ (
    .I3(__454__),
    .I2(__348__),
    .I1(__173__),
    .I0(__233__),
    .O(__536__)
  );
  LUT5 #(
    .INIT(32'hcaaaaaaa)
  ) __1624__ (
    .I4(__504__),
    .I3(__503__),
    .I2(__536__),
    .I1(__38__),
    .I0(__325__),
    .O(__537__)
  );
  LUT3 #(
    .INIT(8'h06)
  ) __1625__ (
    .I2(__380__),
    .I1(__267__),
    .I0(__177__),
    .O(__538__)
  );
  LUT4 #(
    .INIT(16'h0708)
  ) __1626__ (
    .I3(__230__),
    .I2(__332__),
    .I1(__383__),
    .I0(__66__),
    .O(__539__)
  );
  LUT4 #(
    .INIT(16'h0040)
  ) __1627__ (
    .I3(__454__),
    .I2(__348__),
    .I1(__173__),
    .I0(__233__),
    .O(__540__)
  );
  LUT6 #(
    .INIT(64'h0000000000000040)
  ) __1628__ (
    .I5(__156__),
    .I4(__197__),
    .I3(__272__),
    .I2(__503__),
    .I1(__540__),
    .I0(__222__),
    .O(__541__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __1629__ (
    .I2(__541__),
    .I1(__456__),
    .I0(__291__),
    .O(__542__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __1630__ (
    .I1(__233__),
    .I0(__220__),
    .O(__543__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __1631__ (
    .I3(__484__),
    .I2(__443__),
    .I1(__495__),
    .I0(__479__),
    .O(__544__)
  );
  LUT3 #(
    .INIT(8'h1c)
  ) __1632__ (
    .I2(__462__),
    .I1(__334__),
    .I0(__131__),
    .O(__545__)
  );
  LUT2 #(
    .INIT(4'h7)
  ) __1633__ (
    .I1(__312__),
    .I0(__510__),
    .O(__546__)
  );
  LUT3 #(
    .INIT(8'hd5)
  ) __1634__ (
    .I2(__348__),
    .I1(__454__),
    .I0(__503__),
    .O(__547__)
  );
  LUT6 #(
    .INIT(64'hffffffffff35ffff)
  ) __1635__ (
    .I5(__348__),
    .I4(__454__),
    .I3(__173__),
    .I2(__233__),
    .I1(__204__),
    .I0(__495__),
    .O(__548__)
  );
  LUT5 #(
    .INIT(32'h2777ffff)
  ) __1636__ (
    .I4(__504__),
    .I3(__517__),
    .I2(__416__),
    .I1(__294__),
    .I0(__540__),
    .O(__549__)
  );
  LUT4 #(
    .INIT(16'h2777)
  ) __1637__ (
    .I3(__513__),
    .I2(__231__),
    .I1(__236__),
    .I0(__512__),
    .O(__550__)
  );
  LUT5 #(
    .INIT(32'h2777ffff)
  ) __1638__ (
    .I4(__504__),
    .I3(__509__),
    .I2(__105__),
    .I1(__218__),
    .I0(__502__),
    .O(__551__)
  );
  LUT5 #(
    .INIT(32'h00004000)
  ) __1639__ (
    .I4(__454__),
    .I3(__348__),
    .I2(__233__),
    .I1(__303__),
    .I0(__173__),
    .O(__552__)
  );
  LUT5 #(
    .INIT(32'h00000040)
  ) __1640__ (
    .I4(__348__),
    .I3(__454__),
    .I2(__173__),
    .I1(__195__),
    .I0(__233__),
    .O(__553__)
  );
  LUT6 #(
    .INIT(64'h0000000000008000)
  ) __1641__ (
    .I5(__553__),
    .I4(__552__),
    .I3(__551__),
    .I2(__550__),
    .I1(__549__),
    .I0(__548__),
    .O(__554__)
  );
  LUT5 #(
    .INIT(32'h00004000)
  ) __1642__ (
    .I4(__348__),
    .I3(__173__),
    .I2(__233__),
    .I1(__158__),
    .I0(__454__),
    .O(__555__)
  );
  LUT5 #(
    .INIT(32'h00000040)
  ) __1643__ (
    .I4(__348__),
    .I3(__454__),
    .I2(__173__),
    .I1(__323__),
    .I0(__233__),
    .O(__556__)
  );
  LUT5 #(
    .INIT(32'h00004000)
  ) __1644__ (
    .I4(__454__),
    .I3(__348__),
    .I2(__173__),
    .I1(g756),
    .I0(__233__),
    .O(__557__)
  );
  LUT6 #(
    .INIT(64'hffffffffffffff35)
  ) __1645__ (
    .I5(__348__),
    .I4(__454__),
    .I3(__173__),
    .I2(__233__),
    .I1(__142__),
    .I0(g702),
    .O(__558__)
  );
  LUT4 #(
    .INIT(16'h8000)
  ) __1646__ (
    .I3(__348__),
    .I2(__454__),
    .I1(__233__),
    .I0(__402__),
    .O(__559__)
  );
  LUT6 #(
    .INIT(64'h0000000000000040)
  ) __1647__ (
    .I5(__156__),
    .I4(__197__),
    .I3(__272__),
    .I2(__222__),
    .I1(__394__),
    .I0(__233__),
    .O(__560__)
  );
  LUT6 #(
    .INIT(64'h0000000000000100)
  ) __1648__ (
    .I5(__560__),
    .I4(__559__),
    .I3(__558__),
    .I2(__557__),
    .I1(__556__),
    .I0(__555__),
    .O(__561__)
  );
  LUT4 #(
    .INIT(16'h2777)
  ) __1649__ (
    .I3(__513__),
    .I2(__151__),
    .I1(__387__),
    .I0(__515__),
    .O(__562__)
  );
  LUT5 #(
    .INIT(32'h04040704)
  ) __1650__ (
    .I4(__514__),
    .I3(__562__),
    .I2(__531__),
    .I1(__512__),
    .I0(__128__),
    .O(__563__)
  );
  LUT6 #(
    .INIT(64'h0000ff0fbbbbbbbb)
  ) __1651__ (
    .I5(__533__),
    .I4(__563__),
    .I3(__530__),
    .I2(__561__),
    .I1(__554__),
    .I0(__547__),
    .O(__564__)
  );
  LUT2 #(
    .INIT(4'hb)
  ) __1652__ (
    .I1(__313__),
    .I0(__564__),
    .O(__565__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __1653__ (
    .I1(__156__),
    .I0(__444__),
    .O(__566__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __1654__ (
    .I3(__334__),
    .I2(__462__),
    .I1(__302__),
    .I0(__216__),
    .O(__567__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __1655__ (
    .I3(__419__),
    .I2(__82__),
    .I1(__112__),
    .I0(__191__),
    .O(__568__)
  );
  LUT5 #(
    .INIT(32'h80000000)
  ) __1656__ (
    .I4(__190__),
    .I3(__341__),
    .I2(__45__),
    .I1(__267__),
    .I0(__177__),
    .O(__569__)
  );
  LUT4 #(
    .INIT(16'h0708)
  ) __1657__ (
    .I3(__130__),
    .I2(__380__),
    .I1(__319__),
    .I0(__569__),
    .O(__570__)
  );
  LUT6 #(
    .INIT(64'h9009000000009009)
  ) __1658__ (
    .I5(__348__),
    .I4(__124__),
    .I3(__454__),
    .I2(__420__),
    .I1(__173__),
    .I0(__276__),
    .O(__571__)
  );
  LUT6 #(
    .INIT(64'h8100008100000000)
  ) __1659__ (
    .I5(__571__),
    .I4(__197__),
    .I3(__404__),
    .I2(__233__),
    .I1(__138__),
    .I0(__434__),
    .O(__572__)
  );
  LUT6 #(
    .INIT(64'h9009000000009009)
  ) __1660__ (
    .I5(__156__),
    .I4(__202__),
    .I3(__222__),
    .I2(__318__),
    .I1(__173__),
    .I0(__352__),
    .O(__573__)
  );
  LUT6 #(
    .INIT(64'h6ff6ffffffffffff)
  ) __1661__ (
    .I5(__573__),
    .I4(__572__),
    .I3(__272__),
    .I2(__440__),
    .I1(__348__),
    .I0(__108__),
    .O(__574__)
  );
  LUT6 #(
    .INIT(64'h0000000000004000)
  ) __1662__ (
    .I5(__348__),
    .I4(__454__),
    .I3(__173__),
    .I2(__522__),
    .I1(__215__),
    .I0(__233__),
    .O(__575__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __1663__ (
    .I2(__575__),
    .I1(__387__),
    .I0(__323__),
    .O(__576__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __1664__ (
    .I3(__484__),
    .I2(__443__),
    .I1(__38__),
    .I0(__490__),
    .O(__577__)
  );
  LUT6 #(
    .INIT(64'h8000000000000000)
  ) __1665__ (
    .I5(__33__),
    .I4(__372__),
    .I3(__230__),
    .I2(__293__),
    .I1(__335__),
    .I0(__383__),
    .O(__578__)
  );
  LUT4 #(
    .INIT(16'hf7f8)
  ) __1666__ (
    .I3(__14__),
    .I2(__332__),
    .I1(__578__),
    .I0(__66__),
    .O(__579__)
  );
  LUT4 #(
    .INIT(16'hefff)
  ) __1667__ (
    .I3(__35__),
    .I2(__205__),
    .I1(__134__),
    .I0(__260__),
    .O(__580__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __1668__ (
    .I3(__484__),
    .I2(__443__),
    .I1(__496__),
    .I0(__203__),
    .O(__581__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __1669__ (
    .I3(__386__),
    .I2(__147__),
    .I1(__218__),
    .I0(__479__),
    .O(__582__)
  );
  LUT6 #(
    .INIT(64'h0000000000004000)
  ) __1670__ (
    .I5(__156__),
    .I4(__197__),
    .I3(__222__),
    .I2(__512__),
    .I1(__215__),
    .I0(__272__),
    .O(__583__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __1671__ (
    .I2(__583__),
    .I1(__312__),
    .I0(__36__),
    .O(__584__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __1672__ (
    .I1(__30__),
    .I0(__321__),
    .O(__585__)
  );
  LUT5 #(
    .INIT(32'h007f0080)
  ) __1673__ (
    .I4(__293__),
    .I3(__332__),
    .I2(__230__),
    .I1(__383__),
    .I0(__66__),
    .O(__586__)
  );
  LUT5 #(
    .INIT(32'hff7fff80)
  ) __1674__ (
    .I4(__134__),
    .I3(__258__),
    .I2(__35__),
    .I1(__220__),
    .I0(__205__),
    .O(__587__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __1675__ (
    .I3(__386__),
    .I2(__147__),
    .I1(__166__),
    .I0(__364__),
    .O(__588__)
  );
  LUT4 #(
    .INIT(16'h2777)
  ) __1676__ (
    .I3(__515__),
    .I2(__56__),
    .I1(__259__),
    .I0(__514__),
    .O(__589__)
  );
  LUT5 #(
    .INIT(32'h2777ffff)
  ) __1677__ (
    .I4(__504__),
    .I3(__509__),
    .I2(__80__),
    .I1(__310__),
    .I0(__512__),
    .O(__590__)
  );
  LUT4 #(
    .INIT(16'h2777)
  ) __1678__ (
    .I3(__513__),
    .I2(__41__),
    .I1(__110__),
    .I0(__540__),
    .O(__591__)
  );
  LUT4 #(
    .INIT(16'h3dff)
  ) __1679__ (
    .I3(__173__),
    .I2(__348__),
    .I1(__454__),
    .I0(__233__),
    .O(__592__)
  );
  LUT4 #(
    .INIT(16'h0100)
  ) __1680__ (
    .I3(__173__),
    .I2(__348__),
    .I1(__454__),
    .I0(__233__),
    .O(__593__)
  );
  LUT5 #(
    .INIT(32'h2777ffff)
  ) __1681__ (
    .I4(__504__),
    .I3(__517__),
    .I2(__19__),
    .I1(__164__),
    .I0(__593__),
    .O(__594__)
  );
  LUT4 #(
    .INIT(16'h2777)
  ) __1682__ (
    .I3(__502__),
    .I2(__433__),
    .I1(__214__),
    .I0(__536__),
    .O(__595__)
  );
  LUT6 #(
    .INIT(64'h8000000000000000)
  ) __1683__ (
    .I5(__595__),
    .I4(__594__),
    .I3(__592__),
    .I2(__591__),
    .I1(__590__),
    .I0(__589__),
    .O(__596__)
  );
  LUT4 #(
    .INIT(16'h8000)
  ) __1684__ (
    .I3(__348__),
    .I2(__454__),
    .I1(__233__),
    .I0(__152__),
    .O(__597__)
  );
  LUT4 #(
    .INIT(16'h2777)
  ) __1685__ (
    .I3(__517__),
    .I2(g698),
    .I1(g757),
    .I0(__540__),
    .O(__598__)
  );
  LUT4 #(
    .INIT(16'h2777)
  ) __1686__ (
    .I3(__509__),
    .I2(g647),
    .I1(__275__),
    .I0(__515__),
    .O(__599__)
  );
  LUT5 #(
    .INIT(32'h00004000)
  ) __1687__ (
    .I4(__348__),
    .I3(__173__),
    .I2(__233__),
    .I1(__237__),
    .I0(__454__),
    .O(__600__)
  );
  LUT5 #(
    .INIT(32'h00000040)
  ) __1688__ (
    .I4(__348__),
    .I3(__454__),
    .I2(__173__),
    .I1(__246__),
    .I0(__233__),
    .O(__601__)
  );
  LUT6 #(
    .INIT(64'h0000000000000040)
  ) __1689__ (
    .I5(__156__),
    .I4(__197__),
    .I3(__272__),
    .I2(__222__),
    .I1(__301__),
    .I0(__233__),
    .O(__602__)
  );
  LUT6 #(
    .INIT(64'h0000000000000040)
  ) __1690__ (
    .I5(__602__),
    .I4(__601__),
    .I3(__600__),
    .I2(__599__),
    .I1(__598__),
    .I0(__597__),
    .O(__603__)
  );
  LUT4 #(
    .INIT(16'h2777)
  ) __1691__ (
    .I3(__513__),
    .I2(__447__),
    .I1(__89__),
    .I0(__512__),
    .O(__604__)
  );
  LUT4 #(
    .INIT(16'h0040)
  ) __1692__ (
    .I3(__348__),
    .I2(__173__),
    .I1(__233__),
    .I0(__454__),
    .O(__605__)
  );
  LUT5 #(
    .INIT(32'h00000700)
  ) __1693__ (
    .I4(__605__),
    .I3(__604__),
    .I2(__531__),
    .I1(__515__),
    .I0(__216__),
    .O(__606__)
  );
  LUT6 #(
    .INIT(64'h0000ff0fbbbbbbbb)
  ) __1694__ (
    .I5(__533__),
    .I4(__606__),
    .I3(__530__),
    .I2(__603__),
    .I1(__596__),
    .I0(__0__),
    .O(__607__)
  );
  LUT2 #(
    .INIT(4'hb)
  ) __1695__ (
    .I1(__313__),
    .I0(__607__),
    .O(__608__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __1696__ (
    .I3(__386__),
    .I2(__147__),
    .I1(__295__),
    .I0(__109__),
    .O(__609__)
  );
  LUT5 #(
    .INIT(32'h00000100)
  ) __1697__ (
    .I4(__156__),
    .I3(__509__),
    .I2(__197__),
    .I1(__272__),
    .I0(__222__),
    .O(__610__)
  );
  LUT5 #(
    .INIT(32'h2777ffff)
  ) __1698__ (
    .I4(__504__),
    .I3(__517__),
    .I2(__493__),
    .I1(__217__),
    .I0(__515__),
    .O(__611__)
  );
  LUT4 #(
    .INIT(16'h2777)
  ) __1699__ (
    .I3(__514__),
    .I2(__368__),
    .I1(__86__),
    .I0(__512__),
    .O(__612__)
  );
  LUT6 #(
    .INIT(64'h153f000000000000)
  ) __1700__ (
    .I5(__612__),
    .I4(__611__),
    .I3(__513__),
    .I2(__610__),
    .I1(__428__),
    .I0(__209__),
    .O(__613__)
  );
  LUT5 #(
    .INIT(32'h00000040)
  ) __1701__ (
    .I4(__348__),
    .I3(__454__),
    .I2(__233__),
    .I1(g633),
    .I0(__173__),
    .O(__614__)
  );
  LUT5 #(
    .INIT(32'h00004000)
  ) __1702__ (
    .I4(__348__),
    .I3(__173__),
    .I2(__233__),
    .I1(__94__),
    .I0(__454__),
    .O(__615__)
  );
  LUT6 #(
    .INIT(64'h0000000000000777)
  ) __1703__ (
    .I5(__615__),
    .I4(__614__),
    .I3(__523__),
    .I2(g755),
    .I1(__521__),
    .I0(__329__),
    .O(__616__)
  );
  LUT5 #(
    .INIT(32'h00000777)
  ) __1704__ (
    .I4(__531__),
    .I3(__513__),
    .I2(__135__),
    .I1(__515__),
    .I0(__73__),
    .O(__617__)
  );
  LUT6 #(
    .INIT(64'h0000ff0fbbbbbbbb)
  ) __1705__ (
    .I5(__533__),
    .I4(__617__),
    .I3(__530__),
    .I2(__616__),
    .I1(__613__),
    .I0(__0__),
    .O(__618__)
  );
  LUT4 #(
    .INIT(16'h2777)
  ) __1706__ (
    .I3(__514__),
    .I2(__278__),
    .I1(__291__),
    .I0(__512__),
    .O(__619__)
  );
  LUT5 #(
    .INIT(32'h2777ffff)
  ) __1707__ (
    .I4(__504__),
    .I3(__517__),
    .I2(__431__),
    .I1(__362__),
    .I0(__515__),
    .O(__620__)
  );
  LUT6 #(
    .INIT(64'h153f000000000000)
  ) __1708__ (
    .I5(__620__),
    .I4(__619__),
    .I3(__513__),
    .I2(__63__),
    .I1(__610__),
    .I0(__408__),
    .O(__621__)
  );
  LUT5 #(
    .INIT(32'h00004000)
  ) __1709__ (
    .I4(__348__),
    .I3(__173__),
    .I2(__233__),
    .I1(__168__),
    .I0(__454__),
    .O(__622__)
  );
  LUT5 #(
    .INIT(32'h00000040)
  ) __1710__ (
    .I4(__348__),
    .I3(__454__),
    .I2(__233__),
    .I1(g634),
    .I0(__173__),
    .O(__623__)
  );
  LUT6 #(
    .INIT(64'h0000000000000777)
  ) __1711__ (
    .I5(__623__),
    .I4(__622__),
    .I3(__523__),
    .I2(g754),
    .I1(__521__),
    .I0(__184__),
    .O(__624__)
  );
  LUT5 #(
    .INIT(32'h00000777)
  ) __1712__ (
    .I4(__531__),
    .I3(__513__),
    .I2(__23__),
    .I1(__515__),
    .I0(__79__),
    .O(__625__)
  );
  LUT6 #(
    .INIT(64'h0000ff0fbbbbbbbb)
  ) __1713__ (
    .I5(__533__),
    .I4(__625__),
    .I3(__530__),
    .I2(__624__),
    .I1(__621__),
    .I0(__0__),
    .O(__626__)
  );
  LUT4 #(
    .INIT(16'h8000)
  ) __1714__ (
    .I3(__348__),
    .I2(__454__),
    .I1(__233__),
    .I0(__396__),
    .O(__627__)
  );
  LUT6 #(
    .INIT(64'h0000000000000040)
  ) __1715__ (
    .I5(__156__),
    .I4(__197__),
    .I3(__272__),
    .I2(__222__),
    .I1(__67__),
    .I0(__233__),
    .O(__628__)
  );
  LUT6 #(
    .INIT(64'hffffffffffffff35)
  ) __1716__ (
    .I5(__348__),
    .I4(__454__),
    .I3(__173__),
    .I2(__233__),
    .I1(g635),
    .I0(g723),
    .O(__629__)
  );
  LUT4 #(
    .INIT(16'h2777)
  ) __1717__ (
    .I3(__593__),
    .I2(__298__),
    .I1(__143__),
    .I0(__605__),
    .O(__630__)
  );
  LUT6 #(
    .INIT(64'h0007000000000000)
  ) __1718__ (
    .I5(__630__),
    .I4(__629__),
    .I3(__628__),
    .I2(__627__),
    .I1(__523__),
    .I0(g752),
    .O(__631__)
  );
  LUT5 #(
    .INIT(32'h2777ffff)
  ) __1719__ (
    .I4(__504__),
    .I3(__517__),
    .I2(__194__),
    .I1(__95__),
    .I0(__593__),
    .O(__632__)
  );
  LUT4 #(
    .INIT(16'h2777)
  ) __1720__ (
    .I3(__509__),
    .I2(__315__),
    .I1(__123__),
    .I0(__502__),
    .O(__633__)
  );
  LUT4 #(
    .INIT(16'h2777)
  ) __1721__ (
    .I3(__540__),
    .I2(__114__),
    .I1(__459__),
    .I0(__512__),
    .O(__634__)
  );
  LUT4 #(
    .INIT(16'h2777)
  ) __1722__ (
    .I3(__513__),
    .I2(__467__),
    .I1(__421__),
    .I0(__536__),
    .O(__635__)
  );
  LUT4 #(
    .INIT(16'h2777)
  ) __1723__ (
    .I3(__520__),
    .I2(__509__),
    .I1(__57__),
    .I0(__514__),
    .O(__636__)
  );
  LUT5 #(
    .INIT(32'h00004000)
  ) __1724__ (
    .I4(__348__),
    .I3(__454__),
    .I2(__233__),
    .I1(__155__),
    .I0(__173__),
    .O(__637__)
  );
  LUT6 #(
    .INIT(64'h0000000080000000)
  ) __1725__ (
    .I5(__637__),
    .I4(__636__),
    .I3(__635__),
    .I2(__634__),
    .I1(__633__),
    .I0(__632__),
    .O(__638__)
  );
  LUT4 #(
    .INIT(16'hfdf7)
  ) __1726__ (
    .I3(__348__),
    .I2(__454__),
    .I1(__173__),
    .I0(__233__),
    .O(__639__)
  );
  LUT6 #(
    .INIT(64'h0000000015370404)
  ) __1727__ (
    .I5(__531__),
    .I4(__639__),
    .I3(__213__),
    .I2(__355__),
    .I1(__515__),
    .I0(__513__),
    .O(__640__)
  );
  LUT6 #(
    .INIT(64'haaffaabbaaafaaab)
  ) __1728__ (
    .I5(__533__),
    .I4(__530__),
    .I3(__640__),
    .I2(__638__),
    .I1(__631__),
    .I0(__0__),
    .O(__641__)
  );
  LUT4 #(
    .INIT(16'h6996)
  ) __1729__ (
    .I3(__641__),
    .I2(__626__),
    .I1(__534__),
    .I0(__618__),
    .O(__642__)
  );
  LUT5 #(
    .INIT(32'h2777ffff)
  ) __1730__ (
    .I4(__504__),
    .I3(__509__),
    .I2(__247__),
    .I1(__442__),
    .I0(__512__),
    .O(__643__)
  );
  LUT4 #(
    .INIT(16'h2777)
  ) __1731__ (
    .I3(__515__),
    .I2(__414__),
    .I1(__439__),
    .I0(__593__),
    .O(__644__)
  );
  LUT4 #(
    .INIT(16'h2777)
  ) __1732__ (
    .I3(__513__),
    .I2(__193__),
    .I1(__125__),
    .I0(__536__),
    .O(__645__)
  );
  LUT4 #(
    .INIT(16'h2777)
  ) __1733__ (
    .I3(__502__),
    .I2(__353__),
    .I1(__349__),
    .I0(__514__),
    .O(__646__)
  );
  LUT5 #(
    .INIT(32'h2777ffff)
  ) __1734__ (
    .I4(__504__),
    .I3(__517__),
    .I2(__281__),
    .I1(__435__),
    .I0(__540__),
    .O(__647__)
  );
  LUT5 #(
    .INIT(32'h80000000)
  ) __1735__ (
    .I4(__647__),
    .I3(__646__),
    .I2(__645__),
    .I1(__644__),
    .I0(__643__),
    .O(__648__)
  );
  LUT5 #(
    .INIT(32'h00004000)
  ) __1736__ (
    .I4(__348__),
    .I3(__173__),
    .I2(__233__),
    .I1(__206__),
    .I0(__454__),
    .O(__649__)
  );
  LUT5 #(
    .INIT(32'h00000100)
  ) __1737__ (
    .I4(__348__),
    .I3(g722),
    .I2(__454__),
    .I1(__173__),
    .I0(__233__),
    .O(__650__)
  );
  LUT5 #(
    .INIT(32'h00004000)
  ) __1738__ (
    .I4(__454__),
    .I3(__348__),
    .I2(__173__),
    .I1(g753),
    .I0(__233__),
    .O(__651__)
  );
  LUT4 #(
    .INIT(16'h2777)
  ) __1739__ (
    .I3(__509__),
    .I2(g645),
    .I1(__328__),
    .I0(__593__),
    .O(__652__)
  );
  LUT4 #(
    .INIT(16'h8000)
  ) __1740__ (
    .I3(__348__),
    .I2(__454__),
    .I1(__233__),
    .I0(__367__),
    .O(__653__)
  );
  LUT6 #(
    .INIT(64'h0000000000000040)
  ) __1741__ (
    .I5(__156__),
    .I4(__197__),
    .I3(__272__),
    .I2(__222__),
    .I1(__161__),
    .I0(__233__),
    .O(__654__)
  );
  LUT6 #(
    .INIT(64'h0000000000000100)
  ) __1742__ (
    .I5(__654__),
    .I4(__653__),
    .I3(__652__),
    .I2(__651__),
    .I1(__650__),
    .I0(__649__),
    .O(__655__)
  );
  LUT5 #(
    .INIT(32'h00000777)
  ) __1743__ (
    .I4(__531__),
    .I3(__513__),
    .I2(__200__),
    .I1(__515__),
    .I0(__405__),
    .O(__656__)
  );
  LUT6 #(
    .INIT(64'h0000ff0fbbbbbbbb)
  ) __1744__ (
    .I5(__533__),
    .I4(__656__),
    .I3(__530__),
    .I2(__655__),
    .I1(__648__),
    .I0(__547__),
    .O(__657__)
  );
  LUT6 #(
    .INIT(64'h0000000000004000)
  ) __1745__ (
    .I5(__348__),
    .I4(__454__),
    .I3(__173__),
    .I2(__503__),
    .I1(__522__),
    .I0(__233__),
    .O(__658__)
  );
  LUT4 #(
    .INIT(16'h2777)
  ) __1746__ (
    .I3(__333__),
    .I2(__521__),
    .I1(__477__),
    .I0(__605__),
    .O(__659__)
  );
  LUT6 #(
    .INIT(64'h0777ffffffffffff)
  ) __1747__ (
    .I5(__503__),
    .I4(__522__),
    .I3(__515__),
    .I2(__170__),
    .I1(__509__),
    .I0(g648),
    .O(__660__)
  );
  LUT5 #(
    .INIT(32'h27227722)
  ) __1748__ (
    .I4(__517__),
    .I3(__660__),
    .I2(g694),
    .I1(g49),
    .I0(__523__),
    .O(__661__)
  );
  LUT6 #(
    .INIT(64'h153f000000000000)
  ) __1749__ (
    .I5(__661__),
    .I4(__659__),
    .I3(__299__),
    .I2(__470__),
    .I1(__527__),
    .I0(__658__),
    .O(__662__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __1750__ (
    .I5(__52__),
    .I4(__513__),
    .I3(__515__),
    .I2(__312__),
    .I1(__36__),
    .I0(__512__),
    .O(__663__)
  );
  LUT6 #(
    .INIT(64'h4444440444440444)
  ) __1751__ (
    .I5(__348__),
    .I4(__454__),
    .I3(__173__),
    .I2(__233__),
    .I1(__663__),
    .I0(__531__),
    .O(__664__)
  );
  LUT6 #(
    .INIT(64'h0000000000000040)
  ) __1752__ (
    .I5(__156__),
    .I4(__197__),
    .I3(__272__),
    .I2(__503__),
    .I1(__536__),
    .I0(__222__),
    .O(__665__)
  );
  LUT3 #(
    .INIT(8'h7f)
  ) __1753__ (
    .I2(__348__),
    .I1(__454__),
    .I0(__233__),
    .O(__666__)
  );
  LUT5 #(
    .INIT(32'hfff5fff7)
  ) __1754__ (
    .I4(__520__),
    .I3(__348__),
    .I2(__454__),
    .I1(__173__),
    .I0(__233__),
    .O(__667__)
  );
  LUT6 #(
    .INIT(64'h153f000000000000)
  ) __1755__ (
    .I5(__667__),
    .I4(__666__),
    .I3(__100__),
    .I2(__241__),
    .I1(__665__),
    .I0(__541__),
    .O(__668__)
  );
  LUT6 #(
    .INIT(64'h0000000000000040)
  ) __1756__ (
    .I5(__156__),
    .I4(__197__),
    .I3(__272__),
    .I2(__503__),
    .I1(__502__),
    .I0(__222__),
    .O(__669__)
  );
  LUT5 #(
    .INIT(32'h2777ffff)
  ) __1757__ (
    .I4(__504__),
    .I3(__304__),
    .I2(__517__),
    .I1(__481__),
    .I0(__593__),
    .O(__670__)
  );
  LUT5 #(
    .INIT(32'h07770000)
  ) __1758__ (
    .I4(__670__),
    .I3(__512__),
    .I2(__392__),
    .I1(__669__),
    .I0(__60__),
    .O(__671__)
  );
  LUT4 #(
    .INIT(16'h2777)
  ) __1759__ (
    .I3(__270__),
    .I2(__509__),
    .I1(__159__),
    .I0(__514__),
    .O(__672__)
  );
  LUT4 #(
    .INIT(16'h2777)
  ) __1760__ (
    .I3(__513__),
    .I2(__69__),
    .I1(__351__),
    .I0(__515__),
    .O(__673__)
  );
  LUT6 #(
    .INIT(64'h00000000bfffffff)
  ) __1761__ (
    .I5(__533__),
    .I4(__673__),
    .I3(__672__),
    .I2(__671__),
    .I1(__668__),
    .I0(__0__),
    .O(__674__)
  );
  LUT6 #(
    .INIT(64'h0000f2ffffff0d00)
  ) __1762__ (
    .I5(__607__),
    .I4(__674__),
    .I3(__533__),
    .I2(__664__),
    .I1(__530__),
    .I0(__662__),
    .O(__675__)
  );
  LUT3 #(
    .INIT(8'hb0)
  ) __1763__ (
    .I2(__314__),
    .I1(g44),
    .I0(g45),
    .O(__676__)
  );
  LUT4 #(
    .INIT(16'h9669)
  ) __1764__ (
    .I3(__312__),
    .I2(__405__),
    .I1(__216__),
    .I0(__387__),
    .O(__677__)
  );
  LUT6 #(
    .INIT(64'h6996966996696996)
  ) __1765__ (
    .I5(__355__),
    .I4(__79__),
    .I3(__285__),
    .I2(__73__),
    .I1(__677__),
    .I0(__676__),
    .O(__678__)
  );
  LUT6 #(
    .INIT(64'h96699669ffff0000)
  ) __1766__ (
    .I5(g44),
    .I4(__678__),
    .I3(__675__),
    .I2(__564__),
    .I1(__657__),
    .I0(__642__),
    .O(__679__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __1767__ (
    .I2(__541__),
    .I1(__104__),
    .I0(__236__),
    .O(__680__)
  );
  LUT2 #(
    .INIT(4'h7)
  ) __1768__ (
    .I1(__405__),
    .I0(__510__),
    .O(__681__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __1769__ (
    .I3(__386__),
    .I2(__147__),
    .I1(__26__),
    .I0(__490__),
    .O(__682__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __1770__ (
    .I3(__419__),
    .I2(__82__),
    .I1(__292__),
    .I0(__109__),
    .O(__683__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __1771__ (
    .I3(__74__),
    .I2(__489__),
    .I1(__435__),
    .I0(__256__),
    .O(__684__)
  );
  LUT3 #(
    .INIT(8'hf1)
  ) __1772__ (
    .I2(g45),
    .I1(__313__),
    .I0(__284__),
    .O(__685__)
  );
  LUT4 #(
    .INIT(16'hf7f8)
  ) __1773__ (
    .I3(__248__),
    .I2(__258__),
    .I1(__145__),
    .I0(__500__),
    .O(__686__)
  );
  LUT4 #(
    .INIT(16'h4f10)
  ) __1774__ (
    .I3(__449__),
    .I2(__261__),
    .I1(__255__),
    .I0(__472__),
    .O(__687__)
  );
  LUT6 #(
    .INIT(64'h8000000000000000)
  ) __1775__ (
    .I5(__115__),
    .I4(__374__),
    .I3(__29__),
    .I2(__307__),
    .I1(__412__),
    .I0(__464__),
    .O(__688__)
  );
  LUT6 #(
    .INIT(64'h0000000080000000)
  ) __1776__ (
    .I5(__255__),
    .I4(__129__),
    .I3(__244__),
    .I2(__25__),
    .I1(__280__),
    .I0(__688__),
    .O(__689__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __1777__ (
    .I1(__431__),
    .I0(__87__),
    .O(__690__)
  );
  LUT6 #(
    .INIT(64'h0000000000008000)
  ) __1778__ (
    .I5(__255__),
    .I4(__690__),
    .I3(__141__),
    .I2(__129__),
    .I1(__244__),
    .I0(__25__),
    .O(__691__)
  );
  LUT4 #(
    .INIT(16'h8000)
  ) __1779__ (
    .I3(__115__),
    .I2(__374__),
    .I1(__29__),
    .I0(__307__),
    .O(__692__)
  );
  LUT6 #(
    .INIT(64'h88f0000000000000)
  ) __1780__ (
    .I5(__692__),
    .I4(__691__),
    .I3(__194__),
    .I2(__280__),
    .I1(__406__),
    .I0(__412__),
    .O(__693__)
  );
  LUT5 #(
    .INIT(32'h0f0f090f)
  ) __1781__ (
    .I4(__87__),
    .I3(__431__),
    .I2(__693__),
    .I1(__326__),
    .I0(__475__),
    .O(__694__)
  );
  LUT4 #(
    .INIT(16'h7800)
  ) __1782__ (
    .I3(__694__),
    .I2(__406__),
    .I1(__141__),
    .I0(__689__),
    .O(__695__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __1783__ (
    .I3(__386__),
    .I2(__147__),
    .I1(__123__),
    .I0(__485__),
    .O(__696__)
  );
  LUT6 #(
    .INIT(64'h8000000000000000)
  ) __1784__ (
    .I5(__441__),
    .I4(__75__),
    .I3(__245__),
    .I2(__250__),
    .I1(__53__),
    .I0(__449__),
    .O(__697__)
  );
  LUT6 #(
    .INIT(64'h4f5f5f5f10000000)
  ) __1785__ (
    .I5(__187__),
    .I4(__361__),
    .I3(__697__),
    .I2(__261__),
    .I1(__255__),
    .I0(__472__),
    .O(__698__)
  );
  LUT4 #(
    .INIT(16'h0230)
  ) __1786__ (
    .I3(__48__),
    .I2(__62__),
    .I1(__146__),
    .I0(__46__),
    .O(__699__)
  );
  LUT6 #(
    .INIT(64'h0000000080000000)
  ) __1787__ (
    .I5(__255__),
    .I4(__75__),
    .I3(__245__),
    .I2(__250__),
    .I1(__449__),
    .I0(__261__),
    .O(__700__)
  );
  LUT4 #(
    .INIT(16'h152a)
  ) __1788__ (
    .I3(__53__),
    .I2(__261__),
    .I1(__472__),
    .I0(__700__),
    .O(__701__)
  );
  LUT5 #(
    .INIT(32'hcaaaaaaa)
  ) __1789__ (
    .I4(__504__),
    .I3(__503__),
    .I2(__536__),
    .I1(__376__),
    .I0(__362__),
    .O(__702__)
  );
  LUT5 #(
    .INIT(32'hff808080)
  ) __1790__ (
    .I4(__91__),
    .I3(__411__),
    .I2(__122__),
    .I1(__261__),
    .I0(__142__),
    .O(__703__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __1791__ (
    .I2(__40__),
    .I1(__92__),
    .I0(g929),
    .O(__704__)
  );
  LUT6 #(
    .INIT(64'h8000000000000000)
  ) __1792__ (
    .I5(__345__),
    .I4(__167__),
    .I3(__188__),
    .I2(__248__),
    .I1(__145__),
    .I0(__500__),
    .O(__705__)
  );
  LUT5 #(
    .INIT(32'hbfeaaaaa)
  ) __1793__ (
    .I4(__103__),
    .I3(__77__),
    .I2(__300__),
    .I1(__705__),
    .I0(__258__),
    .O(__706__)
  );
  LUT6 #(
    .INIT(64'h8000000000000000)
  ) __1794__ (
    .I5(__124__),
    .I4(__318__),
    .I3(__420__),
    .I2(__202__),
    .I1(__276__),
    .I0(__434__),
    .O(__707__)
  );
  LUT6 #(
    .INIT(64'h7fff800000000000)
  ) __1795__ (
    .I5(__391__),
    .I4(__352__),
    .I3(__138__),
    .I2(__440__),
    .I1(__404__),
    .I0(__707__),
    .O(__708__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __1796__ (
    .I1(__222__),
    .I0(__77__),
    .O(__709__)
  );
  LUT6 #(
    .INIT(64'h8000000000000000)
  ) __1797__ (
    .I5(__156__),
    .I4(__197__),
    .I3(__272__),
    .I2(__222__),
    .I1(__517__),
    .I0(__215__),
    .O(__710__)
  );
  LUT2 #(
    .INIT(4'h7)
  ) __1798__ (
    .I1(__387__),
    .I0(__710__),
    .O(__711__)
  );
  LUT5 #(
    .INIT(32'h134c5f00)
  ) __1799__ (
    .I4(__53__),
    .I3(__441__),
    .I2(__261__),
    .I1(__700__),
    .I0(__472__),
    .O(__712__)
  );
  LUT3 #(
    .INIT(8'hbe)
  ) __1800__ (
    .I2(__220__),
    .I1(__205__),
    .I0(__258__),
    .O(__713__)
  );
  LUT2 #(
    .INIT(4'h7)
  ) __1801__ (
    .I1(__387__),
    .I0(__510__),
    .O(__714__)
  );
  LUT5 #(
    .INIT(32'hcaaaaaaa)
  ) __1802__ (
    .I4(__504__),
    .I3(__517__),
    .I2(__215__),
    .I1(__79__),
    .I0(__431__),
    .O(__715__)
  );
  LUT6 #(
    .INIT(64'h9009000000009009)
  ) __1803__ (
    .I5(__156__),
    .I4(__130__),
    .I3(__272__),
    .I2(__279__),
    .I1(__454__),
    .I0(__190__),
    .O(__716__)
  );
  LUT6 #(
    .INIT(64'h9009000000009009)
  ) __1804__ (
    .I5(__197__),
    .I4(__185__),
    .I3(__348__),
    .I2(__341__),
    .I1(__173__),
    .I0(__45__),
    .O(__717__)
  );
  LUT6 #(
    .INIT(64'h6ff6ffffffffffff)
  ) __1805__ (
    .I5(__717__),
    .I4(__716__),
    .I3(__222__),
    .I2(__319__),
    .I1(__233__),
    .I0(__267__),
    .O(__718__)
  );
  LUT6 #(
    .INIT(64'h8000000000000000)
  ) __1806__ (
    .I5(__156__),
    .I4(__197__),
    .I3(__272__),
    .I2(__222__),
    .I1(__605__),
    .I0(__215__),
    .O(__719__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __1807__ (
    .I2(__719__),
    .I1(__355__),
    .I0(__143__),
    .O(__720__)
  );
  LUT3 #(
    .INIT(8'h40)
  ) __1808__ (
    .I2(__697__),
    .I1(__261__),
    .I0(__255__),
    .O(__721__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __1809__ (
    .I1(__261__),
    .I0(__472__),
    .O(__722__)
  );
  LUT6 #(
    .INIT(64'h00007fff00008000)
  ) __1810__ (
    .I5(__311__),
    .I4(__722__),
    .I3(__232__),
    .I2(__361__),
    .I1(__187__),
    .I0(__721__),
    .O(__723__)
  );
  LUT5 #(
    .INIT(32'h00007800)
  ) __1811__ (
    .I4(__258__),
    .I3(__103__),
    .I2(__35__),
    .I1(__220__),
    .I0(__205__),
    .O(__724__)
  );
  LUT3 #(
    .INIT(8'h01)
  ) __1812__ (
    .I2(g42),
    .I1(g41),
    .I0(g45),
    .O(__725__)
  );
  LUT6 #(
    .INIT(64'h8000000000000000)
  ) __1813__ (
    .I5(__156__),
    .I4(__197__),
    .I3(__272__),
    .I2(__222__),
    .I1(__515__),
    .I0(__215__),
    .O(__726__)
  );
  LUT6 #(
    .INIT(64'hffff0000ff40ff40)
  ) __1814__ (
    .I5(__726__),
    .I4(__216__),
    .I3(__275__),
    .I2(__678__),
    .I1(__725__),
    .I0(g44),
    .O(__727__)
  );
  LUT5 #(
    .INIT(32'h007f0080)
  ) __1815__ (
    .I4(__341__),
    .I3(__380__),
    .I2(__45__),
    .I1(__267__),
    .I0(__177__),
    .O(__728__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __1816__ (
    .I1(__222__),
    .I0(__260__),
    .O(__729__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __1817__ (
    .I3(__74__),
    .I2(__489__),
    .I1(__486__),
    .I0(__191__),
    .O(__730__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __1818__ (
    .I3(__386__),
    .I2(__147__),
    .I1(__403__),
    .I0(__494__),
    .O(__731__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __1819__ (
    .I3(__419__),
    .I2(__82__),
    .I1(__127__),
    .I0(__455__),
    .O(__732__)
  );
  LUT3 #(
    .INIT(8'h60)
  ) __1820__ (
    .I2(__694__),
    .I1(__141__),
    .I0(__689__),
    .O(__733__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __1821__ (
    .I1(__101__),
    .I0(__324__),
    .O(__734__)
  );
  LUT5 #(
    .INIT(32'hcaaaaaaa)
  ) __1822__ (
    .I4(__504__),
    .I3(__503__),
    .I2(__536__),
    .I1(__271__),
    .I0(__204__),
    .O(__735__)
  );
  LUT3 #(
    .INIT(8'hae)
  ) __1823__ (
    .I2(__87__),
    .I1(__281__),
    .I0(__389__),
    .O(__736__)
  );
  LUT3 #(
    .INIT(8'h06)
  ) __1824__ (
    .I2(__332__),
    .I1(__383__),
    .I0(__66__),
    .O(__737__)
  );
  LUT5 #(
    .INIT(32'hcaaaaaaa)
  ) __1825__ (
    .I4(__504__),
    .I3(__503__),
    .I2(__502__),
    .I1(__102__),
    .I0(__303__),
    .O(__738__)
  );
  LUT5 #(
    .INIT(32'hffff9aaa)
  ) __1826__ (
    .I4(__146__),
    .I3(__48__),
    .I2(__62__),
    .I1(__107__),
    .I0(__172__),
    .O(__739__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __1827__ (
    .I1(g43),
    .I0(__19__),
    .O(__740__)
  );
  LUT5 #(
    .INIT(32'hcaaaaaaa)
  ) __1828__ (
    .I4(__504__),
    .I3(__503__),
    .I2(__536__),
    .I1(__496__),
    .I0(__467__),
    .O(__741__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __1829__ (
    .I2(__669__),
    .I1(__375__),
    .I0(__278__),
    .O(__742__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __1830__ (
    .I2(__665__),
    .I1(__76__),
    .I0(__69__),
    .O(__743__)
  );
  LUT4 #(
    .INIT(16'h001c)
  ) __1831__ (
    .I3(__177__),
    .I2(__382__),
    .I1(__393__),
    .I0(__282__),
    .O(__744__)
  );
  LUT5 #(
    .INIT(32'haaaa3fc0)
  ) __1832__ (
    .I4(__322__),
    .I3(__460__),
    .I2(__182__),
    .I1(__157__),
    .I0(__195__),
    .O(__745__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __1833__ (
    .I3(__334__),
    .I2(__462__),
    .I1(__111__),
    .I0(__312__),
    .O(__746__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __1834__ (
    .I1(g698),
    .I0(__246__),
    .O(__747__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __1835__ (
    .I5(g694),
    .I4(__299__),
    .I3(g634),
    .I2(__168__),
    .I1(__94__),
    .I0(g633),
    .O(__748__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __1836__ (
    .I1(__143__),
    .I0(g635),
    .O(__749__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __1837__ (
    .I1(g702),
    .I0(__323__),
    .O(__750__)
  );
  LUT6 #(
    .INIT(64'h0000000000000700)
  ) __1838__ (
    .I5(__750__),
    .I4(__749__),
    .I3(__748__),
    .I2(__747__),
    .I1(__328__),
    .I0(g722),
    .O(__751__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __1839__ (
    .I1(__158__),
    .I0(__142__),
    .O(__752__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __1840__ (
    .I1(g647),
    .I0(__237__),
    .O(__753__)
  );
  LUT6 #(
    .INIT(64'h0000000000000777)
  ) __1841__ (
    .I5(__753__),
    .I4(__752__),
    .I3(g648),
    .I2(__477__),
    .I1(g690),
    .I0(__297__),
    .O(__754__)
  );
  LUT6 #(
    .INIT(64'hf888ffffffffffff)
  ) __1842__ (
    .I5(__754__),
    .I4(__751__),
    .I3(__298__),
    .I2(g723),
    .I1(__206__),
    .I0(g645),
    .O(__755__)
  );
  LUT6 #(
    .INIT(64'h8000000000000000)
  ) __1843__ (
    .I5(__480__),
    .I4(__47__),
    .I3(__413__),
    .I2(__460__),
    .I1(__182__),
    .I0(__157__),
    .O(__756__)
  );
  LUT4 #(
    .INIT(16'haa3c)
  ) __1844__ (
    .I3(__322__),
    .I2(__126__),
    .I1(__756__),
    .I0(__469__),
    .O(__757__)
  );
  LUT6 #(
    .INIT(64'h0000000000000040)
  ) __1845__ (
    .I5(__156__),
    .I4(__197__),
    .I3(__272__),
    .I2(__517__),
    .I1(__215__),
    .I0(__222__),
    .O(__758__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __1846__ (
    .I2(__758__),
    .I1(__73__),
    .I0(__493__),
    .O(__759__)
  );
  LUT2 #(
    .INIT(4'h7)
  ) __1847__ (
    .I1(__216__),
    .I0(__710__),
    .O(__760__)
  );
  LUT3 #(
    .INIT(8'hfd)
  ) __1848__ (
    .I2(__462__),
    .I1(__285__),
    .I0(__334__),
    .O(__761__)
  );
  LUT6 #(
    .INIT(64'h7fff800000000000)
  ) __1849__ (
    .I5(g781),
    .I4(__327__),
    .I3(__378__),
    .I2(__359__),
    .I1(__154__),
    .I0(__463__),
    .O(__762__)
  );
  LUT3 #(
    .INIT(8'h06)
  ) __1850__ (
    .I2(g43),
    .I1(__365__),
    .I0(__254__),
    .O(__763__)
  );
  LUT5 #(
    .INIT(32'h4f5f1000)
  ) __1851__ (
    .I4(__361__),
    .I3(__697__),
    .I2(__261__),
    .I1(__255__),
    .I0(__472__),
    .O(__764__)
  );
  LUT5 #(
    .INIT(32'hcaaaaaaa)
  ) __1852__ (
    .I4(__504__),
    .I3(__503__),
    .I2(__502__),
    .I1(__295__),
    .I0(__368__),
    .O(__765__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __1853__ (
    .I1(__188__),
    .I0(__300__),
    .O(__766__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __1854__ (
    .I1(__345__),
    .I0(__167__),
    .O(__767__)
  );
  LUT6 #(
    .INIT(64'h8000000000000000)
  ) __1855__ (
    .I5(__248__),
    .I4(__145__),
    .I3(__444__),
    .I2(__767__),
    .I1(__77__),
    .I0(__766__),
    .O(__768__)
  );
  LUT2 #(
    .INIT(4'h7)
  ) __1856__ (
    .I1(__768__),
    .I0(__117__),
    .O(__769__)
  );
  LUT5 #(
    .INIT(32'h00004000)
  ) __1857__ (
    .I4(__220__),
    .I3(__134__),
    .I2(__35__),
    .I1(__260__),
    .I0(__205__),
    .O(__770__)
  );
  LUT6 #(
    .INIT(64'h8000000000000000)
  ) __1858__ (
    .I5(__378__),
    .I4(__359__),
    .I3(__417__),
    .I2(__327__),
    .I1(__154__),
    .I0(__463__),
    .O(__771__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __1859__ (
    .I1(__49__),
    .I0(__771__),
    .O(__772__)
  );
  LUT5 #(
    .INIT(32'hcaaaaaaa)
  ) __1860__ (
    .I4(__504__),
    .I3(__503__),
    .I2(__536__),
    .I1(__290__),
    .I0(__56__),
    .O(__773__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __1861__ (
    .I3(__484__),
    .I2(__443__),
    .I1(__426__),
    .I0(__450__),
    .O(__774__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __1862__ (
    .I1(__378__),
    .I0(__359__),
    .O(__775__)
  );
  LUT6 #(
    .INIT(64'hec6c6c6cffffffff)
  ) __1863__ (
    .I5(g781),
    .I4(__417__),
    .I3(__327__),
    .I2(__154__),
    .I1(__463__),
    .I0(__775__),
    .O(__776__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __1864__ (
    .I1(g962),
    .I0(__28__),
    .O(__777__)
  );
  LUT6 #(
    .INIT(64'h0000000000000100)
  ) __1865__ (
    .I5(__316__),
    .I4(__24__),
    .I3(__777__),
    .I2(__55__),
    .I1(__399__),
    .I0(__198__),
    .O(__778__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __1866__ (
    .I2(g43),
    .I1(__778__),
    .I0(__461__),
    .O(__779__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __1867__ (
    .I1(__348__),
    .I0(__345__),
    .O(__780__)
  );
  LUT4 #(
    .INIT(16'hffd5)
  ) __1868__ (
    .I3(__146__),
    .I2(__48__),
    .I1(__62__),
    .I0(__46__),
    .O(__781__)
  );
  LUT3 #(
    .INIT(8'h78)
  ) __1869__ (
    .I2(__371__),
    .I1(__179__),
    .I0(g955),
    .O(__782__)
  );
  LUT6 #(
    .INIT(64'hbfffffffeaaaaaaa)
  ) __1870__ (
    .I5(__335__),
    .I4(__230__),
    .I3(__293__),
    .I2(__383__),
    .I1(__66__),
    .I0(__332__),
    .O(__783__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __1871__ (
    .I3(__419__),
    .I2(__82__),
    .I1(__470__),
    .I0(__274__),
    .O(__784__)
  );
  LUT6 #(
    .INIT(64'hf788778877887788)
  ) __1872__ (
    .I5(g786),
    .I4(__370__),
    .I3(__227__),
    .I2(__133__),
    .I1(__70__),
    .I0(__186__),
    .O(__785__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __1873__ (
    .I3(__74__),
    .I2(__489__),
    .I1(__294__),
    .I0(__479__),
    .O(__786__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __1874__ (
    .I2(__575__),
    .I1(__355__),
    .I0(__298__),
    .O(__787__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __1875__ (
    .I2(__665__),
    .I1(__409__),
    .I0(__193__),
    .O(__788__)
  );
  LUT3 #(
    .INIT(8'he2)
  ) __1876__ (
    .I2(g30),
    .I1(g32),
    .I0(g31),
    .O(__789__)
  );
  LUT5 #(
    .INIT(32'haaaa3fc0)
  ) __1877__ (
    .I4(__322__),
    .I3(__283__),
    .I2(__126__),
    .I1(__756__),
    .I0(__339__),
    .O(__790__)
  );
  LUT5 #(
    .INIT(32'h007f0080)
  ) __1878__ (
    .I4(__185__),
    .I3(__380__),
    .I2(__319__),
    .I1(__130__),
    .I0(__569__),
    .O(__791__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __1879__ (
    .I3(__419__),
    .I2(__82__),
    .I1(__176__),
    .I0(__490__),
    .O(__792__)
  );
  LUT2 #(
    .INIT(4'hb)
  ) __1880__ (
    .I1(__313__),
    .I0(__657__),
    .O(__793__)
  );
  LUT5 #(
    .INIT(32'h4f5f1000)
  ) __1881__ (
    .I4(__250__),
    .I3(__449__),
    .I2(__261__),
    .I1(__255__),
    .I0(__472__),
    .O(__794__)
  );
  LUT3 #(
    .INIT(8'ha3)
  ) __1882__ (
    .I2(__322__),
    .I1(__157__),
    .I0(__481__),
    .O(__795__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __1883__ (
    .I1(__70__),
    .I0(__186__),
    .O(__796__)
  );
  LUT4 #(
    .INIT(16'h0708)
  ) __1884__ (
    .I3(__45__),
    .I2(__380__),
    .I1(__267__),
    .I0(__177__),
    .O(__797__)
  );
  LUT3 #(
    .INIT(8'h10)
  ) __1885__ (
    .I2(__382__),
    .I1(__282__),
    .I0(__393__),
    .O(__798__)
  );
  LUT5 #(
    .INIT(32'h00003700)
  ) __1886__ (
    .I4(__140__),
    .I3(__778__),
    .I2(__340__),
    .I1(g43),
    .I0(__346__),
    .O(__799__)
  );
  LUT6 #(
    .INIT(64'h0000000000000040)
  ) __1887__ (
    .I5(__87__),
    .I4(g1),
    .I3(__779__),
    .I2(__799__),
    .I1(__398__),
    .I0(g1000),
    .O(__800__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __1888__ (
    .I1(__348__),
    .I0(__35__),
    .O(__801__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __1889__ (
    .I3(__484__),
    .I2(__443__),
    .I1(__76__),
    .I0(__452__),
    .O(__802__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __1890__ (
    .I1(__423__),
    .I0(__488__),
    .O(__803__)
  );
  LUT3 #(
    .INIT(8'h40)
  ) __1891__ (
    .I2(g43),
    .I1(g1),
    .I0(__778__),
    .O(__804__)
  );
  LUT5 #(
    .INIT(32'h7fff8000)
  ) __1892__ (
    .I4(__370__),
    .I3(__227__),
    .I2(__133__),
    .I1(__70__),
    .I0(__186__),
    .O(__805__)
  );
  LUT4 #(
    .INIT(16'h4000)
  ) __1893__ (
    .I3(__361__),
    .I2(__697__),
    .I1(__261__),
    .I0(__255__),
    .O(__806__)
  );
  LUT5 #(
    .INIT(32'h134c5f00)
  ) __1894__ (
    .I4(__187__),
    .I3(__232__),
    .I2(__261__),
    .I1(__806__),
    .I0(__472__),
    .O(__807__)
  );
  LUT4 #(
    .INIT(16'h0015)
  ) __1895__ (
    .I3(__258__),
    .I2(__18__),
    .I1(__153__),
    .I0(__468__),
    .O(__808__)
  );
  LUT4 #(
    .INIT(16'hbe00)
  ) __1896__ (
    .I3(__99__),
    .I2(__489__),
    .I1(g1198),
    .I0(__415__),
    .O(__809__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __1897__ (
    .I3(__334__),
    .I2(__462__),
    .I1(__39__),
    .I0(__79__),
    .O(__810__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __1898__ (
    .I1(__25__),
    .I0(__255__),
    .O(__811__)
  );
  LUT6 #(
    .INIT(64'h7fff800000000000)
  ) __1899__ (
    .I5(__694__),
    .I4(__129__),
    .I3(__244__),
    .I2(__811__),
    .I1(__280__),
    .I0(__688__),
    .O(__812__)
  );
  LUT5 #(
    .INIT(32'hcaaaaaaa)
  ) __1900__ (
    .I4(__520__),
    .I3(__512__),
    .I2(__215__),
    .I1(__216__),
    .I0(__89__),
    .O(__813__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __1901__ (
    .I1(__181__),
    .I0(__457__),
    .O(__814__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __1902__ (
    .I3(__419__),
    .I2(__82__),
    .I1(__356__),
    .I0(__410__),
    .O(__815__)
  );
  LUT4 #(
    .INIT(16'h8000)
  ) __1903__ (
    .I3(__445__),
    .I2(__283__),
    .I1(__126__),
    .I0(__756__),
    .O(__816__)
  );
  LUT6 #(
    .INIT(64'haaaaaaaa3fffc000)
  ) __1904__ (
    .I5(__322__),
    .I4(__487__),
    .I3(__90__),
    .I2(__816__),
    .I1(__390__),
    .I0(__85__),
    .O(__817__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __1905__ (
    .I3(__74__),
    .I2(__489__),
    .I1(__110__),
    .I0(__478__),
    .O(__818__)
  );
  LUT5 #(
    .INIT(32'h80000000)
  ) __1906__ (
    .I4(__90__),
    .I3(__445__),
    .I2(__283__),
    .I1(__126__),
    .I0(__756__),
    .O(__819__)
  );
  LUT4 #(
    .INIT(16'haa3c)
  ) __1907__ (
    .I3(__322__),
    .I2(__390__),
    .I1(__819__),
    .I0(__27__),
    .O(__820__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __1908__ (
    .I3(__484__),
    .I2(__443__),
    .I1(__376__),
    .I0(__455__),
    .O(__821__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __1909__ (
    .I3(__419__),
    .I2(__82__),
    .I1(__301__),
    .I0(__478__),
    .O(__822__)
  );
  LUT6 #(
    .INIT(64'h00000000ffff8000)
  ) __1910__ (
    .I5(__322__),
    .I4(__273__),
    .I3(__83__),
    .I2(__390__),
    .I1(__487__),
    .I0(__819__),
    .O(__823__)
  );
  LUT4 #(
    .INIT(16'hf7f8)
  ) __1911__ (
    .I3(__107__),
    .I2(__146__),
    .I1(__48__),
    .I0(__62__),
    .O(__824__)
  );
  LUT2 #(
    .INIT(4'hb)
  ) __1912__ (
    .I1(__313__),
    .I0(__641__),
    .O(__825__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __1913__ (
    .I1(__391__),
    .I0(__434__),
    .O(__826__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __1914__ (
    .I1(__188__),
    .I0(__300__),
    .O(__827__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __1915__ (
    .I1(__167__),
    .I0(__145__),
    .O(__828__)
  );
  LUT6 #(
    .INIT(64'hfffeffffffffffff)
  ) __1916__ (
    .I5(__828__),
    .I4(__827__),
    .I3(__345__),
    .I2(__248__),
    .I1(__444__),
    .I0(__77__),
    .O(__829__)
  );
  LUT4 #(
    .INIT(16'h3700)
  ) __1917__ (
    .I3(__391__),
    .I2(__118__),
    .I1(__768__),
    .I0(__117__),
    .O(__830__)
  );
  LUT6 #(
    .INIT(64'h0000000000004000)
  ) __1918__ (
    .I5(__87__),
    .I4(__779__),
    .I3(g43),
    .I2(__799__),
    .I1(__19__),
    .I0(g1000),
    .O(__831__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __1919__ (
    .I3(__484__),
    .I2(__443__),
    .I1(__125__),
    .I0(__256__),
    .O(__832__)
  );
  LUT4 #(
    .INIT(16'h000b)
  ) __1920__ (
    .I3(g43),
    .I2(__254__),
    .I1(__492__),
    .I0(__365__),
    .O(__833__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __1921__ (
    .I2(__665__),
    .I1(__451__),
    .I0(__351__),
    .O(__834__)
  );
  LUT6 #(
    .INIT(64'hfffffffffffffffe)
  ) __1922__ (
    .I5(__472__),
    .I4(__320__),
    .I3(__437__),
    .I2(__160__),
    .I1(__235__),
    .I0(__65__),
    .O(__835__)
  );
  LUT2 #(
    .INIT(4'h7)
  ) __1923__ (
    .I1(__18__),
    .I0(__264__),
    .O(__836__)
  );
  LUT6 #(
    .INIT(64'hda5a5a5affffffff)
  ) __1924__ (
    .I5(g781),
    .I4(__417__),
    .I3(__327__),
    .I2(__154__),
    .I1(__463__),
    .I0(__775__),
    .O(__837__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __1925__ (
    .I2(__719__),
    .I1(__285__),
    .I0(__297__),
    .O(__838__)
  );
  LUT6 #(
    .INIT(64'h0000000000000001)
  ) __1926__ (
    .I5(__208__),
    .I4(__384__),
    .I3(__189__),
    .I2(__199__),
    .I1(__34__),
    .I0(__64__),
    .O(__839__)
  );
  LUT3 #(
    .INIT(8'h01)
  ) __1927__ (
    .I2(__317__),
    .I1(__171__),
    .I0(__257__),
    .O(__840__)
  );
  LUT6 #(
    .INIT(64'h0000000000000040)
  ) __1928__ (
    .I5(__219__),
    .I4(__150__),
    .I3(__287__),
    .I2(__840__),
    .I1(__839__),
    .I0(__183__),
    .O(__841__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __1929__ (
    .I2(__541__),
    .I1(__58__),
    .I0(__442__),
    .O(__842__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __1930__ (
    .I2(__527__),
    .I1(__21__),
    .I0(__367__),
    .O(__843__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __1931__ (
    .I3(__74__),
    .I2(__489__),
    .I1(__358__),
    .I0(__490__),
    .O(__844__)
  );
  LUT3 #(
    .INIT(8'h04)
  ) __1932__ (
    .I2(__177__),
    .I1(__381__),
    .I0(__119__),
    .O(__845__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __1933__ (
    .I2(g43),
    .I1(__778__),
    .I0(__346__),
    .O(__846__)
  );
  LUT4 #(
    .INIT(16'ha3af)
  ) __1934__ (
    .I3(__18__),
    .I2(__381__),
    .I1(__264__),
    .I0(__226__),
    .O(__847__)
  );
  LUT6 #(
    .INIT(64'hf8f078f078f078f0)
  ) __1935__ (
    .I5(g786),
    .I4(__370__),
    .I3(__227__),
    .I2(__133__),
    .I1(__70__),
    .I0(__186__),
    .O(__848__)
  );
  LUT5 #(
    .INIT(32'h3f7f3333)
  ) __1936__ (
    .I4(__391__),
    .I3(__118__),
    .I2(__768__),
    .I1(__16__),
    .I0(__117__),
    .O(__849__)
  );
  LUT2 #(
    .INIT(4'h7)
  ) __1937__ (
    .I1(__312__),
    .I0(__710__),
    .O(__850__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __1938__ (
    .I3(__386__),
    .I2(__147__),
    .I1(__353__),
    .I0(__256__),
    .O(__851__)
  );
  LUT6 #(
    .INIT(64'haaaaaaaa3fffc000)
  ) __1939__ (
    .I5(__322__),
    .I4(__445__),
    .I3(__283__),
    .I2(__126__),
    .I1(__756__),
    .I0(__249__),
    .O(__852__)
  );
  LUT4 #(
    .INIT(16'hb400)
  ) __1940__ (
    .I3(__694__),
    .I2(__29__),
    .I1(__307__),
    .I0(__255__),
    .O(__853__)
  );
  LUT5 #(
    .INIT(32'h00000001)
  ) __1941__ (
    .I4(__213__),
    .I3(__200__),
    .I2(__447__),
    .I1(__23__),
    .I0(__151__),
    .O(__854__)
  );
  LUT6 #(
    .INIT(64'h8000000000000000)
  ) __1942__ (
    .I5(__52__),
    .I4(__213__),
    .I3(__200__),
    .I2(__447__),
    .I1(__23__),
    .I0(__151__),
    .O(__855__)
  );
  LUT6 #(
    .INIT(64'hf000000000000044)
  ) __1943__ (
    .I5(__344__),
    .I4(__286__),
    .I3(__135__),
    .I2(__855__),
    .I1(__854__),
    .I0(__52__),
    .O(__856__)
  );
  LUT5 #(
    .INIT(32'h00000001)
  ) __1944__ (
    .I4(__42__),
    .I3(__242__),
    .I2(__144__),
    .I1(__49__),
    .I0(__856__),
    .O(__857__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __1945__ (
    .I3(__484__),
    .I2(__443__),
    .I1(__421__),
    .I0(__485__),
    .O(__858__)
  );
  LUT5 #(
    .INIT(32'h7f800000)
  ) __1946__ (
    .I4(__391__),
    .I3(__420__),
    .I2(__124__),
    .I1(__276__),
    .I0(__434__),
    .O(__859__)
  );
  LUT4 #(
    .INIT(16'hbe00)
  ) __1947__ (
    .I3(__99__),
    .I2(__82__),
    .I1(g1202),
    .I0(__61__),
    .O(__860__)
  );
  LUT4 #(
    .INIT(16'h8000)
  ) __1948__ (
    .I3(__378__),
    .I2(__359__),
    .I1(__154__),
    .I0(__463__),
    .O(__861__)
  );
  LUT4 #(
    .INIT(16'h7800)
  ) __1949__ (
    .I3(g781),
    .I2(__417__),
    .I1(__327__),
    .I0(__861__),
    .O(__862__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __1950__ (
    .I2(__575__),
    .I1(__216__),
    .I0(__246__),
    .O(__863__)
  );
  LUT5 #(
    .INIT(32'h80000000)
  ) __1951__ (
    .I4(__14__),
    .I3(__240__),
    .I2(__210__),
    .I1(__225__),
    .I0(__578__),
    .O(__864__)
  );
  LUT5 #(
    .INIT(32'hfffffffe)
  ) __1952__ (
    .I4(__864__),
    .I3(__251__),
    .I2(__221__),
    .I1(__163__),
    .I0(__331__),
    .O(__865__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __1953__ (
    .I3(__74__),
    .I2(__489__),
    .I1(__385__),
    .I0(__364__),
    .O(__866__)
  );
  LUT5 #(
    .INIT(32'h5a5a335a)
  ) __1954__ (
    .I4(__87__),
    .I3(__431__),
    .I2(__693__),
    .I1(__475__),
    .I0(__212__),
    .O(__867__)
  );
  LUT3 #(
    .INIT(8'h40)
  ) __1955__ (
    .I2(g43),
    .I1(__340__),
    .I0(__140__),
    .O(__868__)
  );
  LUT4 #(
    .INIT(16'h4000)
  ) __1956__ (
    .I3(__250__),
    .I2(__449__),
    .I1(__261__),
    .I0(__255__),
    .O(__869__)
  );
  LUT5 #(
    .INIT(32'h134c5f00)
  ) __1957__ (
    .I4(__75__),
    .I3(__245__),
    .I2(__261__),
    .I1(__869__),
    .I0(__472__),
    .O(__870__)
  );
  LUT6 #(
    .INIT(64'hbfff400000000000)
  ) __1958__ (
    .I5(__694__),
    .I4(__374__),
    .I3(__115__),
    .I2(__29__),
    .I1(__307__),
    .I0(__255__),
    .O(__871__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __1959__ (
    .I2(__541__),
    .I1(__385__),
    .I0(__459__),
    .O(__872__)
  );
  LUT5 #(
    .INIT(32'hcaaaaaaa)
  ) __1960__ (
    .I4(__504__),
    .I3(__503__),
    .I2(__536__),
    .I1(__426__),
    .I0(__408__),
    .O(__873__)
  );
  LUT6 #(
    .INIT(64'h8000000000000000)
  ) __1961__ (
    .I5(__357__),
    .I4(__232__),
    .I3(__361__),
    .I2(__311__),
    .I1(__187__),
    .I0(__721__),
    .O(__874__)
  );
  LUT6 #(
    .INIT(64'h135f4c005f5f0000)
  ) __1962__ (
    .I5(__59__),
    .I4(__17__),
    .I3(__98__),
    .I2(__261__),
    .I1(__874__),
    .I0(__472__),
    .O(__875__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __1963__ (
    .I2(__527__),
    .I1(__176__),
    .I0(__458__),
    .O(__876__)
  );
  LUT6 #(
    .INIT(64'hbfffffffeaaaaaaa)
  ) __1964__ (
    .I5(__260__),
    .I4(__134__),
    .I3(__35__),
    .I2(__220__),
    .I1(__205__),
    .I0(__258__),
    .O(__877__)
  );
  LUT5 #(
    .INIT(32'h143c3c3c)
  ) __1965__ (
    .I4(__179__),
    .I3(g955),
    .I2(__334__),
    .I1(__462__),
    .I0(__371__),
    .O(__878__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __1966__ (
    .I3(__419__),
    .I2(__82__),
    .I1(__427__),
    .I0(__364__),
    .O(__879__)
  );
  LUT4 #(
    .INIT(16'h001c)
  ) __1967__ (
    .I3(__146__),
    .I2(__48__),
    .I1(__46__),
    .I0(__62__),
    .O(__880__)
  );
  LUT4 #(
    .INIT(16'h4000)
  ) __1968__ (
    .I3(g43),
    .I2(__778__),
    .I1(__346__),
    .I0(__140__),
    .O(__881__)
  );
  LUT3 #(
    .INIT(8'h60)
  ) __1969__ (
    .I2(__391__),
    .I1(__404__),
    .I0(__707__),
    .O(__882__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __1970__ (
    .I3(__484__),
    .I2(__443__),
    .I1(__290__),
    .I0(__253__),
    .O(__883__)
  );
  LUT5 #(
    .INIT(32'hff7fff80)
  ) __1971__ (
    .I4(__372__),
    .I3(__332__),
    .I2(__33__),
    .I1(__507__),
    .I0(__66__),
    .O(__884__)
  );
  LUT6 #(
    .INIT(64'h00007fff00008000)
  ) __1972__ (
    .I5(__190__),
    .I4(__380__),
    .I3(__341__),
    .I2(__45__),
    .I1(__267__),
    .I0(__177__),
    .O(__885__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __1973__ (
    .I3(__484__),
    .I2(__443__),
    .I1(__116__),
    .I0(__109__),
    .O(__886__)
  );
  LUT2 #(
    .INIT(4'h7)
  ) __1974__ (
    .I1(__216__),
    .I0(__510__),
    .O(__887__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __1975__ (
    .I1(__182__),
    .I0(__157__),
    .O(__888__)
  );
  LUT6 #(
    .INIT(64'haaaaaaaa3fffc000)
  ) __1976__ (
    .I5(__322__),
    .I4(__480__),
    .I3(__413__),
    .I2(__460__),
    .I1(__888__),
    .I0(__95__),
    .O(__889__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __1977__ (
    .I3(__484__),
    .I2(__443__),
    .I1(__409__),
    .I0(__277__),
    .O(__890__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __1978__ (
    .I3(__74__),
    .I2(__489__),
    .I1(__58__),
    .I0(__494__),
    .O(__891__)
  );
  LUT2 #(
    .INIT(4'h7)
  ) __1979__ (
    .I1(__79__),
    .I0(__510__),
    .O(__892__)
  );
  LUT4 #(
    .INIT(16'hbe00)
  ) __1980__ (
    .I3(__99__),
    .I2(__147__),
    .I1(g1194),
    .I0(__446__),
    .O(__893__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __1981__ (
    .I2(__541__),
    .I1(__486__),
    .I0(__392__),
    .O(__894__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __1982__ (
    .I2(__460__),
    .I1(__182__),
    .I0(__157__),
    .O(__895__)
  );
  LUT6 #(
    .INIT(64'haaaaaaaa3fffc000)
  ) __1983__ (
    .I5(__322__),
    .I4(__47__),
    .I3(__480__),
    .I2(__413__),
    .I1(__895__),
    .I0(__201__),
    .O(__896__)
  );
  LUT6 #(
    .INIT(64'h4f5f5f5f10000000)
  ) __1984__ (
    .I5(__75__),
    .I4(__250__),
    .I3(__449__),
    .I2(__261__),
    .I1(__255__),
    .I0(__472__),
    .O(__897__)
  );
  LUT5 #(
    .INIT(32'hbf400000)
  ) __1985__ (
    .I4(__694__),
    .I3(__115__),
    .I2(__29__),
    .I1(__307__),
    .I0(__255__),
    .O(__898__)
  );
  LUT4 #(
    .INIT(16'hba00)
  ) __1986__ (
    .I3(g43),
    .I2(__93__),
    .I1(__425__),
    .I0(__87__),
    .O(__899__)
  );
  LUT5 #(
    .INIT(32'hf0fe0000)
  ) __1987__ (
    .I4(__899__),
    .I3(__476__),
    .I2(__425__),
    .I1(__429__),
    .I0(__121__),
    .O(__900__)
  );
  LUT4 #(
    .INIT(16'hbe00)
  ) __1988__ (
    .I3(__99__),
    .I2(__443__),
    .I1(g1206),
    .I0(__473__),
    .O(__901__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __1989__ (
    .I2(__665__),
    .I1(__262__),
    .I0(__414__),
    .O(__902__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __1990__ (
    .I1(__233__),
    .I0(__188__),
    .O(__903__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __1991__ (
    .I3(__419__),
    .I2(__82__),
    .I1(__394__),
    .I0(__479__),
    .O(__904__)
  );
  LUT6 #(
    .INIT(64'haaaaaaaa3fffc000)
  ) __1992__ (
    .I5(__322__),
    .I4(__413__),
    .I3(__460__),
    .I2(__182__),
    .I1(__157__),
    .I0(__439__),
    .O(__905__)
  );
  LUT6 #(
    .INIT(64'hbfffffffeaaaaaaa)
  ) __1993__ (
    .I5(__225__),
    .I4(__14__),
    .I3(__240__),
    .I2(__578__),
    .I1(__66__),
    .I0(__332__),
    .O(__906__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __1994__ (
    .I2(__694__),
    .I1(__255__),
    .I0(__307__),
    .O(__907__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __1995__ (
    .I3(__334__),
    .I2(__462__),
    .I1(__388__),
    .I0(__387__),
    .O(__908__)
  );
  LUT5 #(
    .INIT(32'h80000000)
  ) __1996__ (
    .I4(__115__),
    .I3(__374__),
    .I2(__29__),
    .I1(__307__),
    .I0(__412__),
    .O(__909__)
  );
  LUT4 #(
    .INIT(16'hb400)
  ) __1997__ (
    .I3(__694__),
    .I2(__464__),
    .I1(__909__),
    .I0(__255__),
    .O(__910__)
  );
  LUT5 #(
    .INIT(32'hcaaaaaaa)
  ) __1998__ (
    .I4(__504__),
    .I3(__517__),
    .I2(__215__),
    .I1(__387__),
    .I0(__416__),
    .O(__911__)
  );
  LUT2 #(
    .INIT(4'h7)
  ) __1999__ (
    .I1(__768__),
    .I0(__88__),
    .O(__912__)
  );
  LUT2 #(
    .INIT(4'h7)
  ) __2000__ (
    .I1(__355__),
    .I0(__510__),
    .O(__913__)
  );
  LUT5 #(
    .INIT(32'h30020000)
  ) __2001__ (
    .I4(__899__),
    .I3(__476__),
    .I2(__121__),
    .I1(__425__),
    .I0(__429__),
    .O(__914__)
  );
  LUT4 #(
    .INIT(16'h0100)
  ) __2002__ (
    .I3(__854__),
    .I2(__344__),
    .I1(__286__),
    .I0(__135__),
    .O(__915__)
  );
  LUT5 #(
    .INIT(32'h0000000e)
  ) __2003__ (
    .I4(__42__),
    .I3(__704__),
    .I2(__144__),
    .I1(__453__),
    .I0(__915__),
    .O(__916__)
  );
  LUT6 #(
    .INIT(64'h0f0e0f0f0f0f000f)
  ) __2004__ (
    .I5(__42__),
    .I4(__144__),
    .I3(__242__),
    .I2(__916__),
    .I1(__453__),
    .I0(__424__),
    .O(__917__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __2005__ (
    .I1(__192__),
    .I0(__917__),
    .O(__918__)
  );
  LUT6 #(
    .INIT(64'hf3faf0f0f0f0f0f0)
  ) __2006__ (
    .I5(__42__),
    .I4(__242__),
    .I3(__144__),
    .I2(__918__),
    .I1(__704__),
    .I0(__181__),
    .O(__919__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __2007__ (
    .I2(__319__),
    .I1(__185__),
    .I0(__130__),
    .O(__920__)
  );
  LUT6 #(
    .INIT(64'h8000000000000000)
  ) __2008__ (
    .I5(__279__),
    .I4(__920__),
    .I3(__190__),
    .I2(__341__),
    .I1(__45__),
    .I0(__267__),
    .O(__921__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __2009__ (
    .I3(__334__),
    .I2(__462__),
    .I1(__483__),
    .I0(__73__),
    .O(__922__)
  );
  LUT5 #(
    .INIT(32'hcaaaaaaa)
  ) __2010__ (
    .I4(__504__),
    .I3(__503__),
    .I2(__536__),
    .I1(__50__),
    .I0(__231__),
    .O(__923__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __2011__ (
    .I2(g43),
    .I1(g1),
    .I0(g10),
    .O(__924__)
  );
  LUT4 #(
    .INIT(16'h0040)
  ) __2012__ (
    .I3(g1),
    .I2(__252__),
    .I1(__398__),
    .I0(g1000),
    .O(__925__)
  );
  LUT6 #(
    .INIT(64'h000000000000efff)
  ) __2013__ (
    .I5(__846__),
    .I4(__925__),
    .I3(__178__),
    .I2(__924__),
    .I1(g1008),
    .I0(g1016),
    .O(__926__)
  );
  LUT3 #(
    .INIT(8'hbf)
  ) __2014__ (
    .I2(g43),
    .I1(__93__),
    .I0(__425__),
    .O(__927__)
  );
  LUT6 #(
    .INIT(64'h0000000010ffffff)
  ) __2015__ (
    .I5(__779__),
    .I4(__927__),
    .I3(__926__),
    .I2(__476__),
    .I1(__429__),
    .I0(__121__),
    .O(__928__)
  );
  LUT5 #(
    .INIT(32'hcaaaaaaa)
  ) __2016__ (
    .I4(__504__),
    .I3(__503__),
    .I2(__536__),
    .I1(__97__),
    .I0(__84__),
    .O(__929__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __2017__ (
    .I3(__386__),
    .I2(__147__),
    .I1(__482__),
    .I0(__191__),
    .O(__930__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __2018__ (
    .I2(__719__),
    .I1(__79__),
    .I0(__168__),
    .O(__931__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __2019__ (
    .I1(__564__),
    .I0(__657__),
    .O(__932__)
  );
  LUT6 #(
    .INIT(64'h3cc3aaaaffffffff)
  ) __2020__ (
    .I5(__313__),
    .I4(g44),
    .I3(__675__),
    .I2(__932__),
    .I1(__642__),
    .I0(__678__),
    .O(__933__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __2021__ (
    .I1(__778__),
    .I0(g1),
    .O(__934__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __2022__ (
    .I1(g1),
    .I0(__778__),
    .O(__935__)
  );
  LUT2 #(
    .INIT(4'h7)
  ) __2023__ (
    .I1(__405__),
    .I0(__710__),
    .O(__936__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __2024__ (
    .I3(__484__),
    .I2(__443__),
    .I1(__271__),
    .I0(__410__),
    .O(__937__)
  );
  LUT5 #(
    .INIT(32'h007f8080)
  ) __2025__ (
    .I4(__91__),
    .I3(__411__),
    .I2(__261__),
    .I1(__142__),
    .I0(__437__),
    .O(__938__)
  );
  LUT2 #(
    .INIT(4'hb)
  ) __2026__ (
    .I1(__313__),
    .I0(__618__),
    .O(__939__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __2027__ (
    .I2(__719__),
    .I1(__216__),
    .I0(__237__),
    .O(__940__)
  );
  LUT4 #(
    .INIT(16'hd0f0)
  ) __2028__ (
    .I3(g43),
    .I2(__87__),
    .I1(__140__),
    .I0(__340__),
    .O(__941__)
  );
  LUT5 #(
    .INIT(32'h51f3ffff)
  ) __2029__ (
    .I4(g43),
    .I3(__778__),
    .I2(__140__),
    .I1(__340__),
    .I0(__346__),
    .O(__942__)
  );
  LUT5 #(
    .INIT(32'h0fbf0f0f)
  ) __2030__ (
    .I4(__942__),
    .I3(__148__),
    .I2(g1),
    .I1(__927__),
    .I0(g10),
    .O(__943__)
  );
  LUT4 #(
    .INIT(16'hffd5)
  ) __2031__ (
    .I3(__177__),
    .I2(__382__),
    .I1(__282__),
    .I0(__393__),
    .O(__944__)
  );
  LUT4 #(
    .INIT(16'hb400)
  ) __2032__ (
    .I3(__694__),
    .I2(__280__),
    .I1(__688__),
    .I0(__255__),
    .O(__945__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __2033__ (
    .I3(__386__),
    .I2(__147__),
    .I1(__60__),
    .I0(__274__),
    .O(__946__)
  );
  LUT6 #(
    .INIT(64'h000080007fff8000)
  ) __2034__ (
    .I5(__261__),
    .I4(__472__),
    .I3(__59__),
    .I2(__98__),
    .I1(__874__),
    .I0(__17__),
    .O(__947__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __2035__ (
    .I3(__484__),
    .I2(__443__),
    .I1(__379__),
    .I0(__149__),
    .O(__948__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __2036__ (
    .I1(g781),
    .I0(__378__),
    .O(__949__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __2037__ (
    .I2(__527__),
    .I1(__292__),
    .I0(__329__),
    .O(__950__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __2038__ (
    .I3(__484__),
    .I2(__443__),
    .I1(__214__),
    .I0(__478__),
    .O(__951__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __2039__ (
    .I3(__484__),
    .I2(__443__),
    .I1(__50__),
    .I0(__438__),
    .O(__952__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __2040__ (
    .I1(__197__),
    .I0(__145__),
    .O(__953__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __2041__ (
    .I2(__35__),
    .I1(__220__),
    .I0(__205__),
    .O(__954__)
  );
  LUT5 #(
    .INIT(32'hff7fff80)
  ) __2042__ (
    .I4(__444__),
    .I3(__258__),
    .I2(__134__),
    .I1(__260__),
    .I0(__954__),
    .O(__955__)
  );
  LUT5 #(
    .INIT(32'h7f800000)
  ) __2043__ (
    .I4(__391__),
    .I3(__138__),
    .I2(__440__),
    .I1(__404__),
    .I0(__707__),
    .O(__956__)
  );
  LUT4 #(
    .INIT(16'h4000)
  ) __2044__ (
    .I3(__42__),
    .I2(__144__),
    .I1(__457__),
    .I0(__242__),
    .O(__957__)
  );
  LUT2 #(
    .INIT(4'h7)
  ) __2045__ (
    .I1(__118__),
    .I0(__768__),
    .O(__958__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __2046__ (
    .I2(__719__),
    .I1(__73__),
    .I0(__94__),
    .O(__959__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __2047__ (
    .I3(__386__),
    .I2(__147__),
    .I1(__375__),
    .I0(__455__),
    .O(__960__)
  );
  LUT3 #(
    .INIT(8'h60)
  ) __2048__ (
    .I2(g781),
    .I1(__378__),
    .I0(__359__),
    .O(__961__)
  );
  LUT4 #(
    .INIT(16'h8000)
  ) __2049__ (
    .I3(__124__),
    .I2(__420__),
    .I1(__276__),
    .I0(__434__),
    .O(__962__)
  );
  LUT4 #(
    .INIT(16'h7800)
  ) __2050__ (
    .I3(__391__),
    .I2(__202__),
    .I1(__318__),
    .I0(__962__),
    .O(__963__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __2051__ (
    .I1(__22__),
    .I0(__343__),
    .O(__964__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __2052__ (
    .I3(__484__),
    .I2(__443__),
    .I1(__165__),
    .I0(__364__),
    .O(__965__)
  );
  LUT2 #(
    .INIT(4'h7)
  ) __2053__ (
    .I1(__73__),
    .I0(__510__),
    .O(__966__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __2054__ (
    .I2(__527__),
    .I1(__112__),
    .I0(__333__),
    .O(__967__)
  );
  LUT5 #(
    .INIT(32'hf0fbf0f0)
  ) __2055__ (
    .I4(__533__),
    .I3(__664__),
    .I2(__674__),
    .I1(__662__),
    .I0(__530__),
    .O(__968__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __2056__ (
    .I2(__758__),
    .I1(__312__),
    .I0(__304__),
    .O(__969__)
  );
  LUT4 #(
    .INIT(16'h0015)
  ) __2057__ (
    .I3(__258__),
    .I2(__264__),
    .I1(__169__),
    .I0(__146__),
    .O(__970__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __2058__ (
    .I2(__575__),
    .I1(__312__),
    .I0(__299__),
    .O(__971__)
  );
  LUT6 #(
    .INIT(64'h0000000000004000)
  ) __2059__ (
    .I5(__87__),
    .I4(__19__),
    .I3(__799__),
    .I2(__81__),
    .I1(__924__),
    .I0(__779__),
    .O(__972__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __2060__ (
    .I3(__419__),
    .I2(__82__),
    .I1(__309__),
    .I0(__253__),
    .O(__973__)
  );
  LUT6 #(
    .INIT(64'h7fffffff80000000)
  ) __2061__ (
    .I5(g786),
    .I4(__370__),
    .I3(__227__),
    .I2(__133__),
    .I1(__70__),
    .I0(__186__),
    .O(__974__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __2062__ (
    .I3(__419__),
    .I2(__82__),
    .I1(__21__),
    .I0(__494__),
    .O(__975__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __2063__ (
    .I1(__578__),
    .I0(__66__),
    .O(__976__)
  );
  LUT6 #(
    .INIT(64'h00007fff00008000)
  ) __2064__ (
    .I5(__210__),
    .I4(__332__),
    .I3(__14__),
    .I2(__240__),
    .I1(__225__),
    .I0(__976__),
    .O(__977__)
  );
  LUT4 #(
    .INIT(16'heffe)
  ) __2065__ (
    .I3(__319__),
    .I2(__569__),
    .I1(__380__),
    .I0(__921__),
    .O(__978__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __2066__ (
    .I1(__92__),
    .I0(g929),
    .O(__979__)
  );
  LUT5 #(
    .INIT(32'hfcff5455)
  ) __2067__ (
    .I4(__87__),
    .I3(__492__),
    .I2(__365__),
    .I1(__254__),
    .I0(__926__),
    .O(__980__)
  );
  LUT3 #(
    .INIT(8'h4f)
  ) __2068__ (
    .I2(g1),
    .I1(__942__),
    .I0(__148__),
    .O(__981__)
  );
  LUT6 #(
    .INIT(64'hbfff400000000000)
  ) __2069__ (
    .I5(__694__),
    .I4(__244__),
    .I3(__280__),
    .I2(__464__),
    .I1(__909__),
    .I0(__255__),
    .O(__982__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __2070__ (
    .I3(__419__),
    .I2(__82__),
    .I1(__67__),
    .I0(__485__),
    .O(__983__)
  );
  LUT6 #(
    .INIT(64'hf0ffffaaff33ffff)
  ) __2071__ (
    .I5(__42__),
    .I4(__242__),
    .I3(__144__),
    .I2(__704__),
    .I1(__453__),
    .I0(__457__),
    .O(__984__)
  );
  LUT5 #(
    .INIT(32'h33733333)
  ) __2072__ (
    .I4(__42__),
    .I3(__242__),
    .I2(__144__),
    .I1(__984__),
    .I0(__424__),
    .O(__985__)
  );
  LUT5 #(
    .INIT(32'hcaaaaaaa)
  ) __2073__ (
    .I4(__504__),
    .I3(__503__),
    .I2(__540__),
    .I1(__358__),
    .I0(__43__),
    .O(__986__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __2074__ (
    .I2(__527__),
    .I1(__309__),
    .I0(__152__),
    .O(__987__)
  );
  LUT4 #(
    .INIT(16'hf0ee)
  ) __2075__ (
    .I3(__583__),
    .I2(__387__),
    .I1(__453__),
    .I0(__128__),
    .O(__988__)
  );
  LUT3 #(
    .INIT(8'h40)
  ) __2076__ (
    .I2(__282__),
    .I1(__393__),
    .I0(__382__),
    .O(__989__)
  );
  LUT4 #(
    .INIT(16'h0230)
  ) __2077__ (
    .I3(__382__),
    .I2(__282__),
    .I1(__177__),
    .I0(__393__),
    .O(__990__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __2078__ (
    .I1(__281__),
    .I0(__87__),
    .O(__991__)
  );
  LUT4 #(
    .INIT(16'h152a)
  ) __2079__ (
    .I3(__98__),
    .I2(__261__),
    .I1(__472__),
    .I0(__874__),
    .O(__992__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __2080__ (
    .I2(__665__),
    .I1(__96__),
    .I0(__41__),
    .O(__993__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __2081__ (
    .I3(__74__),
    .I2(__489__),
    .I1(__114__),
    .I0(__485__),
    .O(__994__)
  );
  LUT2 #(
    .INIT(4'hb)
  ) __2082__ (
    .I1(__220__),
    .I0(__258__),
    .O(__995__)
  );
  LUT6 #(
    .INIT(64'hbfff400000000000)
  ) __2083__ (
    .I5(__694__),
    .I4(__25__),
    .I3(__244__),
    .I2(__280__),
    .I1(__688__),
    .I0(__255__),
    .O(__996__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __2084__ (
    .I3(__334__),
    .I2(__462__),
    .I1(__373__),
    .I0(__405__),
    .O(__997__)
  );
  LUT3 #(
    .INIT(8'h78)
  ) __2085__ (
    .I2(__40__),
    .I1(__92__),
    .I0(g929),
    .O(__998__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __2086__ (
    .I1(__173__),
    .I0(__205__),
    .O(__999__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __2087__ (
    .I1(__173__),
    .I0(__167__),
    .O(__1000__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __2088__ (
    .I2(__758__),
    .I1(__285__),
    .I0(__338__),
    .O(__1001__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __2089__ (
    .I2(__719__),
    .I1(__387__),
    .I0(__158__),
    .O(__1002__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __2090__ (
    .I2(__758__),
    .I1(__216__),
    .I0(__19__),
    .O(__1003__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __2091__ (
    .I3(__74__),
    .I2(__489__),
    .I1(__100__),
    .I0(__274__),
    .O(__1004__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __2092__ (
    .I1(__454__),
    .I0(__300__),
    .O(__1005__)
  );
  LUT4 #(
    .INIT(16'h0060)
  ) __2093__ (
    .I3(__258__),
    .I2(__103__),
    .I1(__300__),
    .I0(__705__),
    .O(__1006__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __2094__ (
    .I2(__669__),
    .I1(__403__),
    .I0(__349__),
    .O(__1007__)
  );
  LUT2 #(
    .INIT(4'hb)
  ) __2095__ (
    .I1(__51__),
    .I0(__36__),
    .O(__1008__)
  );
  LUT5 #(
    .INIT(32'hff00f8f8)
  ) __2096__ (
    .I4(__726__),
    .I3(__312__),
    .I2(__170__),
    .I1(__296__),
    .I0(__725__),
    .O(__1009__)
  );
  LUT5 #(
    .INIT(32'h134c5f00)
  ) __2097__ (
    .I4(__98__),
    .I3(__59__),
    .I2(__261__),
    .I1(__874__),
    .I0(__472__),
    .O(__1010__)
  );
  LUT6 #(
    .INIT(64'haaaaaaaa3fffc000)
  ) __2098__ (
    .I5(__322__),
    .I4(__83__),
    .I3(__390__),
    .I2(__487__),
    .I1(__819__),
    .I0(__113__),
    .O(__1011__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __2099__ (
    .I2(__527__),
    .I1(__427__),
    .I0(__396__),
    .O(__1012__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __2100__ (
    .I3(__74__),
    .I2(__489__),
    .I1(__306__),
    .I0(__109__),
    .O(__1013__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __2101__ (
    .I3(__386__),
    .I2(__147__),
    .I1(__102__),
    .I0(__410__),
    .O(__1014__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __2102__ (
    .I1(__272__),
    .I0(__248__),
    .O(__1015__)
  );
  LUT3 #(
    .INIT(8'hb0)
  ) __2103__ (
    .I2(__207__),
    .I1(__462__),
    .I0(__334__),
    .O(__1016__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __2104__ (
    .I2(__42__),
    .I1(__242__),
    .I0(__144__),
    .O(__1017__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __2105__ (
    .I3(__484__),
    .I2(__443__),
    .I1(__96__),
    .I0(__288__),
    .O(__1018__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __2106__ (
    .I2(__527__),
    .I1(__127__),
    .I0(__184__),
    .O(__1019__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __2107__ (
    .I3(__386__),
    .I2(__147__),
    .I1(__72__),
    .I0(__253__),
    .O(__1020__)
  );
  LUT2 #(
    .INIT(4'he)
  ) __2108__ (
    .I1(__432__),
    .I0(__263__),
    .O(__1021__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __2109__ (
    .I3(__484__),
    .I2(__443__),
    .I1(__241__),
    .I0(__274__),
    .O(__1022__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __2110__ (
    .I3(__386__),
    .I2(__147__),
    .I1(__433__),
    .I0(__478__),
    .O(__1023__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __2111__ (
    .I3(__74__),
    .I2(__489__),
    .I1(__456__),
    .I0(__455__),
    .O(__1024__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __2112__ (
    .I1(__454__),
    .I0(__134__),
    .O(__1025__)
  );
  LUT3 #(
    .INIT(8'hfe)
  ) __2113__ (
    .I2(__258__),
    .I1(__146__),
    .I0(__264__),
    .O(__1026__)
  );
  LUT4 #(
    .INIT(16'hb400)
  ) __2114__ (
    .I3(__694__),
    .I2(__412__),
    .I1(__692__),
    .I0(__255__),
    .O(__1027__)
  );
  LUT5 #(
    .INIT(32'hff7fff80)
  ) __2115__ (
    .I4(__240__),
    .I3(__332__),
    .I2(__14__),
    .I1(__578__),
    .I0(__66__),
    .O(__1028__)
  );
  LUT3 #(
    .INIT(8'hf1)
  ) __2116__ (
    .I2(__177__),
    .I1(__119__),
    .I0(__381__),
    .O(__1029__)
  );
  LUT4 #(
    .INIT(16'h00ca)
  ) __2117__ (
    .I3(__466__),
    .I2(__758__),
    .I1(__405__),
    .I0(__281__),
    .O(__1030__)
  );
  LUT4 #(
    .INIT(16'h0708)
  ) __2118__ (
    .I3(__492__),
    .I2(g43),
    .I1(__365__),
    .I0(__254__),
    .O(__1031__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __2119__ (
    .I3(__484__),
    .I2(__443__),
    .I1(__97__),
    .I0(__71__),
    .O(__1032__)
  );
  LUT5 #(
    .INIT(32'h00008000)
  ) __2120__ (
    .I4(__220__),
    .I3(__134__),
    .I2(__35__),
    .I1(__260__),
    .I0(__205__),
    .O(__1033__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __2121__ (
    .I2(__758__),
    .I1(__355__),
    .I0(__194__),
    .O(__1034__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __2122__ (
    .I1(__401__),
    .I0(__20__),
    .O(__1035__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __2123__ (
    .I2(__669__),
    .I1(__26__),
    .I0(__54__),
    .O(__1036__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __2124__ (
    .I3(__334__),
    .I2(__462__),
    .I1(__136__),
    .I0(__355__),
    .O(__1037__)
  );
  LUT6 #(
    .INIT(64'h7fff800000000000)
  ) __2125__ (
    .I5(__391__),
    .I4(__318__),
    .I3(__124__),
    .I2(__420__),
    .I1(__276__),
    .I0(__434__),
    .O(__1038__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __2126__ (
    .I3(__484__),
    .I2(__443__),
    .I1(__262__),
    .I0(__494__),
    .O(__1039__)
  );
  LUT4 #(
    .INIT(16'haa3c)
  ) __2127__ (
    .I3(__322__),
    .I2(__182__),
    .I1(__157__),
    .I0(__164__),
    .O(__1040__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __2128__ (
    .I2(__527__),
    .I1(__356__),
    .I0(__402__),
    .O(__1041__)
  );
  LUT3 #(
    .INIT(8'h10)
  ) __2129__ (
    .I2(g43),
    .I1(__778__),
    .I0(g1),
    .O(__1042__)
  );
  LUT4 #(
    .INIT(16'h7800)
  ) __2130__ (
    .I3(__391__),
    .I2(__124__),
    .I1(__276__),
    .I0(__434__),
    .O(__1043__)
  );
  LUT5 #(
    .INIT(32'h00008000)
  ) __2131__ (
    .I4(__205__),
    .I3(__134__),
    .I2(__35__),
    .I1(__260__),
    .I0(__220__),
    .O(__1044__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __2132__ (
    .I3(__419__),
    .I2(__82__),
    .I1(__161__),
    .I0(__256__),
    .O(__1045__)
  );
  LUT5 #(
    .INIT(32'hcaaaaaaa)
  ) __2133__ (
    .I4(__504__),
    .I3(__503__),
    .I2(__502__),
    .I1(__166__),
    .I0(__57__),
    .O(__1046__)
  );
  LUT6 #(
    .INIT(64'h9009000000009009)
  ) __2134__ (
    .I5(__156__),
    .I4(__440__),
    .I3(__348__),
    .I2(__318__),
    .I1(__233__),
    .I0(__124__),
    .O(__1047__)
  );
  LUT6 #(
    .INIT(64'h0000000000009009)
  ) __2135__ (
    .I5(__276__),
    .I4(__434__),
    .I3(__197__),
    .I2(__138__),
    .I1(__173__),
    .I0(__420__),
    .O(__1048__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __2136__ (
    .I1(__1048__),
    .I0(__1047__),
    .O(__1049__)
  );
  LUT4 #(
    .INIT(16'h9009)
  ) __2137__ (
    .I3(__272__),
    .I2(__352__),
    .I1(__222__),
    .I0(__404__),
    .O(__1050__)
  );
  LUT6 #(
    .INIT(64'h6ff6ffffffffffff)
  ) __2138__ (
    .I5(__1050__),
    .I4(__1049__),
    .I3(__454__),
    .I2(__202__),
    .I1(__233__),
    .I0(__108__),
    .O(__1051__)
  );
  LUT6 #(
    .INIT(64'hbfffffffeaaaaaaa)
  ) __2139__ (
    .I5(__167__),
    .I4(__188__),
    .I3(__248__),
    .I2(__145__),
    .I1(__500__),
    .I0(__258__),
    .O(__1052__)
  );
  LUT4 #(
    .INIT(16'haa3c)
  ) __2140__ (
    .I3(__322__),
    .I2(__90__),
    .I1(__816__),
    .I0(__360__),
    .O(__1053__)
  );
  LUT4 #(
    .INIT(16'h7800)
  ) __2141__ (
    .I3(__391__),
    .I2(__440__),
    .I1(__404__),
    .I0(__707__),
    .O(__1054__)
  );
  LUT5 #(
    .INIT(32'hcaaaaaaa)
  ) __2142__ (
    .I4(__504__),
    .I3(__503__),
    .I2(__536__),
    .I1(__379__),
    .I0(__209__),
    .O(__1055__)
  );
  LUT3 #(
    .INIT(8'h60)
  ) __2143__ (
    .I2(__391__),
    .I1(__276__),
    .I0(__434__),
    .O(__1056__)
  );
  LUT5 #(
    .INIT(32'hcaaaaaaa)
  ) __2144__ (
    .I4(__504__),
    .I3(__503__),
    .I2(__502__),
    .I1(__482__),
    .I0(__159__),
    .O(__1057__)
  );
  LUT2 #(
    .INIT(4'he)
  ) __2145__ (
    .I1(__215__),
    .I0(__284__),
    .O(__1058__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __2146__ (
    .I2(__719__),
    .I1(__405__),
    .I0(__206__),
    .O(__1059__)
  );
  LUT5 #(
    .INIT(32'h00004000)
  ) __2147__ (
    .I4(__425__),
    .I3(g43),
    .I2(__93__),
    .I1(__87__),
    .I0(__338__),
    .O(__1060__)
  );
  LUT3 #(
    .INIT(8'hfe)
  ) __2148__ (
    .I2(__258__),
    .I1(__468__),
    .I0(__18__),
    .O(__1061__)
  );
  LUT6 #(
    .INIT(64'h00007fff00008000)
  ) __2149__ (
    .I5(__279__),
    .I4(__380__),
    .I3(__319__),
    .I2(__185__),
    .I1(__130__),
    .I0(__569__),
    .O(__1062__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __2150__ (
    .I2(__665__),
    .I1(__116__),
    .I0(__217__),
    .O(__1063__)
  );
  LUT2 #(
    .INIT(4'hb)
  ) __2151__ (
    .I1(__313__),
    .I0(__626__),
    .O(__1064__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __2152__ (
    .I2(__575__),
    .I1(__405__),
    .I0(__328__),
    .O(__1065__)
  );
  LUT4 #(
    .INIT(16'h8000)
  ) __2153__ (
    .I3(__188__),
    .I2(__248__),
    .I1(__145__),
    .I0(__500__),
    .O(__1066__)
  );
  LUT4 #(
    .INIT(16'hf7f8)
  ) __2154__ (
    .I3(__345__),
    .I2(__258__),
    .I1(__167__),
    .I0(__1066__),
    .O(__1067__)
  );
  LUT3 #(
    .INIT(8'he2)
  ) __2155__ (
    .I2(__223__),
    .I1(__89__),
    .I0(g11),
    .O(__1068__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __2156__ (
    .I2(__719__),
    .I1(__312__),
    .I0(__477__),
    .O(__1069__)
  );
  LUT4 #(
    .INIT(16'h8000)
  ) __2157__ (
    .I3(__138__),
    .I2(__440__),
    .I1(__404__),
    .I0(__707__),
    .O(__1070__)
  );
  LUT4 #(
    .INIT(16'h7800)
  ) __2158__ (
    .I3(__391__),
    .I2(__108__),
    .I1(__352__),
    .I0(__1070__),
    .O(__1071__)
  );
  LUT5 #(
    .INIT(32'hfeff0000)
  ) __2159__ (
    .I4(__453__),
    .I3(__854__),
    .I2(__344__),
    .I1(__286__),
    .I0(__135__),
    .O(__1072__)
  );
  LUT6 #(
    .INIT(64'h3f3fffff33000302)
  ) __2160__ (
    .I5(__42__),
    .I4(__242__),
    .I3(__192__),
    .I2(__704__),
    .I1(__144__),
    .I0(__1072__),
    .O(__1073__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __2161__ (
    .I1(__334__),
    .I0(__462__),
    .O(__1074__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __2162__ (
    .I3(__74__),
    .I2(__489__),
    .I1(__104__),
    .I0(__410__),
    .O(__1075__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __2163__ (
    .I3(__484__),
    .I2(__443__),
    .I1(__451__),
    .I0(__191__),
    .O(__1076__)
  );
  LUT6 #(
    .INIT(64'h0000000000008000)
  ) __2164__ (
    .I5(__87__),
    .I4(__779__),
    .I3(__799__),
    .I2(__81__),
    .I1(g1),
    .I0(__19__),
    .O(__1077__)
  );
  LUT5 #(
    .INIT(32'hfef00000)
  ) __2165__ (
    .I4(__899__),
    .I3(__429__),
    .I2(__425__),
    .I1(__476__),
    .I0(__121__),
    .O(__1078__)
  );
  LUT5 #(
    .INIT(32'hcaaaaaaa)
  ) __2166__ (
    .I4(__504__),
    .I3(__503__),
    .I2(__536__),
    .I1(__165__),
    .I0(__155__),
    .O(__1079__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __2167__ (
    .I2(__541__),
    .I1(__306__),
    .I0(__86__),
    .O(__1080__)
  );
  LUT5 #(
    .INIT(32'h80000000)
  ) __2168__ (
    .I4(__232__),
    .I3(__361__),
    .I2(__311__),
    .I1(__187__),
    .I0(__721__),
    .O(__1081__)
  );
  LUT4 #(
    .INIT(16'h152a)
  ) __2169__ (
    .I3(__357__),
    .I2(__261__),
    .I1(__472__),
    .I0(__1081__),
    .O(__1082__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __2170__ (
    .I2(__541__),
    .I1(__377__),
    .I0(__310__),
    .O(__1083__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __2171__ (
    .I2(__162__),
    .I1(__122__),
    .I0(g1080),
    .O(__1084__)
  );
  LUT6 #(
    .INIT(64'hf0fbf0f0ffffffff)
  ) __2172__ (
    .I5(__313__),
    .I4(__533__),
    .I3(__664__),
    .I2(__674__),
    .I1(__662__),
    .I0(__530__),
    .O(__1085__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __2173__ (
    .I1(__179__),
    .I0(g955),
    .O(__1086__)
  );
  assign g4657 = __841__;
  assign g3191 = __82__;
  assign g785 = __144__;
  assign g6308 = g45;
  assign g4664 = __734__;
  assign g1195 = __31__;
  assign g7048 = __1008__;
  assign g7763 = __974__;
  assign g6909 = g1008;
  assign g6289 = g1;
  assign g9378 = __933__;
  assign g6212 = __354__;
  assign g7730 = __354__;
  assign g1817 = __23__;
  assign g206 = __78__;
  assign g291 = __78__;
  assign g372 = __78__;
  assign g453 = __78__;
  assign g534 = __78__;
  assign g594 = __78__;
  assign g7294 = __936__;
  assign g7295 = __936__;
  assign g7283 = __966__;
  assign g4663 = __1035__;
  assign g8872 = __981__;
  assign g6298 = g28;
  assign g6303 = g32;
  assign g6293 = g23;
  assign g6305 = g41;
  assign g3856 = __10__;
  assign g8661 = 1'b0;
  assign g6269 = g1000;
  assign g8958 = __943__;
  assign g8234 = __927__;
  assign g9132 = __927__;
  assign g3857 = __11__;
  assign g6425 = __87__;
  assign g8218 = __87__;
  assign g6236 = __1021__;
  assign g7731 = __1021__;
  assign g4372 = __320__;
  assign g4371 = __65__;
  assign g1894 = __239__;
  assign g4660 = __964__;
  assign g5669 = __273__;
  assign g7504 = __273__;
  assign g1201 = __234__;
  assign g6302 = g31;
  assign g3130 = __489__;
  assign g7424 = __221__;
  assign g6300 = g29;
  assign g9128 = __789__;
  assign g9204 = __789__;
  assign g6295 = g25;
  assign g6376 = g25;
  assign g9310 = __1064__;
  assign g7063 = __836__;
  assign g8663 = __836__;
  assign g5571 = __389__;
  assign g6849 = __857__;
  assign g6288 = g9;
  assign g9312 = __939__;
  assign g1824 = __135__;
  assign g9297 = __608__;
  assign g6290 = g11;
  assign g4316 = __457__;
  assign g1205 = __395__;
  assign g9299 = __565__;
  assign g5678 = __432__;
  assign g7505 = __432__;
  assign g3854 = __12__;
  assign g1911 = __475__;
  assign g5687 = __172__;
  assign g7508 = __172__;
  assign g3096 = __147__;
  assign g7290 = __511__;
  assign g6207 = __493__;
  assign g7729 = __493__;
  assign g1724 = __226__;
  assign g1944 = __162__;
  assign g7289 = __546__;
  assign g5729 = g49;
  assign g1804 = __200__;
  assign g7474 = __685__;
  assign g2662 = __103__;
  assign g6304 = g37;
  assign g1015 = __1077__;
  assign g6648 = __255__;
  assign g8216 = __255__;
  assign g1783 = __344__;
  assign g7425 = __251__;
  assign g2844 = __443__;
  assign g3159 = __443__;
  assign g7292 = __760__;
  assign g7288 = __887__;
  assign g6292 = g22;
  assign g7284 = __892__;
  assign g5143 = g1554;
  assign g7514 = __941__;
  assign g1810 = __213__;
  assign g9305 = __793__;
  assign g6306 = g42;
  assign g1870 = __24__;
  assign g6297 = g27;
  assign g1197 = __350__;
  assign g3829 = __366__;
  assign g3859 = __366__;
  assign g3860 = __366__;
  assign g6850 = __8__;
  assign g7293 = __711__;
  assign g6895 = __1__;
  assign g7103 = __934__;
  assign g9280 = __1085__;
  assign g4373 = __160__;
  assign g6223 = __6__;
  assign g7732 = __6__;
  assign g1006 = __831__;
  assign g6307 = g44;
  assign g9314 = __535__;
  assign g4267 = __472__;
  assign g1871 = __55__;
  assign g7298 = __935__;
  assign g1829 = __286__;
  assign g6675 = __4__;
  assign g8219 = __4__;
  assign g7423 = __163__;
  assign g6299 = g21;
  assign g6291 = g10;
  assign g7285 = __913__;
  assign g7286 = __681__;
  assign g4661 = __585__;
  assign g5682 = __418__;
  assign g7506 = __418__;
  assign g9308 = __825__;
  assign g7287 = __714__;
  assign g1017 = __425__;
  assign g3077 = __425__;
  assign g6294 = g24;
  assign g5164 = __1017__;
  assign g7291 = __850__;
  assign g6301 = g30;
  assign g1246 = __471__;
  assign g2888 = __91__;
  assign g1193 = __407__;
  assign g1798 = __151__;
  assign g6653 = __308__;
  assign g8217 = __308__;
  assign g4655 = __1074__;
  assign g5684 = __107__;
  assign g7507 = __107__;
  assign g6296 = g26;
  assign g4370 = __235__;
endmodule
