module s5378 (
  CK,
  n3065gat,
  n3066gat,
  n3067gat,
  n3068gat,
  n3069gat,
  n3070gat,
  n3071gat,
  n3072gat,
  n3073gat,
  n3074gat,
  n3075gat,
  n3076gat,
  n3077gat,
  n3078gat,
  n3079gat,
  n3080gat,
  n3081gat,
  n3082gat,
  n3083gat,
  n3084gat,
  n3085gat,
  n3086gat,
  n3087gat,
  n3088gat,
  n3089gat,
  n3090gat,
  n3091gat,
  n3092gat,
  n3093gat,
  n3094gat,
  n3095gat,
  n3097gat,
  n3098gat,
  n3099gat,
  n3100gat,
  n3150gat,
  n3127gat,
  n3133gat,
  n3149gat,
  n3125gat,
  n3118gat,
  n3143gat,
  n3146gat,
  n3123gat,
  n3132gat,
  n3106gat,
  n3119gat,
  n3124gat,
  n3136gat,
  n3145gat,
  n3117gat,
  n3114gat,
  n3104gat,
  n3134gat,
  n3128gat,
  n3116gat,
  n3105gat,
  n3120gat,
  n3126gat,
  n3121gat,
  n3135gat,
  n3144gat,
  n3108gat,
  n3113gat,
  n3107gat,
  n3109gat,
  n3131gat,
  n3137gat,
  n3111gat,
  n3110gat,
  n3138gat,
  n3130gat,
  n3129gat,
  n3151gat,
  n3141gat,
  n3142gat,
  n3112gat,
  n3115gat,
  n3147gat,
  n3148gat,
  n3152gat,
  n3139gat,
  n3140gat,
  n3122gat
);
  input CK;
  wire CK;
  input n3065gat;
  wire n3065gat;
  input n3066gat;
  wire n3066gat;
  input n3067gat;
  wire n3067gat;
  input n3068gat;
  wire n3068gat;
  input n3069gat;
  wire n3069gat;
  input n3070gat;
  wire n3070gat;
  input n3071gat;
  wire n3071gat;
  input n3072gat;
  wire n3072gat;
  input n3073gat;
  wire n3073gat;
  input n3074gat;
  wire n3074gat;
  input n3075gat;
  wire n3075gat;
  input n3076gat;
  wire n3076gat;
  input n3077gat;
  wire n3077gat;
  input n3078gat;
  wire n3078gat;
  input n3079gat;
  wire n3079gat;
  input n3080gat;
  wire n3080gat;
  input n3081gat;
  wire n3081gat;
  input n3082gat;
  wire n3082gat;
  input n3083gat;
  wire n3083gat;
  input n3084gat;
  wire n3084gat;
  input n3085gat;
  wire n3085gat;
  input n3086gat;
  wire n3086gat;
  input n3087gat;
  wire n3087gat;
  input n3088gat;
  wire n3088gat;
  input n3089gat;
  wire n3089gat;
  input n3090gat;
  wire n3090gat;
  input n3091gat;
  wire n3091gat;
  input n3092gat;
  wire n3092gat;
  input n3093gat;
  wire n3093gat;
  input n3094gat;
  wire n3094gat;
  input n3095gat;
  wire n3095gat;
  input n3097gat;
  wire n3097gat;
  input n3098gat;
  wire n3098gat;
  input n3099gat;
  wire n3099gat;
  input n3100gat;
  wire n3100gat;
  output n3150gat;
  wire n3150gat;
  output n3127gat;
  wire n3127gat;
  output n3133gat;
  wire n3133gat;
  output n3149gat;
  wire n3149gat;
  output n3125gat;
  wire n3125gat;
  output n3118gat;
  wire n3118gat;
  output n3143gat;
  wire n3143gat;
  output n3146gat;
  wire n3146gat;
  output n3123gat;
  wire n3123gat;
  output n3132gat;
  wire n3132gat;
  output n3106gat;
  wire n3106gat;
  output n3119gat;
  wire n3119gat;
  output n3124gat;
  wire n3124gat;
  output n3136gat;
  wire n3136gat;
  output n3145gat;
  wire n3145gat;
  output n3117gat;
  wire n3117gat;
  output n3114gat;
  wire n3114gat;
  output n3104gat;
  wire n3104gat;
  output n3134gat;
  wire n3134gat;
  output n3128gat;
  wire n3128gat;
  output n3116gat;
  wire n3116gat;
  output n3105gat;
  wire n3105gat;
  output n3120gat;
  wire n3120gat;
  output n3126gat;
  wire n3126gat;
  output n3121gat;
  wire n3121gat;
  output n3135gat;
  wire n3135gat;
  output n3144gat;
  wire n3144gat;
  output n3108gat;
  wire n3108gat;
  output n3113gat;
  wire n3113gat;
  output n3107gat;
  wire n3107gat;
  output n3109gat;
  wire n3109gat;
  output n3131gat;
  wire n3131gat;
  output n3137gat;
  wire n3137gat;
  output n3111gat;
  wire n3111gat;
  output n3110gat;
  wire n3110gat;
  output n3138gat;
  wire n3138gat;
  output n3130gat;
  wire n3130gat;
  output n3129gat;
  wire n3129gat;
  output n3151gat;
  wire n3151gat;
  output n3141gat;
  wire n3141gat;
  output n3142gat;
  wire n3142gat;
  output n3112gat;
  wire n3112gat;
  output n3115gat;
  wire n3115gat;
  output n3147gat;
  wire n3147gat;
  output n3148gat;
  wire n3148gat;
  output n3152gat;
  wire n3152gat;
  output n3139gat;
  wire n3139gat;
  output n3140gat;
  wire n3140gat;
  output n3122gat;
  wire n3122gat;
  wire __0__;
  wire __1__;
  wire __2__;
  wire __3__;
  wire __4__;
  wire __5__;
  wire __6__;
  wire __7__;
  wire __8__;
  wire __9__;
  wire __10__;
  wire __11__;
  wire __12__;
  wire __13__;
  wire __14__;
  wire __15__;
  wire __16__;
  wire __17__;
  wire __18__;
  wire __19__;
  wire __20__;
  wire __21__;
  wire __22__;
  wire __23__;
  wire __24__;
  wire __25__;
  wire __26__;
  wire __27__;
  wire __28__;
  wire __29__;
  wire __30__;
  wire __31__;
  wire __32__;
  wire __33__;
  wire __34__;
  wire __35__;
  wire __36__;
  wire __37__;
  wire __38__;
  wire __39__;
  wire __40__;
  wire __41__;
  wire __42__;
  wire __43__;
  wire __44__;
  wire __45__;
  wire __46__;
  wire __47__;
  wire __48__;
  wire __49__;
  wire __50__;
  wire __51__;
  wire __52__;
  wire __53__;
  wire __54__;
  wire __55__;
  wire __56__;
  wire __57__;
  wire __58__;
  wire __59__;
  wire __60__;
  wire __61__;
  wire __62__;
  wire __63__;
  wire __64__;
  wire __65__;
  wire __66__;
  wire __67__;
  wire __68__;
  wire __69__;
  wire __70__;
  wire __71__;
  wire __72__;
  wire __73__;
  wire __74__;
  wire __75__;
  wire __76__;
  wire __77__;
  wire __78__;
  wire __79__;
  wire __80__;
  wire __81__;
  wire __82__;
  wire __83__;
  wire __84__;
  wire __85__;
  wire __86__;
  wire __87__;
  wire __88__;
  wire __89__;
  wire __90__;
  wire __91__;
  wire __92__;
  wire __93__;
  wire __94__;
  wire __95__;
  wire __96__;
  wire __97__;
  wire __98__;
  wire __99__;
  wire __100__;
  wire __101__;
  wire __102__;
  wire __103__;
  wire __104__;
  wire __105__;
  wire __106__;
  wire __107__;
  wire __108__;
  wire __109__;
  wire __110__;
  wire __111__;
  wire __112__;
  wire __113__;
  wire __114__;
  wire __115__;
  wire __116__;
  wire __117__;
  wire __118__;
  wire __119__;
  wire __120__;
  wire __121__;
  wire __122__;
  wire __123__;
  wire __124__;
  wire __125__;
  wire __126__;
  wire __127__;
  wire __128__;
  wire __129__;
  wire __130__;
  wire __131__;
  wire __132__;
  wire __133__;
  wire __134__;
  wire __135__;
  wire __136__;
  wire __137__;
  wire __138__;
  wire __139__;
  wire __140__;
  wire __141__;
  wire __142__;
  wire __143__;
  wire __144__;
  wire __145__;
  wire __146__;
  wire __147__;
  wire __148__;
  wire __149__;
  wire __150__;
  wire __151__;
  wire __152__;
  wire __153__;
  wire __154__;
  wire __155__;
  wire __156__;
  wire __157__;
  wire __158__;
  wire __159__;
  wire __160__;
  wire __161__;
  wire __162__;
  wire __163__;
  wire __164__;
  wire __165__;
  wire __166__;
  wire __167__;
  wire __168__;
  wire __169__;
  wire __170__;
  wire __171__;
  wire __172__;
  wire __173__;
  wire __174__;
  wire __175__;
  wire __176__;
  wire __177__;
  wire __178__;
  wire __179__;
  wire __180__;
  wire __181__;
  wire __182__;
  wire __183__;
  wire __184__;
  wire __185__;
  wire __186__;
  wire __187__;
  wire __188__;
  wire __189__;
  wire __190__;
  wire __191__;
  wire __192__;
  wire __193__;
  wire __194__;
  wire __195__;
  wire __196__;
  wire __197__;
  wire __198__;
  wire __199__;
  wire __200__;
  wire __201__;
  wire __202__;
  wire __203__;
  wire __204__;
  wire __205__;
  wire __206__;
  wire __209__;
  wire __210__;
  wire __211__;
  wire __212__;
  wire __213__;
  wire __214__;
  wire __215__;
  wire __216__;
  wire __217__;
  wire __218__;
  wire __219__;
  wire __220__;
  wire __221__;
  wire __222__;
  wire __223__;
  wire __224__;
  wire __225__;
  wire __226__;
  wire __227__;
  wire __228__;
  wire __229__;
  wire __230__;
  wire __231__;
  wire __232__;
  wire __233__;
  wire __234__;
  wire __235__;
  wire __236__;
  wire __237__;
  wire __238__;
  wire __239__;
  wire __240__;
  wire __241__;
  wire __242__;
  wire __243__;
  wire __244__;
  wire __245__;
  wire __246__;
  wire __247__;
  wire __248__;
  wire __249__;
  wire __250__;
  wire __251__;
  wire __252__;
  wire __253__;
  wire __254__;
  wire __255__;
  wire __256__;
  wire __257__;
  wire __258__;
  wire __259__;
  wire __260__;
  wire __261__;
  wire __262__;
  wire __263__;
  wire __264__;
  wire __265__;
  wire __266__;
  wire __267__;
  wire __268__;
  wire __269__;
  wire __270__;
  wire __271__;
  wire __272__;
  wire __273__;
  wire __274__;
  wire __275__;
  wire __276__;
  wire __277__;
  wire __278__;
  wire __279__;
  wire __280__;
  wire __281__;
  wire __282__;
  wire __283__;
  wire __284__;
  wire __285__;
  wire __286__;
  wire __287__;
  wire __288__;
  wire __289__;
  wire __290__;
  wire __291__;
  wire __292__;
  wire __293__;
  wire __294__;
  wire __295__;
  wire __296__;
  wire __297__;
  wire __298__;
  wire __299__;
  wire __300__;
  wire __301__;
  wire __302__;
  wire __303__;
  wire __304__;
  wire __305__;
  wire __306__;
  wire __307__;
  wire __308__;
  wire __309__;
  wire __310__;
  wire __311__;
  wire __312__;
  wire __313__;
  wire __314__;
  wire __315__;
  wire __316__;
  wire __317__;
  wire __318__;
  wire __319__;
  wire __320__;
  wire __321__;
  wire __322__;
  wire __323__;
  wire __324__;
  wire __325__;
  wire __326__;
  wire __327__;
  wire __328__;
  wire __329__;
  wire __330__;
  wire __331__;
  wire __332__;
  wire __333__;
  wire __334__;
  wire __335__;
  wire __336__;
  wire __337__;
  wire __338__;
  wire __339__;
  wire __340__;
  wire __341__;
  wire __342__;
  wire __343__;
  wire __344__;
  wire __345__;
  wire __346__;
  wire __347__;
  wire __348__;
  wire __349__;
  wire __350__;
  wire __351__;
  wire __352__;
  wire __353__;
  wire __354__;
  wire __355__;
  wire __356__;
  wire __357__;
  wire __358__;
  wire __359__;
  wire __360__;
  wire __361__;
  wire __362__;
  wire __363__;
  wire __364__;
  wire __365__;
  wire __366__;
  wire __367__;
  wire __368__;
  wire __369__;
  wire __370__;
  wire __371__;
  wire __372__;
  wire __373__;
  wire __374__;
  wire __375__;
  wire __376__;
  wire __377__;
  wire __378__;
  wire __379__;
  wire __380__;
  wire __381__;
  wire __382__;
  wire __383__;
  wire __384__;
  wire __385__;
  wire __386__;
  wire __387__;
  wire __388__;
  wire __389__;
  wire __390__;
  wire __391__;
  wire __392__;
  wire __393__;
  wire __394__;
  wire __395__;
  wire __396__;
  wire __397__;
  wire __398__;
  wire __399__;
  wire __400__;
  wire __401__;
  wire __402__;
  wire __403__;
  wire __404__;
  wire __405__;
  wire __406__;
  wire __407__;
  wire __408__;
  wire __409__;
  wire __410__;
  wire __411__;
  wire __412__;
  wire __413__;
  wire __414__;
  wire __415__;
  wire __416__;
  wire __417__;
  wire __418__;
  wire __419__;
  wire __420__;
  wire __421__;
  wire __422__;
  wire __423__;
  wire __424__;
  wire __425__;
  wire __426__;
  wire __427__;
  wire __428__;
  wire __429__;
  wire __430__;
  wire __431__;
  wire __432__;
  wire __433__;
  wire __434__;
  wire __435__;
  wire __436__;
  wire __437__;
  wire __438__;
  wire __439__;
  wire __440__;
  wire __441__;
  wire __442__;
  wire __443__;
  wire __444__;
  wire __445__;
  wire __446__;
  wire __447__;
  wire __448__;
  wire __449__;
  wire __450__;
  wire __451__;
  wire __452__;
  wire __453__;
  wire __454__;
  wire __455__;
  wire __456__;
  wire __457__;
  wire __458__;
  wire __459__;
  wire __460__;
  wire __461__;
  wire __462__;
  wire __463__;
  wire __464__;
  wire __465__;
  wire __466__;
  wire __467__;
  wire __468__;
  wire __469__;
  wire __470__;
  wire __471__;
  wire __472__;
  wire __473__;
  wire __474__;
  wire __475__;
  wire __476__;
  wire __477__;
  wire __478__;
  wire __479__;
  wire __480__;
  wire __481__;
  wire __482__;
  wire __483__;
  wire __484__;
  wire __485__;
  wire __486__;
  wire __487__;
  wire __488__;
  wire __489__;
  wire __490__;
  wire __491__;
  wire __492__;
  wire __493__;
  wire __494__;
  wire __495__;
  wire __496__;
  wire __497__;
  wire __498__;
  wire __499__;
  wire __500__;
  wire __501__;
  wire __502__;
  wire __503__;
  wire __504__;
  wire __505__;
  wire __506__;
  wire __507__;
  wire __508__;
  wire __509__;
  wire __510__;
  INV __511__ (
    .I(__196__),
    .O(__0__)
  );
  INV __512__ (
    .I(__192__),
    .O(__1__)
  );
  INV __513__ (
    .I(__189__),
    .O(__2__)
  );
  INV __514__ (
    .I(__50__),
    .O(__3__)
  );
  INV __515__ (
    .I(__180__),
    .O(__4__)
  );
  INV __516__ (
    .I(__53__),
    .O(__5__)
  );
  INV __517__ (
    .I(__174__),
    .O(__6__)
  );
  INV __518__ (
    .I(__170__),
    .O(__7__)
  );
  INV __519__ (
    .I(__124__),
    .O(__8__)
  );
  INV __520__ (
    .I(__52__),
    .O(__9__)
  );
  INV __521__ (
    .I(__141__),
    .O(__10__)
  );
  INV __522__ (
    .I(__56__),
    .O(__11__)
  );
  INV __523__ (
    .I(__197__),
    .O(__12__)
  );
  INV __524__ (
    .I(__193__),
    .O(__13__)
  );
  INV __525__ (
    .I(__191__),
    .O(__14__)
  );
  INV __526__ (
    .I(__190__),
    .O(__15__)
  );
  INV __527__ (
    .I(__187__),
    .O(__16__)
  );
  INV __528__ (
    .I(__184__),
    .O(__17__)
  );
  INV __529__ (
    .I(__183__),
    .O(__18__)
  );
  INV __530__ (
    .I(__185__),
    .O(__19__)
  );
  INV __531__ (
    .I(__177__),
    .O(__20__)
  );
  INV __532__ (
    .I(__182__),
    .O(__21__)
  );
  INV __533__ (
    .I(__123__),
    .O(__22__)
  );
  INV __534__ (
    .I(__135__),
    .O(__23__)
  );
  INV __535__ (
    .I(__134__),
    .O(__24__)
  );
  INV __536__ (
    .I(__133__),
    .O(__25__)
  );
  INV __537__ (
    .I(__49__),
    .O(__26__)
  );
  INV __538__ (
    .I(__186__),
    .O(__27__)
  );
  INV __539__ (
    .I(__129__),
    .O(__28__)
  );
  INV __540__ (
    .I(__113__),
    .O(__29__)
  );
  INV __541__ (
    .I(__145__),
    .O(__30__)
  );
  INV __542__ (
    .I(__100__),
    .O(__31__)
  );
  INV __543__ (
    .I(__102__),
    .O(__32__)
  );
  INV __544__ (
    .I(__101__),
    .O(__33__)
  );
  INV __545__ (
    .I(__98__),
    .O(__34__)
  );
  INV __546__ (
    .I(__97__),
    .O(__35__)
  );
  INV __547__ (
    .I(__93__),
    .O(__36__)
  );
  INV __548__ (
    .I(__92__),
    .O(__37__)
  );
  INV __549__ (
    .I(__88__),
    .O(__38__)
  );
  INV __550__ (
    .I(__87__),
    .O(__39__)
  );
  INV __551__ (
    .I(__86__),
    .O(__40__)
  );
  INV __552__ (
    .I(__144__),
    .O(__41__)
  );
  INV __553__ (
    .I(__55__),
    .O(__42__)
  );
  INV __554__ (
    .I(__54__),
    .O(__43__)
  );
  INV __555__ (
    .I(__85__),
    .O(__44__)
  );
  INV __556__ (
    .I(__94__),
    .O(__45__)
  );
  INV __557__ (
    .I(__72__),
    .O(__46__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __558__ (
    .D(n3070gat),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__47__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __559__ (
    .D(__451__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__48__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __560__ (
    .D(__283__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__49__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __561__ (
    .D(__489__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__50__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __562__ (
    .D(__390__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__51__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __563__ (
    .D(__505__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__52__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __564__ (
    .D(__357__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__53__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __565__ (
    .D(__42__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__54__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __566__ (
    .D(__41__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__55__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __567__ (
    .D(__239__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__56__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __568__ (
    .D(__228__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__57__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __569__ (
    .D(__412__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__58__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __570__ (
    .D(__40__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__59__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __571__ (
    .D(__46__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__60__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __572__ (
    .D(__3__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__61__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __573__ (
    .D(__501__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__62__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __574__ (
    .D(__269__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__63__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __575__ (
    .D(__272__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__64__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __576__ (
    .D(__446__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__65__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __577__ (
    .D(__431__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__66__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __578__ (
    .D(__460__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__67__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __579__ (
    .D(__481__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__68__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __580__ (
    .D(__426__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__69__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __581__ (
    .D(__265__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__70__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __582__ (
    .D(__467__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__71__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __583__ (
    .D(__45__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__72__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __584__ (
    .D(__5__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__73__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __585__ (
    .D(__6__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__74__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __586__ (
    .D(__4__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__75__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __587__ (
    .D(__12__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__76__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __588__ (
    .D(__11__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__77__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __589__ (
    .D(__8__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__78__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __590__ (
    .D(__9__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__79__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __591__ (
    .D(__10__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__80__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __592__ (
    .D(__7__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__81__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __593__ (
    .D(__28__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__82__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __594__ (
    .D(__44__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__83__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __595__ (
    .D(__22__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__84__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __596__ (
    .D(__43__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__85__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __597__ (
    .D(__411__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__86__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __598__ (
    .D(__38__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__87__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __599__ (
    .D(__421__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__88__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __600__ (
    .D(__398__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__89__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __601__ (
    .D(__224__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__90__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __602__ (
    .D(__37__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__91__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __603__ (
    .D(__36__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__92__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __604__ (
    .D(__483__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__93__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __605__ (
    .D(__34__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__94__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __606__ (
    .D(__478__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__95__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __607__ (
    .D(__261__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__96__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __608__ (
    .D(__422__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__97__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __609__ (
    .D(__388__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__98__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __610__ (
    .D(__33__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__99__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __611__ (
    .D(__270__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__100__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __612__ (
    .D(__32__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__101__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __613__ (
    .D(__31__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__102__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __614__ (
    .D(__482__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__103__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __615__ (
    .D(__24__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__104__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __616__ (
    .D(__26__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__105__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __617__ (
    .D(__25__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__106__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __618__ (
    .D(__30__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__107__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __619__ (
    .D(__231__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__108__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __620__ (
    .D(__504__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__109__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __621__ (
    .D(__500__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__110__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __622__ (
    .D(__229__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__111__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __623__ (
    .D(__29__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__112__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __624__ (
    .D(__361__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__113__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __625__ (
    .D(__424__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__114__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __626__ (
    .D(__15__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__115__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __627__ (
    .D(__17__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__116__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __628__ (
    .D(__16__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__117__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __629__ (
    .D(__13__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__118__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __630__ (
    .D(__19__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__119__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __631__ (
    .D(__18__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__120__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __632__ (
    .D(__21__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__121__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __633__ (
    .D(__27__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__122__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __634__ (
    .D(__485__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__123__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __635__ (
    .D(__414__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__124__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __636__ (
    .D(__20__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__125__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __637__ (
    .D(__372__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__126__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __638__ (
    .D(__385__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__127__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __639__ (
    .D(__209__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__128__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __640__ (
    .D(__280__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__129__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __641__ (
    .D(__220__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__130__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __642__ (
    .D(__230__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__131__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __643__ (
    .D(__346__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__132__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __644__ (
    .D(__406__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__133__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __645__ (
    .D(__275__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__134__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __646__ (
    .D(__353__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__135__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __647__ (
    .D(__336__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__136__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __648__ (
    .D(__470__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__137__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __649__ (
    .D(__285__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__138__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __650__ (
    .D(__378__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__139__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __651__ (
    .D(__391__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__140__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __652__ (
    .D(__366__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__141__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __653__ (
    .D(__490__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__142__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __654__ (
    .D(__23__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__143__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __655__ (
    .D(__39__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__144__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __656__ (
    .D(__284__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__145__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __657__ (
    .D(__14__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__146__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __658__ (
    .D(__458__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__147__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __659__ (
    .D(__395__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__148__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __660__ (
    .D(n3069gat),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__149__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __661__ (
    .D(__497__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__150__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __662__ (
    .D(__499__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__151__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __663__ (
    .D(__423__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__152__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __664__ (
    .D(__341__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__153__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __665__ (
    .D(__425__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__154__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __666__ (
    .D(__510__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__155__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __667__ (
    .D(__370__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__156__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __668__ (
    .D(__226__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__157__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __669__ (
    .D(__443__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__158__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __670__ (
    .D(__409__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__159__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __671__ (
    .D(__455__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__160__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __672__ (
    .D(__471__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__161__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __673__ (
    .D(__493__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__162__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __674__ (
    .D(__445__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__163__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __675__ (
    .D(__509__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__164__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __676__ (
    .D(__377__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__165__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __677__ (
    .D(__389__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__166__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __678__ (
    .D(__487__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__167__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __679__ (
    .D(__210__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__168__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __680__ (
    .D(__456__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__169__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __681__ (
    .D(__437__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__170__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __682__ (
    .D(__386__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__171__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __683__ (
    .D(__407__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__172__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __684__ (
    .D(__219__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__173__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __685__ (
    .D(__492__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__174__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __686__ (
    .D(__362__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__175__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __687__ (
    .D(__392__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__176__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __688__ (
    .D(__461__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__177__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __689__ (
    .D(__459__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__178__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __690__ (
    .D(__457__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__179__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __691__ (
    .D(__477__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__180__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __692__ (
    .D(__440__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__181__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __693__ (
    .D(__282__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__182__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __694__ (
    .D(__358__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__183__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __695__ (
    .D(__379__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__184__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __696__ (
    .D(__276__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__185__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __697__ (
    .D(__488__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__186__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __698__ (
    .D(__301__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__187__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __699__ (
    .D(__2__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__188__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __700__ (
    .D(__1__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__189__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __701__ (
    .D(__503__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__190__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __702__ (
    .D(__486__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__191__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __703__ (
    .D(__472__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__192__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __704__ (
    .D(__506__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__193__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __705__ (
    .D(__474__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__194__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __706__ (
    .D(__0__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__195__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __707__ (
    .D(__479__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__196__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __708__ (
    .D(__496__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__197__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __709__ (
    .D(__247__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__198__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __710__ (
    .D(n3068gat),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__199__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __711__ (
    .D(n3073gat),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__200__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __712__ (
    .D(n3066gat),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__201__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __713__ (
    .D(n3067gat),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__202__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __714__ (
    .D(n3065gat),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__203__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __715__ (
    .D(__434__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__204__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __716__ (
    .D(n3071gat),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__205__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __717__ (
    .D(n3072gat),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__206__)
  );
  LUT6 #(
    .INIT(64'h9669699669969669)
  ) __720__ (
    .I5(__185__),
    .I4(__182__),
    .I3(__177__),
    .I2(__183__),
    .I1(__186__),
    .I0(__129__),
    .O(__209__)
  );
  LUT4 #(
    .INIT(16'heac0)
  ) __721__ (
    .I3(n3093gat),
    .I2(n3095gat),
    .I1(n3082gat),
    .I0(n3073gat),
    .O(__210__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __722__ (
    .I1(__149__),
    .I0(__47__),
    .O(__211__)
  );
  LUT6 #(
    .INIT(64'hbeffffbeffffffff)
  ) __723__ (
    .I5(__211__),
    .I4(__117__),
    .I3(__206__),
    .I2(__146__),
    .I1(__205__),
    .I0(__116__),
    .O(__212__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __724__ (
    .I1(__149__),
    .I0(__47__),
    .O(__213__)
  );
  LUT6 #(
    .INIT(64'hbeffffbeffffffff)
  ) __725__ (
    .I5(__213__),
    .I4(__117__),
    .I3(__206__),
    .I2(__146__),
    .I1(__205__),
    .I0(__116__),
    .O(__214__)
  );
  LUT3 #(
    .INIT(8'h40)
  ) __726__ (
    .I2(__117__),
    .I1(__146__),
    .I0(__116__),
    .O(__215__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __727__ (
    .I1(__121__),
    .I0(__120__),
    .O(__216__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __728__ (
    .I1(__125__),
    .I0(__122__),
    .O(__217__)
  );
  LUT5 #(
    .INIT(32'h00000040)
  ) __729__ (
    .I4(__121__),
    .I3(__120__),
    .I2(__125__),
    .I1(__119__),
    .I0(__122__),
    .O(__218__)
  );
  LUT3 #(
    .INIT(8'h1f)
  ) __730__ (
    .I2(__176__),
    .I1(__178__),
    .I0(__57__),
    .O(__219__)
  );
  LUT3 #(
    .INIT(8'h7f)
  ) __731__ (
    .I2(__57__),
    .I1(__131__),
    .I0(__126__),
    .O(__220__)
  );
  LUT6 #(
    .INIT(64'h4040ff0000000000)
  ) __732__ (
    .I5(__220__),
    .I4(__219__),
    .I3(__218__),
    .I2(__217__),
    .I1(__216__),
    .I0(__119__),
    .O(__221__)
  );
  LUT6 #(
    .INIT(64'h3355f00000000000)
  ) __733__ (
    .I5(__221__),
    .I4(__115__),
    .I3(__118__),
    .I2(__215__),
    .I1(__214__),
    .I0(__212__),
    .O(__222__)
  );
  LUT6 #(
    .INIT(64'h000000007fffffff)
  ) __734__ (
    .I5(n3100gat),
    .I4(__128__),
    .I3(__132__),
    .I2(__136__),
    .I1(__137__),
    .I0(__204__),
    .O(__223__)
  );
  LUT4 #(
    .INIT(16'h0004)
  ) __735__ (
    .I3(__223__),
    .I2(__222__),
    .I1(__99__),
    .I0(__91__),
    .O(__224__)
  );
  LUT6 #(
    .INIT(64'h9669699669969669)
  ) __736__ (
    .I5(__155__),
    .I4(__168__),
    .I3(__164__),
    .I2(__159__),
    .I1(__161__),
    .I0(__169__),
    .O(__225__)
  );
  LUT4 #(
    .INIT(16'h9669)
  ) __737__ (
    .I3(__181__),
    .I2(__175__),
    .I1(__179__),
    .I0(__225__),
    .O(__226__)
  );
  LUT3 #(
    .INIT(8'h70)
  ) __738__ (
    .I2(__97__),
    .I1(__147__),
    .I0(__98__),
    .O(__227__)
  );
  LUT3 #(
    .INIT(8'h40)
  ) __739__ (
    .I2(n3100gat),
    .I1(__83__),
    .I0(__54__),
    .O(__228__)
  );
  LUT5 #(
    .INIT(32'h07080000)
  ) __740__ (
    .I4(__205__),
    .I3(__149__),
    .I2(__90__),
    .I1(__206__),
    .I0(__47__),
    .O(__229__)
  );
  LUT5 #(
    .INIT(32'h00000040)
  ) __741__ (
    .I4(__205__),
    .I3(__90__),
    .I2(__206__),
    .I1(__149__),
    .I0(__47__),
    .O(__230__)
  );
  LUT5 #(
    .INIT(32'h10001000)
  ) __742__ (
    .I4(__206__),
    .I3(__205__),
    .I2(__149__),
    .I1(__90__),
    .I0(__47__),
    .O(__231__)
  );
  LUT5 #(
    .INIT(32'h00004000)
  ) __743__ (
    .I4(__90__),
    .I3(__206__),
    .I2(__205__),
    .I1(__149__),
    .I0(__47__),
    .O(__232__)
  );
  LUT3 #(
    .INIT(8'h04)
  ) __744__ (
    .I2(__79__),
    .I1(__232__),
    .I0(__80__),
    .O(__233__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __745__ (
    .I1(n3092gat),
    .I0(n3091gat),
    .O(__234__)
  );
  LUT4 #(
    .INIT(16'h0040)
  ) __746__ (
    .I3(n3083gat),
    .I2(n3093gat),
    .I1(__97__),
    .I0(n3084gat),
    .O(__235__)
  );
  LUT6 #(
    .INIT(64'h0000000000004000)
  ) __747__ (
    .I5(n3086gat),
    .I4(n3088gat),
    .I3(n3087gat),
    .I2(n3085gat),
    .I1(__235__),
    .I0(__234__),
    .O(__236__)
  );
  LUT6 #(
    .INIT(64'h0000000000004000)
  ) __748__ (
    .I5(n3085gat),
    .I4(n3083gat),
    .I3(n3095gat),
    .I2(n3088gat),
    .I1(__97__),
    .I0(n3084gat),
    .O(__237__)
  );
  LUT4 #(
    .INIT(16'h4000)
  ) __749__ (
    .I3(n3086gat),
    .I2(n3094gat),
    .I1(__237__),
    .I0(n3087gat),
    .O(__238__)
  );
  LUT6 #(
    .INIT(64'heeeeaaaaccccf00f)
  ) __750__ (
    .I5(__238__),
    .I4(__236__),
    .I3(__77__),
    .I2(__233__),
    .I1(n3070gat),
    .I0(n3079gat),
    .O(__239__)
  );
  LUT6 #(
    .INIT(64'h033000a000000000)
  ) __751__ (
    .I5(n3086gat),
    .I4(n3095gat),
    .I3(n3087gat),
    .I2(n3093gat),
    .I1(n3088gat),
    .I0(n3085gat),
    .O(__240__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __752__ (
    .I1(__240__),
    .I0(__151__),
    .O(__241__)
  );
  LUT6 #(
    .INIT(64'h033000a000000000)
  ) __753__ (
    .I5(n3087gat),
    .I4(n3093gat),
    .I3(n3086gat),
    .I2(n3095gat),
    .I1(n3085gat),
    .I0(n3088gat),
    .O(__242__)
  );
  LUT6 #(
    .INIT(64'hfcc0a000a0000000)
  ) __754__ (
    .I5(n3093gat),
    .I4(n3087gat),
    .I3(n3095gat),
    .I2(n3086gat),
    .I1(n3085gat),
    .I0(n3088gat),
    .O(__243__)
  );
  LUT4 #(
    .INIT(16'hb0bb)
  ) __755__ (
    .I3(__243__),
    .I2(__201__),
    .I1(__242__),
    .I0(__175__),
    .O(__244__)
  );
  LUT2 #(
    .INIT(4'h9)
  ) __756__ (
    .I1(__206__),
    .I0(__205__),
    .O(__245__)
  );
  LUT3 #(
    .INIT(8'h96)
  ) __757__ (
    .I2(__203__),
    .I1(__201__),
    .I0(__202__),
    .O(__246__)
  );
  LUT6 #(
    .INIT(64'h9669699669969669)
  ) __758__ (
    .I5(__200__),
    .I4(__149__),
    .I3(__47__),
    .I2(__199__),
    .I1(__246__),
    .I0(__245__),
    .O(__247__)
  );
  LUT4 #(
    .INIT(16'h0004)
  ) __759__ (
    .I3(n3085gat),
    .I2(n3083gat),
    .I1(n3095gat),
    .I0(n3084gat),
    .O(__248__)
  );
  LUT6 #(
    .INIT(64'h00080c0000a00000)
  ) __760__ (
    .I5(n3093gat),
    .I4(n3095gat),
    .I3(n3087gat),
    .I2(n3086gat),
    .I1(n3085gat),
    .I0(n3088gat),
    .O(__249__)
  );
  LUT6 #(
    .INIT(64'hbfff0f0fbfbf0f0f)
  ) __761__ (
    .I5(__249__),
    .I4(__248__),
    .I3(__127__),
    .I2(__247__),
    .I1(__244__),
    .I0(__241__),
    .O(__250__)
  );
  LUT6 #(
    .INIT(64'h6996966996696996)
  ) __762__ (
    .I5(__110__),
    .I4(__140__),
    .I3(__139__),
    .I2(__148__),
    .I1(__150__),
    .I0(__152__),
    .O(__251__)
  );
  LUT3 #(
    .INIT(8'h69)
  ) __763__ (
    .I2(__154__),
    .I1(__151__),
    .I0(__251__),
    .O(__252__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __764__ (
    .I1(__249__),
    .I0(__124__),
    .O(__253__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __765__ (
    .I1(__242__),
    .I0(__168__),
    .O(__254__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __766__ (
    .I1(__243__),
    .I0(__200__),
    .O(__255__)
  );
  LUT6 #(
    .INIT(64'h0011000000000c00)
  ) __767__ (
    .I5(n3093gat),
    .I4(n3086gat),
    .I3(n3095gat),
    .I2(n3088gat),
    .I1(n3087gat),
    .I0(n3085gat),
    .O(__256__)
  );
  LUT6 #(
    .INIT(64'h0000007000440000)
  ) __768__ (
    .I5(n3093gat),
    .I4(n3086gat),
    .I3(n3087gat),
    .I2(n3085gat),
    .I1(n3095gat),
    .I0(n3088gat),
    .O(__257__)
  );
  LUT3 #(
    .INIT(8'h07)
  ) __769__ (
    .I2(__257__),
    .I1(__256__),
    .I0(__155__),
    .O(__258__)
  );
  LUT6 #(
    .INIT(64'h0000000700000000)
  ) __770__ (
    .I5(__258__),
    .I4(__255__),
    .I3(__254__),
    .I2(__253__),
    .I1(__252__),
    .I0(__240__),
    .O(__259__)
  );
  LUT6 #(
    .INIT(64'h69966996ffff6996)
  ) __771__ (
    .I5(__259__),
    .I4(__248__),
    .I3(__49__),
    .I2(__133__),
    .I1(__134__),
    .I0(__135__),
    .O(__260__)
  );
  LUT6 #(
    .INIT(64'h0000000000008000)
  ) __772__ (
    .I5(__125__),
    .I4(__120__),
    .I3(__219__),
    .I2(__119__),
    .I1(__121__),
    .I0(__122__),
    .O(__261__)
  );
  LUT6 #(
    .INIT(64'hfffbfeffffffffff)
  ) __773__ (
    .I5(__118__),
    .I4(__117__),
    .I3(__146__),
    .I2(__115__),
    .I1(__219__),
    .I0(__116__),
    .O(__262__)
  );
  LUT6 #(
    .INIT(64'h000000000001ffff)
  ) __774__ (
    .I5(__262__),
    .I4(__103__),
    .I3(__106__),
    .I2(__104__),
    .I1(__105__),
    .I0(__108__),
    .O(__263__)
  );
  LUT6 #(
    .INIT(64'h0000000000004000)
  ) __775__ (
    .I5(__119__),
    .I4(__120__),
    .I3(__219__),
    .I2(__121__),
    .I1(__217__),
    .I0(__107__),
    .O(__264__)
  );
  LUT5 #(
    .INIT(32'h00000004)
  ) __776__ (
    .I4(__125__),
    .I3(__121__),
    .I2(__120__),
    .I1(__119__),
    .I0(__122__),
    .O(__265__)
  );
  LUT5 #(
    .INIT(32'h00088888)
  ) __777__ (
    .I4(__176__),
    .I3(__178__),
    .I2(__57__),
    .I1(__265__),
    .I0(__107__),
    .O(__266__)
  );
  LUT4 #(
    .INIT(16'he000)
  ) __778__ (
    .I3(__176__),
    .I2(__218__),
    .I1(__178__),
    .I0(__57__),
    .O(__267__)
  );
  LUT5 #(
    .INIT(32'h000000e0)
  ) __779__ (
    .I4(__111__),
    .I3(__112__),
    .I2(__176__),
    .I1(__178__),
    .I0(__57__),
    .O(__268__)
  );
  LUT5 #(
    .INIT(32'h00004000)
  ) __780__ (
    .I4(__120__),
    .I3(__125__),
    .I2(__119__),
    .I1(__121__),
    .I0(__122__),
    .O(__269__)
  );
  LUT6 #(
    .INIT(64'haaaaaaa8a8a8aaa8)
  ) __781__ (
    .I5(__269__),
    .I4(__268__),
    .I3(__267__),
    .I2(__266__),
    .I1(__264__),
    .I0(__263__),
    .O(__270__)
  );
  LUT5 #(
    .INIT(32'h00000040)
  ) __782__ (
    .I4(__118__),
    .I3(__146__),
    .I2(__117__),
    .I1(__116__),
    .I0(__115__),
    .O(__271__)
  );
  LUT6 #(
    .INIT(64'h4000000000000000)
  ) __783__ (
    .I5(__125__),
    .I4(__119__),
    .I3(__121__),
    .I2(__120__),
    .I1(__271__),
    .I0(__122__),
    .O(__272__)
  );
  LUT5 #(
    .INIT(32'hff00fe01)
  ) __784__ (
    .I4(__125__),
    .I3(__119__),
    .I2(__121__),
    .I1(__120__),
    .I0(__122__),
    .O(__273__)
  );
  LUT6 #(
    .INIT(64'h0000000000008000)
  ) __785__ (
    .I5(__119__),
    .I4(__120__),
    .I3(__219__),
    .I2(__125__),
    .I1(__121__),
    .I0(__122__),
    .O(__274__)
  );
  LUT6 #(
    .INIT(64'h0d00000005000000)
  ) __786__ (
    .I5(__57__),
    .I4(__93__),
    .I3(__87__),
    .I2(__223__),
    .I1(__109__),
    .I0(__59__),
    .O(__275__)
  );
  LUT6 #(
    .INIT(64'h020700000a0f0000)
  ) __787__ (
    .I5(__219__),
    .I4(__275__),
    .I3(__274__),
    .I2(__273__),
    .I1(__265__),
    .I0(__107__),
    .O(__276__)
  );
  LUT6 #(
    .INIT(64'ha8a8a80000000000)
  ) __788__ (
    .I5(__176__),
    .I4(__178__),
    .I3(__57__),
    .I2(__111__),
    .I1(__112__),
    .I0(__218__),
    .O(__277__)
  );
  LUT6 #(
    .INIT(64'h000000000000e000)
  ) __789__ (
    .I5(__111__),
    .I4(__112__),
    .I3(__176__),
    .I2(__269__),
    .I1(__178__),
    .I0(__57__),
    .O(__278__)
  );
  LUT5 #(
    .INIT(32'h00f4ff0b)
  ) __790__ (
    .I4(__82__),
    .I3(__120__),
    .I2(__121__),
    .I1(__125__),
    .I0(__122__),
    .O(__279__)
  );
  LUT6 #(
    .INIT(64'hfffeffffffffffff)
  ) __791__ (
    .I5(__275__),
    .I4(__279__),
    .I3(__278__),
    .I2(__277__),
    .I1(__266__),
    .I0(__264__),
    .O(__280__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __792__ (
    .I1(__121__),
    .I0(__120__),
    .O(__281__)
  );
  LUT6 #(
    .INIT(64'h0000000000000004)
  ) __793__ (
    .I5(__278__),
    .I4(__277__),
    .I3(__266__),
    .I2(__264__),
    .I1(__275__),
    .I0(__281__),
    .O(__282__)
  );
  LUT4 #(
    .INIT(16'h02a8)
  ) __794__ (
    .I3(__105__),
    .I2(__106__),
    .I1(__104__),
    .I0(__275__),
    .O(__283__)
  );
  LUT6 #(
    .INIT(64'h0000000000008000)
  ) __795__ (
    .I5(__121__),
    .I4(__120__),
    .I3(__125__),
    .I2(__119__),
    .I1(__122__),
    .I0(__271__),
    .O(__284__)
  );
  LUT4 #(
    .INIT(16'hf888)
  ) __796__ (
    .I3(__238__),
    .I2(n3076gat),
    .I1(__236__),
    .I0(n3067gat),
    .O(__285__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __797__ (
    .I5(__242__),
    .I4(__199__),
    .I3(__249__),
    .I2(__170__),
    .I1(__240__),
    .I0(__163__),
    .O(__286__)
  );
  LUT5 #(
    .INIT(32'h000000e0)
  ) __798__ (
    .I4(n3083gat),
    .I3(n3084gat),
    .I2(n3093gat),
    .I1(n3086gat),
    .I0(n3085gat),
    .O(__287__)
  );
  LUT6 #(
    .INIT(64'h55ff54fc55ff55ff)
  ) __799__ (
    .I5(n3095gat),
    .I4(n3085gat),
    .I3(n3088gat),
    .I2(n3083gat),
    .I1(n3084gat),
    .I0(__287__),
    .O(__288__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __800__ (
    .I1(__240__),
    .I0(__110__),
    .O(__289__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __801__ (
    .I1(__243__),
    .I0(__199__),
    .O(__290__)
  );
  LUT4 #(
    .INIT(16'hb0bb)
  ) __802__ (
    .I3(__242__),
    .I2(__164__),
    .I1(__249__),
    .I0(__58__),
    .O(__291__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __803__ (
    .I1(n3085gat),
    .I0(n3083gat),
    .O(__292__)
  );
  LUT6 #(
    .INIT(64'h4000000000000000)
  ) __804__ (
    .I5(n3095gat),
    .I4(n3086gat),
    .I3(n3087gat),
    .I2(n3088gat),
    .I1(__292__),
    .I0(n3084gat),
    .O(__293__)
  );
  LUT3 #(
    .INIT(8'h0b)
  ) __805__ (
    .I2(__293__),
    .I1(__287__),
    .I0(n3088gat),
    .O(__294__)
  );
  LUT6 #(
    .INIT(64'h11111111fff1ffff)
  ) __806__ (
    .I5(__294__),
    .I4(__291__),
    .I3(__290__),
    .I2(__289__),
    .I1(__288__),
    .I0(__286__),
    .O(__295__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __807__ (
    .I1(__97__),
    .I0(n3084gat),
    .O(__296__)
  );
  LUT6 #(
    .INIT(64'h0000000000008000)
  ) __808__ (
    .I5(n3086gat),
    .I4(__237__),
    .I3(n3095gat),
    .I2(n3087gat),
    .I1(__292__),
    .I0(__296__),
    .O(__297__)
  );
  LUT6 #(
    .INIT(64'h0000000000004000)
  ) __809__ (
    .I5(n3087gat),
    .I4(n3083gat),
    .I3(n3093gat),
    .I2(n3088gat),
    .I1(__97__),
    .I0(n3084gat),
    .O(__298__)
  );
  LUT6 #(
    .INIT(64'hafffefffafffafff)
  ) __810__ (
    .I5(n3086gat),
    .I4(n3085gat),
    .I3(__121__),
    .I2(__120__),
    .I1(__298__),
    .I0(__297__),
    .O(__299__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __811__ (
    .I1(__57__),
    .I0(__109__),
    .O(__300__)
  );
  LUT6 #(
    .INIT(64'h0d00000000000000)
  ) __812__ (
    .I5(__262__),
    .I4(__93__),
    .I3(__87__),
    .I2(__223__),
    .I1(__300__),
    .I0(__59__),
    .O(__301__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __813__ (
    .I1(__242__),
    .I0(__249__),
    .O(__302__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __814__ (
    .I1(__240__),
    .I0(__166__),
    .O(__303__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __815__ (
    .I1(__240__),
    .I0(__150__),
    .O(__304__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __816__ (
    .I1(__249__),
    .I0(__141__),
    .O(__305__)
  );
  LUT6 #(
    .INIT(64'h000000000000b0bb)
  ) __817__ (
    .I5(__305__),
    .I4(__304__),
    .I3(__243__),
    .I2(__205__),
    .I1(__242__),
    .I0(__169__),
    .O(__306__)
  );
  LUT6 #(
    .INIT(64'h000000fff1f1f1ff)
  ) __818__ (
    .I5(__288__),
    .I4(__294__),
    .I3(__306__),
    .I2(__303__),
    .I1(__205__),
    .I0(__302__),
    .O(__307__)
  );
  LUT6 #(
    .INIT(64'haaffffccf0ffffff)
  ) __819__ (
    .I5(__191__),
    .I4(__187__),
    .I3(__193__),
    .I2(__203__),
    .I1(__199__),
    .I0(__169__),
    .O(__308__)
  );
  LUT6 #(
    .INIT(64'hffaaffccf0ffffff)
  ) __820__ (
    .I5(__193__),
    .I4(__191__),
    .I3(__187__),
    .I2(__202__),
    .I1(__201__),
    .I0(__155__),
    .O(__309__)
  );
  LUT5 #(
    .INIT(32'hfcfaffff)
  ) __821__ (
    .I4(__193__),
    .I3(__187__),
    .I2(__191__),
    .I1(__53__),
    .I0(__180__),
    .O(__310__)
  );
  LUT3 #(
    .INIT(8'h40)
  ) __822__ (
    .I2(__191__),
    .I1(__193__),
    .I0(__187__),
    .O(__311__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __823__ (
    .I2(__187__),
    .I1(__191__),
    .I0(__193__),
    .O(__312__)
  );
  LUT5 #(
    .INIT(32'hfcfaffff)
  ) __824__ (
    .I4(__191__),
    .I3(__187__),
    .I2(__193__),
    .I1(__50__),
    .I0(__170__),
    .O(__313__)
  );
  LUT5 #(
    .INIT(32'hbb0b0000)
  ) __825__ (
    .I4(__313__),
    .I3(__141__),
    .I2(__312__),
    .I1(__311__),
    .I0(__52__),
    .O(__314__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __826__ (
    .I1(__184__),
    .I0(__190__),
    .O(__315__)
  );
  LUT6 #(
    .INIT(64'h777700000fff0000)
  ) __827__ (
    .I5(__220__),
    .I4(__315__),
    .I3(__314__),
    .I2(__310__),
    .I1(__309__),
    .I0(__308__),
    .O(__316__)
  );
  LUT5 #(
    .INIT(32'h00004000)
  ) __828__ (
    .I4(__149__),
    .I3(__206__),
    .I2(__205__),
    .I1(__47__),
    .I0(__90__),
    .O(__317__)
  );
  LUT5 #(
    .INIT(32'hb0000000)
  ) __829__ (
    .I4(__187__),
    .I3(__191__),
    .I2(__193__),
    .I1(__130__),
    .I0(__317__),
    .O(__318__)
  );
  LUT6 #(
    .INIT(64'h0003000500000000)
  ) __830__ (
    .I5(__187__),
    .I4(__220__),
    .I3(__191__),
    .I2(__193__),
    .I1(__159__),
    .I0(__197__),
    .O(__319__)
  );
  LUT6 #(
    .INIT(64'h0000000300000005)
  ) __831__ (
    .I5(__220__),
    .I4(__187__),
    .I3(__191__),
    .I2(__193__),
    .I1(__161__),
    .I0(__56__),
    .O(__320__)
  );
  LUT6 #(
    .INIT(64'h0008080000000800)
  ) __832__ (
    .I5(__206__),
    .I4(__205__),
    .I3(__149__),
    .I2(__90__),
    .I1(__47__),
    .I0(__311__),
    .O(__321__)
  );
  LUT6 #(
    .INIT(64'hffffffaaccf0ffff)
  ) __833__ (
    .I5(__191__),
    .I4(__193__),
    .I3(__187__),
    .I2(__127__),
    .I1(__142__),
    .I0(__58__),
    .O(__322__)
  );
  LUT6 #(
    .INIT(64'hffffffaaccf0ffff)
  ) __834__ (
    .I5(__191__),
    .I4(__193__),
    .I3(__187__),
    .I2(__175__),
    .I1(__181__),
    .I0(__164__),
    .O(__323__)
  );
  LUT3 #(
    .INIT(8'h40)
  ) __835__ (
    .I2(__187__),
    .I1(__191__),
    .I0(__193__),
    .O(__324__)
  );
  LUT6 #(
    .INIT(64'h33ff00ff5f5f0f0f)
  ) __836__ (
    .I5(__220__),
    .I4(__324__),
    .I3(__323__),
    .I2(__322__),
    .I1(__179__),
    .I0(__138__),
    .O(__325__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __837__ (
    .I1(__184__),
    .I0(__190__),
    .O(__326__)
  );
  LUT6 #(
    .INIT(64'hfffffffe00000000)
  ) __838__ (
    .I5(__326__),
    .I4(__325__),
    .I3(__321__),
    .I2(__320__),
    .I1(__319__),
    .I0(__318__),
    .O(__327__)
  );
  LUT5 #(
    .INIT(32'hfcfaffff)
  ) __839__ (
    .I4(__187__),
    .I3(__193__),
    .I2(__191__),
    .I1(__152__),
    .I0(__150__),
    .O(__328__)
  );
  LUT6 #(
    .INIT(64'hf0c0f0f0f0f0f0a0)
  ) __840__ (
    .I5(__187__),
    .I4(__191__),
    .I3(__193__),
    .I2(__328__),
    .I1(__140__),
    .I0(__148__),
    .O(__329__)
  );
  LUT5 #(
    .INIT(32'hcffaffff)
  ) __841__ (
    .I4(__193__),
    .I3(__187__),
    .I2(__191__),
    .I1(__154__),
    .I0(__110__),
    .O(__330__)
  );
  LUT6 #(
    .INIT(64'hf0c0f0a0f0f0f0f0)
  ) __842__ (
    .I5(__191__),
    .I4(__193__),
    .I3(__187__),
    .I2(__330__),
    .I1(__151__),
    .I0(__139__),
    .O(__331__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __843__ (
    .I1(__184__),
    .I0(__190__),
    .O(__332__)
  );
  LUT6 #(
    .INIT(64'h6900000096000000)
  ) __844__ (
    .I5(__154__),
    .I4(__332__),
    .I3(__312__),
    .I2(__151__),
    .I1(__251__),
    .I0(__206__),
    .O(__333__)
  );
  LUT4 #(
    .INIT(16'hefff)
  ) __845__ (
    .I3(__149__),
    .I2(__47__),
    .I1(__205__),
    .I0(__90__),
    .O(__334__)
  );
  LUT6 #(
    .INIT(64'h00000000f0f7f0f0)
  ) __846__ (
    .I5(__334__),
    .I4(__190__),
    .I3(__184__),
    .I2(__333__),
    .I1(__331__),
    .I0(__329__),
    .O(__335__)
  );
  LUT6 #(
    .INIT(64'h9669699669969669)
  ) __847__ (
    .I5(__184__),
    .I4(__187__),
    .I3(__191__),
    .I2(__193__),
    .I1(__190__),
    .I0(__123__),
    .O(__336__)
  );
  LUT3 #(
    .INIT(8'h04)
  ) __848__ (
    .I2(__155__),
    .I1(__97__),
    .I0(__94__),
    .O(__337__)
  );
  LUT6 #(
    .INIT(64'h0f0c0f0a0f0f0f0f)
  ) __849__ (
    .I5(__220__),
    .I4(__219__),
    .I3(__113__),
    .I2(__337__),
    .I1(__96__),
    .I0(__95__),
    .O(__338__)
  );
  LUT6 #(
    .INIT(64'hffe0ffffffffffff)
  ) __850__ (
    .I5(__338__),
    .I4(__336__),
    .I3(__335__),
    .I2(__114__),
    .I1(__327__),
    .I0(__316__),
    .O(__339__)
  );
  LUT3 #(
    .INIT(8'h96)
  ) __851__ (
    .I2(__149__),
    .I1(__47__),
    .I0(__170__),
    .O(__340__)
  );
  LUT6 #(
    .INIT(64'h9669699669969669)
  ) __852__ (
    .I5(__174__),
    .I4(__245__),
    .I3(__180__),
    .I2(__50__),
    .I1(__53__),
    .I0(__340__),
    .O(__341__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __853__ (
    .I1(__249__),
    .I0(__56__),
    .O(__342__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __854__ (
    .I1(__242__),
    .I0(__161__),
    .O(__343__)
  );
  LUT6 #(
    .INIT(64'h000000000000b0bb)
  ) __855__ (
    .I5(__343__),
    .I4(__342__),
    .I3(__243__),
    .I2(__47__),
    .I1(__240__),
    .I0(__139__),
    .O(__344__)
  );
  LUT6 #(
    .INIT(64'h5555555755555555)
  ) __856__ (
    .I5(n3095gat),
    .I4(n3085gat),
    .I3(n3083gat),
    .I2(n3084gat),
    .I1(__344__),
    .I0(__341__),
    .O(__345__)
  );
  LUT4 #(
    .INIT(16'h9669)
  ) __857__ (
    .I3(__49__),
    .I2(__133__),
    .I1(__134__),
    .I0(__135__),
    .O(__346__)
  );
  LUT6 #(
    .INIT(64'hdc7373dc73dcdc73)
  ) __858__ (
    .I5(__154__),
    .I4(__151__),
    .I3(__251__),
    .I2(__248__),
    .I1(__156__),
    .I0(__306__),
    .O(__347__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __859__ (
    .I5(__242__),
    .I4(__202__),
    .I3(__249__),
    .I2(__50__),
    .I1(__240__),
    .I0(__171__),
    .O(__348__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __860__ (
    .I1(__243__),
    .I0(__202__),
    .O(__349__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __861__ (
    .I1(__249__),
    .I0(__138__),
    .O(__350__)
  );
  LUT4 #(
    .INIT(16'hb0bb)
  ) __862__ (
    .I3(__242__),
    .I2(__179__),
    .I1(__240__),
    .I0(__152__),
    .O(__351__)
  );
  LUT6 #(
    .INIT(64'h11111111fff1ffff)
  ) __863__ (
    .I5(__294__),
    .I4(__351__),
    .I3(__350__),
    .I2(__349__),
    .I1(__288__),
    .I0(__348__),
    .O(__352__)
  );
  LUT4 #(
    .INIT(16'hb4ff)
  ) __864__ (
    .I3(__275__),
    .I2(__143__),
    .I1(__106__),
    .I0(__104__),
    .O(__353__)
  );
  LUT6 #(
    .INIT(64'h0000000000000040)
  ) __865__ (
    .I5(__206__),
    .I4(__90__),
    .I3(__47__),
    .I2(__205__),
    .I1(__149__),
    .I0(__81__),
    .O(__354__)
  );
  LUT4 #(
    .INIT(16'h00e0)
  ) __866__ (
    .I3(n3086gat),
    .I2(n3085gat),
    .I1(n3092gat),
    .I0(n3091gat),
    .O(__355__)
  );
  LUT5 #(
    .INIT(32'h00007fff)
  ) __867__ (
    .I4(__238__),
    .I3(n3087gat),
    .I2(n3088gat),
    .I1(__235__),
    .I0(__355__),
    .O(__356__)
  );
  LUT6 #(
    .INIT(64'h0300fcffaaaaaaaa)
  ) __868__ (
    .I5(__356__),
    .I4(__73__),
    .I3(__354__),
    .I2(__75__),
    .I1(__61__),
    .I0(n3065gat),
    .O(__357__)
  );
  LUT6 #(
    .INIT(64'h0003000500000000)
  ) __869__ (
    .I5(__275__),
    .I4(__268__),
    .I3(__266__),
    .I2(__264__),
    .I1(__269__),
    .I0(__267__),
    .O(__358__)
  );
  LUT5 #(
    .INIT(32'h333c777d)
  ) __870__ (
    .I4(__90__),
    .I3(__121__),
    .I2(__120__),
    .I1(__122__),
    .I0(__201__),
    .O(__359__)
  );
  LUT3 #(
    .INIT(8'h40)
  ) __871__ (
    .I2(__119__),
    .I1(__121__),
    .I0(__120__),
    .O(__360__)
  );
  LUT6 #(
    .INIT(64'h8000000000000000)
  ) __872__ (
    .I5(__118__),
    .I4(__115__),
    .I3(__125__),
    .I2(__122__),
    .I1(__360__),
    .I0(__215__),
    .O(__361__)
  );
  LUT4 #(
    .INIT(16'hf888)
  ) __873__ (
    .I3(n3093gat),
    .I2(n3066gat),
    .I1(n3095gat),
    .I0(n3075gat),
    .O(__362__)
  );
  LUT6 #(
    .INIT(64'h8000000000000000)
  ) __874__ (
    .I5(__93__),
    .I4(__87__),
    .I3(__91__),
    .I2(__55__),
    .I1(__144__),
    .I0(__92__),
    .O(__363__)
  );
  LUT5 #(
    .INIT(32'h2aaaaaaa)
  ) __875__ (
    .I4(__97__),
    .I3(__60__),
    .I2(__147__),
    .I1(__98__),
    .I0(__363__),
    .O(__364__)
  );
  LUT6 #(
    .INIT(64'h0000000000004000)
  ) __876__ (
    .I5(__79__),
    .I4(__90__),
    .I3(__206__),
    .I2(__205__),
    .I1(__149__),
    .I0(__47__),
    .O(__365__)
  );
  LUT6 #(
    .INIT(64'heeeeaaaaccccf00f)
  ) __877__ (
    .I5(__238__),
    .I4(__236__),
    .I3(__365__),
    .I2(__80__),
    .I1(n3071gat),
    .I0(n3080gat),
    .O(__366__)
  );
  LUT6 #(
    .INIT(64'heffffffbffffffff)
  ) __878__ (
    .I5(__185__),
    .I4(__173__),
    .I3(__182__),
    .I2(__177__),
    .I1(__183__),
    .I0(__186__),
    .O(__367__)
  );
  LUT6 #(
    .INIT(64'h000000000000fbbf)
  ) __879__ (
    .I5(__184__),
    .I4(__367__),
    .I3(__187__),
    .I2(__191__),
    .I1(__193__),
    .I0(__190__),
    .O(__368__)
  );
  LUT6 #(
    .INIT(64'h020800000a000000)
  ) __880__ (
    .I5(__206__),
    .I4(__205__),
    .I3(__149__),
    .I2(__90__),
    .I1(__47__),
    .I0(__368__),
    .O(__369__)
  );
  LUT5 #(
    .INIT(32'hfefcfaf0)
  ) __881__ (
    .I4(n3093gat),
    .I3(n3095gat),
    .I2(__369__),
    .I1(n3073gat),
    .I0(n3082gat),
    .O(__370__)
  );
  LUT4 #(
    .INIT(16'h56ff)
  ) __882__ (
    .I3(__162__),
    .I2(__106__),
    .I1(__104__),
    .I0(__105__),
    .O(__371__)
  );
  LUT5 #(
    .INIT(32'h00000004)
  ) __883__ (
    .I4(__206__),
    .I3(__205__),
    .I2(__90__),
    .I1(__149__),
    .I0(__47__),
    .O(__372__)
  );
  LUT6 #(
    .INIT(64'h0000000000004000)
  ) __884__ (
    .I5(n3085gat),
    .I4(n3083gat),
    .I3(n3095gat),
    .I2(n3086gat),
    .I1(__97__),
    .I0(n3084gat),
    .O(__373__)
  );
  LUT6 #(
    .INIT(64'h0000000000004000)
  ) __885__ (
    .I5(n3085gat),
    .I4(n3083gat),
    .I3(n3095gat),
    .I2(n3087gat),
    .I1(__97__),
    .I0(n3084gat),
    .O(__374__)
  );
  LUT4 #(
    .INIT(16'he000)
  ) __886__ (
    .I3(n3086gat),
    .I2(n3085gat),
    .I1(n3092gat),
    .I0(n3091gat),
    .O(__375__)
  );
  LUT6 #(
    .INIT(64'h0000bfffbfffbfff)
  ) __887__ (
    .I5(__375__),
    .I4(__298__),
    .I3(n3094gat),
    .I2(__374__),
    .I1(__373__),
    .I0(__237__),
    .O(__376__)
  );
  LUT3 #(
    .INIT(8'hf4)
  ) __888__ (
    .I2(__369__),
    .I1(n3072gat),
    .I0(__376__),
    .O(__377__)
  );
  LUT6 #(
    .INIT(64'hfeeefcccfaaaf000)
  ) __889__ (
    .I5(n3093gat),
    .I4(n3095gat),
    .I3(__229__),
    .I2(__368__),
    .I1(n3070gat),
    .I0(n3079gat),
    .O(__378__)
  );
  LUT6 #(
    .INIT(64'h2222222222222228)
  ) __890__ (
    .I5(__118__),
    .I4(__117__),
    .I3(__146__),
    .I2(__115__),
    .I1(__116__),
    .I0(__301__),
    .O(__379__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __891__ (
    .I1(__240__),
    .I0(__48__),
    .O(__380__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __892__ (
    .I1(__243__),
    .I0(__149__),
    .O(__381__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __893__ (
    .I1(__249__),
    .I0(__197__),
    .O(__382__)
  );
  LUT6 #(
    .INIT(64'h000000000000b0bb)
  ) __894__ (
    .I5(__382__),
    .I4(__381__),
    .I3(__242__),
    .I2(__159__),
    .I1(__240__),
    .I0(__140__),
    .O(__383__)
  );
  LUT6 #(
    .INIT(64'h000000fff1f1f1ff)
  ) __895__ (
    .I5(__288__),
    .I4(__294__),
    .I3(__383__),
    .I2(__380__),
    .I1(__149__),
    .I0(__302__),
    .O(__384__)
  );
  LUT4 #(
    .INIT(16'hf888)
  ) __896__ (
    .I3(__238__),
    .I2(n3075gat),
    .I1(__236__),
    .I0(n3066gat),
    .O(__385__)
  );
  LUT3 #(
    .INIT(8'hf4)
  ) __897__ (
    .I2(__369__),
    .I1(n3067gat),
    .I0(__376__),
    .O(__386__)
  );
  LUT4 #(
    .INIT(16'hb000)
  ) __898__ (
    .I3(n3100gat),
    .I2(__196__),
    .I1(__192__),
    .I0(__188__),
    .O(__387__)
  );
  LUT6 #(
    .INIT(64'h0000000000004000)
  ) __899__ (
    .I5(__205__),
    .I4(__90__),
    .I3(__206__),
    .I2(__149__),
    .I1(__387__),
    .I0(__47__),
    .O(__388__)
  );
  LUT3 #(
    .INIT(8'hf4)
  ) __900__ (
    .I2(__369__),
    .I1(n3071gat),
    .I0(__376__),
    .O(__389__)
  );
  LUT4 #(
    .INIT(16'h6996)
  ) __901__ (
    .I3(__154__),
    .I2(__151__),
    .I1(__251__),
    .I0(__156__),
    .O(__390__)
  );
  LUT6 #(
    .INIT(64'hfeeefcccfaaaf000)
  ) __902__ (
    .I5(n3093gat),
    .I4(n3095gat),
    .I3(__229__),
    .I2(__368__),
    .I1(n3069gat),
    .I0(n3078gat),
    .O(__391__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __903__ (
    .I1(__90__),
    .I0(__203__),
    .O(__392__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __904__ (
    .I1(__240__),
    .I0(__162__),
    .O(__393__)
  );
  LUT6 #(
    .INIT(64'h000000fff1f1f1ff)
  ) __905__ (
    .I5(__288__),
    .I4(__294__),
    .I3(__344__),
    .I2(__393__),
    .I1(__47__),
    .I0(__302__),
    .O(__394__)
  );
  LUT6 #(
    .INIT(64'hfeeefcccfaaaf000)
  ) __906__ (
    .I5(n3072gat),
    .I4(n3095gat),
    .I3(__229__),
    .I2(__368__),
    .I1(n3093gat),
    .I0(n3081gat),
    .O(__395__)
  );
  LUT5 #(
    .INIT(32'h0000e000)
  ) __907__ (
    .I4(__113__),
    .I3(__176__),
    .I2(__229__),
    .I1(__178__),
    .I0(__57__),
    .O(__396__)
  );
  LUT5 #(
    .INIT(32'h00000040)
  ) __908__ (
    .I4(__184__),
    .I3(__191__),
    .I2(__187__),
    .I1(__193__),
    .I0(__190__),
    .O(__397__)
  );
  LUT5 #(
    .INIT(32'h12203020)
  ) __909__ (
    .I4(__206__),
    .I3(__205__),
    .I2(__149__),
    .I1(__90__),
    .I0(__47__),
    .O(__398__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __910__ (
    .I1(__113__),
    .I0(__66__),
    .O(__399__)
  );
  LUT6 #(
    .INIT(64'h00efefefffffffff)
  ) __911__ (
    .I5(__219__),
    .I4(__220__),
    .I3(__399__),
    .I2(__398__),
    .I1(__64__),
    .I0(__397__),
    .O(__400__)
  );
  LUT6 #(
    .INIT(64'h0000f0f0000000bb)
  ) __912__ (
    .I5(__219__),
    .I4(__95__),
    .I3(__65__),
    .I2(__66__),
    .I1(__334__),
    .I0(__113__),
    .O(__401__)
  );
  LUT5 #(
    .INIT(32'h0000e000)
  ) __913__ (
    .I4(__62__),
    .I3(__176__),
    .I2(__65__),
    .I1(__178__),
    .I0(__57__),
    .O(__402__)
  );
  LUT3 #(
    .INIT(8'h04)
  ) __914__ (
    .I2(__98__),
    .I1(__97__),
    .I0(n3098gat),
    .O(__403__)
  );
  LUT6 #(
    .INIT(64'h00007f000000ffff)
  ) __915__ (
    .I5(__403__),
    .I4(__402__),
    .I3(__192__),
    .I2(__300__),
    .I1(__188__),
    .I0(n3097gat),
    .O(__404__)
  );
  LUT6 #(
    .INIT(64'hffff444fffffffff)
  ) __916__ (
    .I5(__404__),
    .I4(__401__),
    .I3(__96__),
    .I2(__400__),
    .I1(__396__),
    .I0(__67__),
    .O(__405__)
  );
  LUT3 #(
    .INIT(8'h70)
  ) __917__ (
    .I2(__275__),
    .I1(__106__),
    .I0(__104__),
    .O(__406__)
  );
  LUT3 #(
    .INIT(8'hf4)
  ) __918__ (
    .I2(__369__),
    .I1(n3065gat),
    .I0(__376__),
    .O(__407__)
  );
  LUT4 #(
    .INIT(16'h56ff)
  ) __919__ (
    .I3(__171__),
    .I2(__117__),
    .I1(__146__),
    .I0(__118__),
    .O(__408__)
  );
  LUT4 #(
    .INIT(16'hf888)
  ) __920__ (
    .I3(n3093gat),
    .I2(n3069gat),
    .I1(n3095gat),
    .I0(n3078gat),
    .O(__409__)
  );
  LUT6 #(
    .INIT(64'h55555556ffffffff)
  ) __921__ (
    .I5(__172__),
    .I4(__118__),
    .I3(__117__),
    .I2(__146__),
    .I1(__115__),
    .I0(__116__),
    .O(__410__)
  );
  LUT3 #(
    .INIT(8'h07)
  ) __922__ (
    .I2(__222__),
    .I1(__57__),
    .I0(__109__),
    .O(__411__)
  );
  LUT4 #(
    .INIT(16'hf888)
  ) __923__ (
    .I3(n3068gat),
    .I2(__236__),
    .I1(n3077gat),
    .I0(__238__),
    .O(__412__)
  );
  LUT5 #(
    .INIT(32'h0bfff400)
  ) __924__ (
    .I4(__78__),
    .I3(__232__),
    .I2(__79__),
    .I1(__77__),
    .I0(__80__),
    .O(__413__)
  );
  LUT5 #(
    .INIT(32'hfcccf055)
  ) __925__ (
    .I4(__238__),
    .I3(__236__),
    .I2(n3073gat),
    .I1(n3082gat),
    .I0(__413__),
    .O(__414__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __926__ (
    .I5(__242__),
    .I4(__203__),
    .I3(__249__),
    .I2(__53__),
    .I1(__240__),
    .I0(__172__),
    .O(__415__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __927__ (
    .I1(__249__),
    .I0(__142__),
    .O(__416__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __928__ (
    .I1(__240__),
    .I0(__154__),
    .O(__417__)
  );
  LUT4 #(
    .INIT(16'hb0bb)
  ) __929__ (
    .I3(__243__),
    .I2(__203__),
    .I1(__242__),
    .I0(__181__),
    .O(__418__)
  );
  LUT6 #(
    .INIT(64'h11111111fff1ffff)
  ) __930__ (
    .I5(__294__),
    .I4(__418__),
    .I3(__417__),
    .I2(__416__),
    .I1(__288__),
    .I0(__415__),
    .O(__419__)
  );
  LUT3 #(
    .INIT(8'h7f)
  ) __931__ (
    .I2(__166__),
    .I1(__106__),
    .I0(__104__),
    .O(__420__)
  );
  LUT3 #(
    .INIT(8'h01)
  ) __932__ (
    .I2(__98__),
    .I1(__89__),
    .I0(__102__),
    .O(__421__)
  );
  LUT6 #(
    .INIT(64'h0000003100003131)
  ) __933__ (
    .I5(__57__),
    .I4(__223__),
    .I3(__109__),
    .I2(__99__),
    .I1(__222__),
    .I0(__98__),
    .O(__422__)
  );
  LUT6 #(
    .INIT(64'hfeeefcccfaaaf000)
  ) __934__ (
    .I5(n3093gat),
    .I4(n3095gat),
    .I3(__229__),
    .I2(__368__),
    .I1(n3067gat),
    .I0(n3076gat),
    .O(__423__)
  );
  LUT6 #(
    .INIT(64'h4040ff0000000000)
  ) __935__ (
    .I5(__271__),
    .I4(__219__),
    .I3(__218__),
    .I2(__217__),
    .I1(__216__),
    .I0(__119__),
    .O(__424__)
  );
  LUT5 #(
    .INIT(32'hfefcfaf0)
  ) __936__ (
    .I4(n3093gat),
    .I3(n3095gat),
    .I2(__369__),
    .I1(n3065gat),
    .I0(n3074gat),
    .O(__425__)
  );
  LUT6 #(
    .INIT(64'h0000000000000040)
  ) __937__ (
    .I5(__121__),
    .I4(__120__),
    .I3(__122__),
    .I2(__125__),
    .I1(__119__),
    .I0(__222__),
    .O(__426__)
  );
  LUT6 #(
    .INIT(64'h4000000000000000)
  ) __938__ (
    .I5(n3095gat),
    .I4(n3086gat),
    .I3(__292__),
    .I2(n3094gat),
    .I1(__97__),
    .I0(n3084gat),
    .O(__427__)
  );
  LUT4 #(
    .INIT(16'h01fe)
  ) __939__ (
    .I3(__125__),
    .I2(__121__),
    .I1(__120__),
    .I0(__122__),
    .O(__428__)
  );
  LUT6 #(
    .INIT(64'hffffffffff101010)
  ) __940__ (
    .I5(__428__),
    .I4(__355__),
    .I3(__298__),
    .I2(__427__),
    .I1(__237__),
    .I0(__374__),
    .O(__429__)
  );
  LUT5 #(
    .INIT(32'h00000040)
  ) __941__ (
    .I4(__118__),
    .I3(__117__),
    .I2(__146__),
    .I1(__116__),
    .I0(__115__),
    .O(__430__)
  );
  LUT6 #(
    .INIT(64'h0000000000000040)
  ) __942__ (
    .I5(__125__),
    .I4(__121__),
    .I3(__120__),
    .I2(__119__),
    .I1(__430__),
    .I0(__122__),
    .O(__431__)
  );
  LUT6 #(
    .INIT(64'hbfff0f0fbfbf0f0f)
  ) __943__ (
    .I5(__243__),
    .I4(__248__),
    .I3(__199__),
    .I2(__247__),
    .I1(__291__),
    .I0(__289__),
    .O(__432__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __944__ (
    .I1(n3083gat),
    .I0(n3084gat),
    .O(__433__)
  );
  LUT6 #(
    .INIT(64'h9669699669969669)
  ) __945__ (
    .I5(n3086gat),
    .I4(n3087gat),
    .I3(n3085gat),
    .I2(n3088gat),
    .I1(n3089gat),
    .I0(__433__),
    .O(__434__)
  );
  LUT6 #(
    .INIT(64'hbfff0f0fbfbf0f0f)
  ) __946__ (
    .I5(__249__),
    .I4(__248__),
    .I3(__142__),
    .I2(__434__),
    .I1(__418__),
    .I0(__417__),
    .O(__435__)
  );
  LUT5 #(
    .INIT(32'h00000040)
  ) __947__ (
    .I4(__206__),
    .I3(__90__),
    .I2(__205__),
    .I1(__149__),
    .I0(__47__),
    .O(__436__)
  );
  LUT4 #(
    .INIT(16'hc3aa)
  ) __948__ (
    .I3(__356__),
    .I2(__436__),
    .I1(__81__),
    .I0(n3068gat),
    .O(__437__)
  );
  LUT3 #(
    .INIT(8'h40)
  ) __949__ (
    .I2(n3086gat),
    .I1(__298__),
    .I0(n3085gat),
    .O(__438__)
  );
  LUT6 #(
    .INIT(64'hefefefcfafafaf0f)
  ) __950__ (
    .I5(n3094gat),
    .I4(n3092gat),
    .I3(n3091gat),
    .I2(__273__),
    .I1(__297__),
    .I0(__438__),
    .O(__439__)
  );
  LUT4 #(
    .INIT(16'hf888)
  ) __951__ (
    .I3(n3093gat),
    .I2(n3065gat),
    .I1(n3095gat),
    .I0(n3074gat),
    .O(__440__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __952__ (
    .I5(__243__),
    .I4(__206__),
    .I3(__249__),
    .I2(__52__),
    .I1(__240__),
    .I0(__148__),
    .O(__441__)
  );
  LUT6 #(
    .INIT(64'h6996966996696996)
  ) __953__ (
    .I5(__163__),
    .I4(__48__),
    .I3(__162__),
    .I2(__165__),
    .I1(__166__),
    .I0(__171__),
    .O(__442__)
  );
  LUT4 #(
    .INIT(16'h6996)
  ) __954__ (
    .I3(__160__),
    .I2(__172__),
    .I1(__167__),
    .I0(__442__),
    .O(__443__)
  );
  LUT6 #(
    .INIT(64'h44cc44c4ffffffff)
  ) __955__ (
    .I5(__443__),
    .I4(__256__),
    .I3(__155__),
    .I2(__242__),
    .I1(__248__),
    .I0(__441__),
    .O(__444__)
  );
  LUT3 #(
    .INIT(8'hf4)
  ) __956__ (
    .I2(__369__),
    .I1(n3068gat),
    .I0(__376__),
    .O(__445__)
  );
  LUT6 #(
    .INIT(64'h0000000000004000)
  ) __957__ (
    .I5(__118__),
    .I4(__117__),
    .I3(__146__),
    .I2(__116__),
    .I1(__218__),
    .I0(__115__),
    .O(__446__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __958__ (
    .I1(__240__),
    .I0(__165__),
    .O(__447__)
  );
  LUT4 #(
    .INIT(16'hf100)
  ) __959__ (
    .I3(__441__),
    .I2(__155__),
    .I1(__256__),
    .I0(__242__),
    .O(__448__)
  );
  LUT6 #(
    .INIT(64'h000000fff1f1f1ff)
  ) __960__ (
    .I5(__288__),
    .I4(__294__),
    .I3(__448__),
    .I2(__447__),
    .I1(__206__),
    .I0(__302__),
    .O(__449__)
  );
  LUT6 #(
    .INIT(64'hffe0ffffffffffff)
  ) __961__ (
    .I5(__338__),
    .I4(__209__),
    .I3(__335__),
    .I2(__114__),
    .I1(__327__),
    .I0(__316__),
    .O(__450__)
  );
  LUT3 #(
    .INIT(8'hf4)
  ) __962__ (
    .I2(__369__),
    .I1(n3069gat),
    .I0(__376__),
    .O(__451__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __963__ (
    .I5(__242__),
    .I4(__201__),
    .I3(__249__),
    .I2(__180__),
    .I1(__240__),
    .I0(__167__),
    .O(__452__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __964__ (
    .I1(__249__),
    .I0(__127__),
    .O(__453__)
  );
  LUT6 #(
    .INIT(64'h11111111fff1ffff)
  ) __965__ (
    .I5(__294__),
    .I4(__244__),
    .I3(__453__),
    .I2(__241__),
    .I1(__288__),
    .I0(__452__),
    .O(__454__)
  );
  LUT3 #(
    .INIT(8'hf4)
  ) __966__ (
    .I2(__369__),
    .I1(n3073gat),
    .I0(__376__),
    .O(__455__)
  );
  LUT4 #(
    .INIT(16'hf888)
  ) __967__ (
    .I3(n3093gat),
    .I2(n3071gat),
    .I1(n3095gat),
    .I0(n3080gat),
    .O(__456__)
  );
  LUT4 #(
    .INIT(16'hf888)
  ) __968__ (
    .I3(n3093gat),
    .I2(n3067gat),
    .I1(n3095gat),
    .I0(n3076gat),
    .O(__457__)
  );
  LUT6 #(
    .INIT(64'h0000000000000040)
  ) __969__ (
    .I5(__206__),
    .I4(__205__),
    .I3(__90__),
    .I2(__149__),
    .I1(__387__),
    .I0(__47__),
    .O(__458__)
  );
  LUT6 #(
    .INIT(64'h000000000d000000)
  ) __970__ (
    .I5(__90__),
    .I4(n3100gat),
    .I3(__196__),
    .I2(__203__),
    .I1(__188__),
    .I0(__192__),
    .O(__459__)
  );
  LUT5 #(
    .INIT(32'h00008000)
  ) __971__ (
    .I4(__121__),
    .I3(__125__),
    .I2(__119__),
    .I1(__120__),
    .I0(__122__),
    .O(__460__)
  );
  LUT6 #(
    .INIT(64'h0000000022222228)
  ) __972__ (
    .I5(__277__),
    .I4(__121__),
    .I3(__120__),
    .I2(__122__),
    .I1(__125__),
    .I0(__275__),
    .O(__461__)
  );
  LUT6 #(
    .INIT(64'h000000000000ff8f)
  ) __973__ (
    .I5(__219__),
    .I4(__69__),
    .I3(__220__),
    .I2(__334__),
    .I1(__229__),
    .I0(__71__),
    .O(__462__)
  );
  LUT6 #(
    .INIT(64'hffff00ffefefefef)
  ) __974__ (
    .I5(__219__),
    .I4(__70__),
    .I3(__64__),
    .I2(__229__),
    .I1(__63__),
    .I0(__113__),
    .O(__463__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __975__ (
    .I1(__463__),
    .I0(__462__),
    .O(__464__)
  );
  LUT6 #(
    .INIT(64'h00fff4ff00ff00ff)
  ) __976__ (
    .I5(__219__),
    .I4(__68__),
    .I3(__464__),
    .I2(__220__),
    .I1(__398__),
    .I0(__64__),
    .O(__465__)
  );
  LUT5 #(
    .INIT(32'h00008000)
  ) __977__ (
    .I4(__183__),
    .I3(__185__),
    .I2(__182__),
    .I1(__177__),
    .I0(__186__),
    .O(__466__)
  );
  LUT6 #(
    .INIT(64'h4000000000000000)
  ) __978__ (
    .I5(__187__),
    .I4(__191__),
    .I3(__193__),
    .I2(__190__),
    .I1(__466__),
    .I0(__184__),
    .O(__467__)
  );
  LUT3 #(
    .INIT(8'h69)
  ) __979__ (
    .I2(__172__),
    .I1(__167__),
    .I0(__442__),
    .O(__468__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __980__ (
    .I1(__51__),
    .I0(__158__),
    .O(__469__)
  );
  LUT6 #(
    .INIT(64'hbfffffffffffffff)
  ) __981__ (
    .I5(__469__),
    .I4(__194__),
    .I3(__153__),
    .I2(__157__),
    .I1(__198__),
    .I0(n3090gat),
    .O(__470__)
  );
  LUT4 #(
    .INIT(16'hf888)
  ) __982__ (
    .I3(n3093gat),
    .I2(n3070gat),
    .I1(n3095gat),
    .I0(n3079gat),
    .O(__471__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __983__ (
    .I1(__195__),
    .I0(n3099gat),
    .O(__472__)
  );
  LUT5 #(
    .INIT(32'h96696996)
  ) __984__ (
    .I4(__124__),
    .I3(__58__),
    .I2(__197__),
    .I1(__141__),
    .I0(__52__),
    .O(__473__)
  );
  LUT5 #(
    .INIT(32'h96696996)
  ) __985__ (
    .I4(__138__),
    .I3(__56__),
    .I2(__142__),
    .I1(__127__),
    .I0(__473__),
    .O(__474__)
  );
  LUT6 #(
    .INIT(64'h5555555755555555)
  ) __986__ (
    .I5(n3095gat),
    .I4(n3085gat),
    .I3(n3083gat),
    .I2(n3084gat),
    .I1(__383__),
    .I0(__474__),
    .O(__475__)
  );
  LUT4 #(
    .INIT(16'h007f)
  ) __987__ (
    .I3(__398__),
    .I2(__60__),
    .I1(__147__),
    .I0(__98__),
    .O(__476__)
  );
  LUT5 #(
    .INIT(32'h30cfaaaa)
  ) __988__ (
    .I4(__356__),
    .I3(__75__),
    .I2(__354__),
    .I1(__61__),
    .I0(n3066gat),
    .O(__477__)
  );
  LUT5 #(
    .INIT(32'h00008000)
  ) __989__ (
    .I4(__122__),
    .I3(__125__),
    .I2(__119__),
    .I1(__121__),
    .I0(__120__),
    .O(__478__)
  );
  LUT4 #(
    .INIT(16'h8000)
  ) __990__ (
    .I3(__206__),
    .I2(__205__),
    .I1(__149__),
    .I0(__47__),
    .O(__479__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __991__ (
    .I1(__118__),
    .I0(__115__),
    .O(__480__)
  );
  LUT6 #(
    .INIT(64'h00000000efff0000)
  ) __992__ (
    .I5(__222__),
    .I4(__274__),
    .I3(__117__),
    .I2(__480__),
    .I1(__146__),
    .I0(__116__),
    .O(__481__)
  );
  LUT5 #(
    .INIT(32'h07080000)
  ) __993__ (
    .I4(__47__),
    .I3(__149__),
    .I2(__90__),
    .I1(__206__),
    .I0(__205__),
    .O(__482__)
  );
  LUT6 #(
    .INIT(64'haa00c0c000000000)
  ) __994__ (
    .I5(n3087gat),
    .I4(n3088gat),
    .I3(n3094gat),
    .I2(__235__),
    .I1(__375__),
    .I0(__373__),
    .O(__483__)
  );
  LUT3 #(
    .INIT(8'h7f)
  ) __995__ (
    .I2(__163__),
    .I1(__117__),
    .I0(__146__),
    .O(__484__)
  );
  LUT6 #(
    .INIT(64'hff0b00f4ffffffff)
  ) __996__ (
    .I5(__301__),
    .I4(__84__),
    .I3(__117__),
    .I2(__146__),
    .I1(__115__),
    .I0(__118__),
    .O(__485__)
  );
  LUT6 #(
    .INIT(64'h00008aaaa8aaaaaa)
  ) __997__ (
    .I5(__117__),
    .I4(__146__),
    .I3(__480__),
    .I2(__219__),
    .I1(__116__),
    .I0(__275__),
    .O(__486__)
  );
  LUT3 #(
    .INIT(8'hf4)
  ) __998__ (
    .I2(__369__),
    .I1(n3066gat),
    .I0(__376__),
    .O(__487__)
  );
  LUT5 #(
    .INIT(32'h000002a8)
  ) __999__ (
    .I4(__278__),
    .I3(__122__),
    .I2(__121__),
    .I1(__120__),
    .I0(__275__),
    .O(__488__)
  );
  LUT4 #(
    .INIT(16'hc3aa)
  ) __1000__ (
    .I3(__356__),
    .I2(__61__),
    .I1(__354__),
    .I0(n3067gat),
    .O(__489__)
  );
  LUT4 #(
    .INIT(16'hf888)
  ) __1001__ (
    .I3(__238__),
    .I2(n3074gat),
    .I1(__236__),
    .I0(n3065gat),
    .O(__490__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __1002__ (
    .I1(__75__),
    .I0(__61__),
    .O(__491__)
  );
  LUT6 #(
    .INIT(64'hfc0003ffaaaaaaaa)
  ) __1003__ (
    .I5(__356__),
    .I4(__74__),
    .I3(__436__),
    .I2(__81__),
    .I1(__491__),
    .I0(n3073gat),
    .O(__492__)
  );
  LUT3 #(
    .INIT(8'hf4)
  ) __1004__ (
    .I2(__369__),
    .I1(n3070gat),
    .I0(__376__),
    .O(__493__)
  );
  LUT6 #(
    .INIT(64'h4000000000000000)
  ) __1005__ (
    .I5(__191__),
    .I4(__193__),
    .I3(__332__),
    .I2(__466__),
    .I1(__231__),
    .I0(__187__),
    .O(__494__)
  );
  LUT4 #(
    .INIT(16'h0004)
  ) __1006__ (
    .I3(__79__),
    .I2(__77__),
    .I1(__232__),
    .I0(__80__),
    .O(__495__)
  );
  LUT6 #(
    .INIT(64'heeeeaaaaccccf00f)
  ) __1007__ (
    .I5(__238__),
    .I4(__236__),
    .I3(__76__),
    .I2(__495__),
    .I1(n3069gat),
    .I0(n3078gat),
    .O(__496__)
  );
  LUT6 #(
    .INIT(64'hfeeefcccfaaaf000)
  ) __1008__ (
    .I5(n3093gat),
    .I4(n3095gat),
    .I3(__229__),
    .I2(__368__),
    .I1(n3071gat),
    .I0(n3080gat),
    .O(__497__)
  );
  LUT6 #(
    .INIT(64'hbfff0f0fbfbf0f0f)
  ) __1009__ (
    .I5(__249__),
    .I4(__248__),
    .I3(__138__),
    .I2(__226__),
    .I1(__351__),
    .I0(__349__),
    .O(__498__)
  );
  LUT6 #(
    .INIT(64'hfeeefcccfaaaf000)
  ) __1010__ (
    .I5(n3093gat),
    .I4(n3095gat),
    .I3(__229__),
    .I2(__368__),
    .I1(n3066gat),
    .I0(n3075gat),
    .O(__499__)
  );
  LUT6 #(
    .INIT(64'hfeeefcccfaaaf000)
  ) __1011__ (
    .I5(n3093gat),
    .I4(n3095gat),
    .I3(__229__),
    .I2(__368__),
    .I1(n3068gat),
    .I0(n3077gat),
    .O(__500__)
  );
  LUT6 #(
    .INIT(64'h4000000000000000)
  ) __1012__ (
    .I5(__125__),
    .I4(__119__),
    .I3(__121__),
    .I2(__122__),
    .I1(__99__),
    .I0(__120__),
    .O(__501__)
  );
  LUT5 #(
    .INIT(32'h5556ffff)
  ) __1013__ (
    .I4(__167__),
    .I3(__118__),
    .I2(__117__),
    .I1(__146__),
    .I0(__115__),
    .O(__502__)
  );
  LUT6 #(
    .INIT(64'h0808080808080880)
  ) __1014__ (
    .I5(__118__),
    .I4(__117__),
    .I3(__146__),
    .I2(__115__),
    .I1(__262__),
    .I0(__275__),
    .O(__503__)
  );
  LUT5 #(
    .INIT(32'h13203300)
  ) __1015__ (
    .I4(__206__),
    .I3(__149__),
    .I2(__205__),
    .I1(__90__),
    .I0(__47__),
    .O(__504__)
  );
  LUT6 #(
    .INIT(64'heeeeaaaaccccf00f)
  ) __1016__ (
    .I5(__238__),
    .I4(__236__),
    .I3(__79__),
    .I2(__232__),
    .I1(n3072gat),
    .I0(n3081gat),
    .O(__505__)
  );
  LUT5 #(
    .INIT(32'h00088880)
  ) __1017__ (
    .I4(__118__),
    .I3(__117__),
    .I2(__146__),
    .I1(__262__),
    .I0(__275__),
    .O(__506__)
  );
  LUT6 #(
    .INIT(64'h0000b0bbb0bbb0bb)
  ) __1018__ (
    .I5(__468__),
    .I4(__240__),
    .I3(__242__),
    .I2(__200__),
    .I1(__249__),
    .I0(__174__),
    .O(__507__)
  );
  LUT6 #(
    .INIT(64'h3232ff322222fff2)
  ) __1019__ (
    .I5(n3088gat),
    .I4(__259__),
    .I3(__293__),
    .I2(__287__),
    .I1(__507__),
    .I0(__248__),
    .O(__508__)
  );
  LUT4 #(
    .INIT(16'hf888)
  ) __1020__ (
    .I3(n3093gat),
    .I2(n3068gat),
    .I1(n3095gat),
    .I0(n3077gat),
    .O(__509__)
  );
  LUT4 #(
    .INIT(16'hf888)
  ) __1021__ (
    .I3(n3072gat),
    .I2(n3093gat),
    .I1(n3095gat),
    .I0(n3081gat),
    .O(__510__)
  );
  assign n3150gat = __359__;
  assign n3127gat = __25__;
  assign n3133gat = __295__;
  assign n3149gat = __220__;
  assign n3125gat = __260__;
  assign n3118gat = __250__;
  assign n3143gat = __450__;
  assign n3146gat = __364__;
  assign n3123gat = __347__;
  assign n3132gat = __352__;
  assign n3106gat = __35__;
  assign n3119gat = __498__;
  assign n3124gat = __444__;
  assign n3136gat = __307__;
  assign n3145gat = __476__;
  assign n3117gat = __435__;
  assign n3114gat = __420__;
  assign n3104gat = __439__;
  assign n3134gat = __384__;
  assign n3128gat = __24__;
  assign n3116gat = __468__;
  assign n3105gat = __429__;
  assign n3120gat = __432__;
  assign n3126gat = __26__;
  assign n3121gat = __475__;
  assign n3135gat = __394__;
  assign n3144gat = __339__;
  assign n3108gat = __410__;
  assign n3113gat = __371__;
  assign n3107gat = __227__;
  assign n3109gat = __502__;
  assign n3131gat = __454__;
  assign n3137gat = __449__;
  assign n3111gat = __484__;
  assign n3110gat = __408__;
  assign n3138gat = __494__;
  assign n3130gat = __419__;
  assign n3129gat = __508__;
  assign n3151gat = __299__;
  assign n3141gat = __465__;
  assign n3142gat = __465__;
  assign n3112gat = 1'b1;
  assign n3115gat = 1'b1;
  assign n3147gat = 1'b1;
  assign n3148gat = 1'b1;
  assign n3152gat = 1'b1;
  assign n3139gat = __405__;
  assign n3140gat = __405__;
  assign n3122gat = __345__;
endmodule
