// IWLS benchmark module "CM162" printed on Wed May 29 16:31:28 2002
module cm162a(a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s);
input
  a,
  b,
  c,
  d,
  e,
  f,
  g,
  h,
  i,
  j,
  k,
  l,
  m,
  n;
output
  o,
  p,
  q,
  r,
  s;
wire
  o0,
  d0,
  p0,
  e0,
  q0,
  f0,
  r0,
  g0,
  s0,
  \[0] ,
  \[1] ,
  j0,
  \[2] ,
  k0,
  \[3] ,
  l0,
  \[4] ,
  m0,
  n0;
assign
  o0 = ~l0 & ~n0,
  d0 = ~o0 & ~j0,
  p0 = (~l & ~r0) | (l & r0),
  e0 = (~i & l0) | (i & ~l0),
  q0 = (~m & ~s0) | (m & s0),
  f0 = ~o0 & ~k0,
  r0 = ~k & (~i & ~l0),
  g0 = (~k & ~m0) | (k & m0),
  s0 = ~k & (~i & (~l0 & ~l)),
  \[0]  = (~f0 & ~d0) | ((~f0 & ~a) | ((~e0 & ~d0) | (~e0 & ~a))),
  \[1]  = (~f0 & ~d0) | ((~f0 & ~b) | ((~g0 & ~d0) | (~g0 & ~b))),
  o = \[0] ,
  p = \[1] ,
  q = \[2] ,
  r = \[3] ,
  s = \[4] ,
  j0 = ~f | d,
  \[2]  = (~f0 & ~d0) | ((~f0 & ~g) | ((~p0 & ~d0) | (~p0 & ~g))),
  k0 = ~f | ~d,
  \[3]  = (~f0 & ~d0) | ((~f0 & ~h) | ((~q0 & ~d0) | (~q0 & ~h))),
  l0 = ~e | (~d | ~c),
  \[4]  = e & ~n0,
  m0 = ~l0 & ~i,
  n0 = ~n | ~j;
endmodule

