// IWLS benchmark module "x3.blif" printed on Wed May 29 17:30:37 2002
module x3 (b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, \xx , y, z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0, o0, r0, s0, t0, u0, v0, w0, x0, y0, z0, a1, b1, c1, d1, e1, f1, g1, h1, i1, j1, k1, l1, m1, n1, o1, p1, q1, r1, s1, t1, u1, v1, w1, x1, y1, z1, a2, b2, c2, d2, e2, f2, g2, h2, i2, j2, k2, l2, m2, n2, o2, p2, q2, r2, s2, t2, u2, v2, w2, x2, y2, z2, a3, b3, c3, d3, e3, f3, g3, h3, i3, j3, k3, l3, m3, n3, o3, p3, q3, r3, s3, t3, u3, v3, w3, x3, y3, z3, a4, b4, c4, d4, e4, f4, g4, h4, i4, j4, k4, l4, m4, n4, o4, p4, q4, r4, s4, t4, u4, v4, w4, x4, y4, z4, a5, b5, c5, d5, e5, f5, g5, h5, i5, j5, k5, l5, m5, n5, o5, p5, q5, r5, s5, t5, u5, v5, w5, x5, y5, z5, a6, b6, c6, d6, e6, f6, g6, h6, i6, j6, k6, l6, m6, n6, o6, p6, q6, r6, s6, t6, u6, v6, w6, x6, y6, z6, a7, b7, c7, d7, e7, f7, g7, h7, i7, j7, k7, l7, m7, n7, o7, p7, q7, r7, s7, t7, u7, v7, w7, x7, y7, z7, a8, b8, c8);
input
  b,
  c,
  d,
  e,
  f,
  g,
  h,
  i,
  j,
  k,
  l,
  m,
  n,
  o,
  p,
  q,
  r,
  s,
  t,
  u,
  v,
  w,
  \xx ,
  y,
  z,
  a0,
  a1,
  a2,
  a3,
  a4,
  b0,
  b1,
  b2,
  b3,
  b4,
  c0,
  c1,
  c2,
  c3,
  c4,
  d0,
  d1,
  d2,
  d3,
  d4,
  e0,
  e1,
  e2,
  e3,
  e4,
  f0,
  f1,
  f2,
  f3,
  f4,
  g0,
  g1,
  g2,
  g3,
  g4,
  h0,
  h1,
  h2,
  h3,
  h4,
  i0,
  i1,
  i2,
  i3,
  j0,
  j1,
  j2,
  j3,
  k0,
  k1,
  k2,
  k3,
  l0,
  l1,
  l2,
  l3,
  m0,
  m1,
  m2,
  m3,
  n0,
  n1,
  n2,
  n3,
  o0,
  o1,
  o2,
  o3,
  p1,
  p2,
  p3,
  q1,
  q2,
  q3,
  r0,
  r1,
  r2,
  r3,
  s0,
  s1,
  s2,
  s3,
  t0,
  t1,
  t2,
  t3,
  u0,
  u1,
  u2,
  u3,
  v0,
  v1,
  v2,
  v3,
  w0,
  w1,
  w2,
  w3,
  x0,
  x1,
  x2,
  x3,
  y0,
  y1,
  y2,
  y3,
  z0,
  z1,
  z2,
  z3;
output
  a5,
  a6,
  a7,
  a8,
  b5,
  b6,
  b7,
  b8,
  c5,
  c6,
  c7,
  c8,
  d5,
  d6,
  d7,
  e5,
  e6,
  e7,
  f5,
  f6,
  f7,
  g5,
  g6,
  g7,
  h5,
  h6,
  h7,
  i4,
  i5,
  i6,
  i7,
  j4,
  j5,
  j6,
  j7,
  k4,
  k5,
  k6,
  k7,
  l4,
  l5,
  l6,
  l7,
  m4,
  m5,
  m6,
  m7,
  n4,
  n5,
  n6,
  n7,
  o4,
  o5,
  o6,
  o7,
  p4,
  p5,
  p6,
  p7,
  q4,
  q5,
  q6,
  q7,
  r4,
  r5,
  r6,
  r7,
  s4,
  s5,
  s6,
  s7,
  t4,
  t5,
  t6,
  t7,
  u4,
  u5,
  u6,
  u7,
  v4,
  v5,
  v6,
  v7,
  w4,
  w5,
  w6,
  w7,
  x4,
  x5,
  x6,
  x7,
  y4,
  y5,
  y6,
  y7,
  z4,
  z5,
  z6,
  z7;
wire
  \[77] ,
  \[78] ,
  \[79] ,
  h16,
  h17,
  h18,
  h19,
  h20,
  h21,
  h22,
  h23,
  h24,
  h25,
  \[80] ,
  \[81] ,
  \[82] ,
  \[83] ,
  \[84] ,
  x16,
  x17,
  x18,
  x19,
  \[85] ,
  x21,
  x22,
  x23,
  x24,
  \[86] ,
  \[87] ,
  \[88] ,
  \[89] ,
  i12,
  i14,
  i15,
  i16,
  i17,
  i18,
  i19,
  i21,
  i22,
  i23,
  i25,
  \[90] ,
  \[91] ,
  \[92] ,
  \[93] ,
  \[94] ,
  y11,
  y13,
  y14,
  y15,
  y16,
  y17,
  y19,
  \[95] ,
  y20,
  y21,
  y22,
  y23,
  y24,
  \[96] ,
  \[97] ,
  \[98] ,
  j12,
  j16,
  j17,
  j18,
  j19,
  j20,
  j21,
  j22,
  j23,
  j24,
  j25,
  \[0] ,
  \[1] ,
  \[2] ,
  \[3] ,
  \[4] ,
  z11,
  z12,
  \[5] ,
  z17,
  z18,
  z21,
  z22,
  z24,
  \[6] ,
  \[7] ,
  \[8] ,
  \[9] ,
  k12,
  k14,
  k15,
  k17,
  k18,
  k21,
  k22,
  k24,
  l12,
  l16,
  l19,
  l20,
  l21,
  l23,
  l24,
  l25,
  m13,
  m14,
  m15,
  m16,
  m21,
  m22,
  m23,
  m24,
  m25,
  n12,
  n16,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  o12,
  o14,
  o15,
  o16,
  o18,
  o19,
  o21,
  o22,
  o23,
  o24,
  o25,
  p12,
  p16,
  p18,
  p20,
  p21,
  p22,
  p24,
  a13,
  a14,
  a15,
  a16,
  a18,
  a19,
  a20,
  a21,
  a22,
  a24,
  a25,
  \[10] ,
  \[11] ,
  \[12] ,
  \[13] ,
  \[14] ,
  q12,
  q13,
  q14,
  q15,
  q16,
  q18,
  q19,
  \[15] ,
  q21,
  q23,
  q24,
  \[16] ,
  \[17] ,
  \[18] ,
  \[19] ,
  b13,
  b18,
  b19,
  b23,
  b24,
  b25,
  \[20] ,
  \[21] ,
  \[22] ,
  \[23] ,
  \[24] ,
  r12,
  r16,
  r17,
  r18,
  r19,
  \[25] ,
  r22,
  r23,
  r24,
  \[26] ,
  \[27] ,
  \[28] ,
  \[29] ,
  c12,
  c13,
  c14,
  c15,
  c16,
  c17,
  c19,
  c21,
  c22,
  c23,
  c24,
  c25,
  \[30] ,
  \[31] ,
  \[32] ,
  \[33] ,
  \[34] ,
  s13,
  s14,
  s15,
  s16,
  s18,
  s19,
  \[35] ,
  s20,
  s21,
  s22,
  s23,
  s24,
  \[36] ,
  \[37] ,
  \[38] ,
  \[39] ,
  d16,
  d17,
  d18,
  d20,
  d22,
  d23,
  d24,
  d25,
  \[40] ,
  \[41] ,
  \[42] ,
  \[43] ,
  \[44] ,
  t16,
  \[45] ,
  t21,
  t22,
  t23,
  t24,
  \[46] ,
  \[47] ,
  \[48] ,
  \[49] ,
  e14,
  e15,
  e17,
  e18,
  e19,
  e21,
  e22,
  e23,
  e25,
  \[50] ,
  \[51] ,
  \[52] ,
  \[53] ,
  \[54] ,
  u13,
  u14,
  u15,
  u17,
  u18,
  u19,
  \[55] ,
  u20,
  u21,
  u22,
  u24,
  \[56] ,
  \[57] ,
  \[58] ,
  \[59] ,
  f16,
  f18,
  f20,
  f22,
  f24,
  f25,
  \[60] ,
  \[61] ,
  \[62] ,
  \[63] ,
  \[64] ,
  v16,
  v17,
  v19,
  \[65] ,
  v21,
  v23,
  v24,
  \[66] ,
  \[67] ,
  \[68] ,
  \[69] ,
  g14,
  g15,
  g16,
  g17,
  g18,
  g21,
  g23,
  g24,
  g25,
  \[70] ,
  \[71] ,
  \[72] ,
  \[73] ,
  \[74] ,
  w12,
  w13,
  w15,
  w16,
  w17,
  w18,
  w19,
  \[75] ,
  w20,
  w22,
  w23,
  w24,
  \[76] ;
assign
  \[77]  = (~d22 & (~y1 & ~c22)) | ((~d22 & (~y1 & ~h21)) | (~d22 & (~y1 & c))),
  \[78]  = (~i22 & (~y1 & ~h22)) | ((~i22 & (~y1 & ~h21)) | (~i22 & (~y1 & c))),
  \[79]  = (~n22 & (~y1 & ~m22)) | ((~n22 & (~y1 & ~h21)) | (~n22 & (~y1 & c))),
  h16 = (~o16 & (~n16 & ~z12)) | ((~o16 & (~n16 & ~l16)) | ((~o16 & (~n16 & q12)) | ((~o16 & (~m16 & ~z12)) | ((~o16 & (~m16 & ~l16)) | ((~o16 & (~m16 & q12)) | ((~o16 & (q2 & ~z12)) | ((~o16 & (q2 & ~l16)) | (~o16 & (q2 & q12))))))))),
  h17 = l0 | n0,
  h18 = (~i18 & (~a2 & ~w16)) | ((~i18 & (~a2 & ~v16)) | (~i18 & (~a2 & h0))),
  h19 = (~i19 & (~c & ~d)) | y1,
  h20 = (~w2 & (~h & f)) | ((~v2 & ~f) | y1),
  h21 = ~d & ~e,
  h22 = (~k22 & ~n16) | ((~k22 & x1) | (~k22 & ~o3)),
  h23 = (~b1 & (~e & d)) | ((~r1 & e) | ~i23),
  h24 = ~l21 | h3,
  h25 = o2 | p2,
  \[80]  = (~s22 & (~y1 & ~r22)) | ((~s22 & (~y1 & ~h21)) | (~s22 & (~y1 & c))),
  \[81]  = (~x22 & (~y1 & ~w22)) | ((~x22 & (~y1 & ~h21)) | (~x22 & (~y1 & c))),
  \[82]  = (~c23 & (~y1 & ~b23)) | ((~c23 & (~y1 & ~h21)) | (~c23 & (~y1 & c))),
  \[83]  = (~h23 & (~y1 & ~g23)) | ((~h23 & (~y1 & ~h21)) | (~h23 & (~y1 & c))),
  \[84]  = (~m23 & (~y1 & ~l23)) | ((~m23 & (~y1 & ~h21)) | (~m23 & (~y1 & c))),
  x16 = (h4 & ~y16) | ((a2 & ~f2) | (a2 & ~e2)),
  x17 = n0 | ~c2,
  x18 = (z18 & (k2 & ~x1)) | ((~z18 & ~k2) | y1),
  x19 = (~i25 & (j2 & ~p2)) | (~i25 & ~o2),
  \[85]  = (~r23 & (~y1 & ~q23)) | ((~r23 & (~y1 & ~h21)) | (~r23 & (~y1 & c))),
  x21 = (~a22 & ~n16) | ((~a22 & x1) | (~a22 & ~m3)),
  x22 = (~z0 & (~e & d)) | ((~p1 & e) | ~y22),
  x23 = ~l21 | f3,
  x24 = ~u24 | (~m24 | ~t24),
  \[86]  = (~w23 & (~y1 & ~v23)) | ((~w23 & (~y1 & ~h21)) | (~w23 & (~y1 & c))),
  \[87]  = (~b24 & (~y1 & ~a24)) | ((~b24 & (~y1 & ~h21)) | (~b24 & (~y1 & c))),
  \[88]  = (~g24 & (~y1 & ~f24)) | ((~g24 & (~y1 & ~h21)) | (~g24 & (~y1 & c))),
  \[89]  = ~l0 & (~n0 & ~y3),
  i12 = ~q12 | y1,
  i14 = (r & (~l & i)) | ((~b1 & ~r) | ((~b1 & ~l) | (~b1 & ~i))),
  i15 = (~b0 & (~z & s)) | ((~n1 & b0) | ((~n1 & ~z) | (~n1 & ~s))),
  i16 = ~j16 | (~q2 | ~r2),
  i17 = y3 & (z3 & a4),
  i18 = ~y16 & h4,
  i19 = e | (~x1 | m2),
  i21 = (~m21 & ~n16) | ((~m21 & x1) | (~m21 & ~j3)),
  i22 = (~w0 & (~e & d)) | ((~m1 & e) | ~j22),
  i23 = ~l21 | c3,
  i25 = ~j25 | ~n2,
  \[90]  = (~j24 & y3) | (~j24 & z3),
  \[91]  = (~k24 & (y3 & z3)) | (~k24 & a4),
  \[92]  = (~h17 & (~w17 & ~l24)) | ((~h17 & (~w17 & ~y3)) | ((~h17 & (~w17 & ~z3)) | ((~h17 & (b4 & ~l24)) | ((~h17 & (b4 & ~y3)) | (~h17 & (b4 & ~z3)))))),
  \[93]  = (~h17 & (~n24 & ~m24)) | ((~h17 & (~n24 & ~y3)) | ((~h17 & (~n24 & ~z3)) | ((~h17 & (c4 & ~m24)) | ((~h17 & (c4 & ~y3)) | (~h17 & (c4 & ~z3)))))),
  \[94]  = (~h17 & (~p24 & ~j17)) | ((~h17 & (~p24 & ~o24)) | ((~h17 & (~p24 & ~y3)) | ((~h17 & (d4 & ~j17)) | ((~h17 & (d4 & ~o24)) | (~h17 & (d4 & ~y3)))))),
  y11 = d | e,
  y13 = (~r & (~o & i)) | ((~w0 & r) | ((~w0 & ~o) | (~w0 & ~i))),
  y14 = (~b0 & (~u & s)) | ((~i1 & b0) | ((~i1 & ~u) | (~i1 & ~s))),
  y15 = (b0 & (~z & s)) | ((~v1 & ~b0) | ((~v1 & ~z) | (~v1 & ~s))),
  y16 = ~a25 | (~z3 | ~y3),
  y17 = ~b18 & (~a18 & ~z17),
  y19 = (~i2 & ~x19) | (~q2 | x1),
  \[95]  = (~h17 & (~r24 & ~q24)) | ((~h17 & (~r24 & ~d17)) | ((~h17 & (~r24 & ~y3)) | ((~h17 & (e4 & ~q24)) | ((~h17 & (e4 & ~d17)) | (~h17 & (e4 & ~y3)))))),
  y20 = (h & (~e3 & f)) | ((~d3 & ~f) | y1),
  y21 = (~u0 & (~e & d)) | ((~k1 & e) | ~z21),
  y22 = ~l21 | a3,
  y23 = (v3 & (~k2 & ~j2)) | (v3 & x1),
  y24 = (h2 & g2) | (~b | n0),
  \[96]  = (~h17 & (~v24 & ~u24)) | ((~h17 & (~v24 & ~m24)) | ((~h17 & (~v24 & ~t24)) | ((~h17 & (f4 & ~u24)) | ((~h17 & (f4 & ~m24)) | (~h17 & (f4 & ~t24)))))),
  \[97]  = (~h17 & (~x24 & ~w24)) | ((~h17 & (~x24 & ~s24)) | ((~h17 & (~x24 & ~i17)) | ((~h17 & (g4 & ~w24)) | ((~h17 & (g4 & ~s24)) | (~h17 & (g4 & ~i17)))))),
  \[98]  = (~y24 & (l0 & d2)) | (~y24 & h4),
  j12 = a2 | (j2 | k2),
  j16 = ~x1 & (~y1 & i2),
  j17 = b4 & (c4 & d4),
  j18 = i0 | j0,
  j19 = m2 & n2,
  j20 = (~x2 & (~h & f)) | ((~w2 & ~f) | y1),
  j21 = (~r0 & (~e & d)) | ((~h1 & e) | ~k21),
  j22 = ~l21 | x2,
  j23 = (s3 & (~k2 & ~j2)) | (s3 & x1),
  j24 = (z3 & y3) | (l0 | n0),
  j25 = (~m2 & (l2 & p2)) | ((~m2 & (l2 & o2)) | (~m2 & (l2 & ~g0))),
  \[0]  = ~z24,
  \[1]  = (~z11 & (~y11 & ~c)) | y1,
  \[2]  = (w12 & (~l12 & ~x1)) | ((~k12 & (~j12 & ~i12)) | ~n12),
  \[3]  = (g2 & (h2 & ~n0)) | (c2 & ~n0),
  \[4]  = ~m13 & ~y1,
  z11 = (~o0 & ~c12) | ((~o0 & x1) | (~o0 & ~i2)),
  z12 = (~r2 & ~q2) | ~i2,
  \[5]  = ~q13 & ~y1,
  z17 = ~d18 | (~b2 | ~y3),
  z18 = (~o25 & (~o2 & ~n25)) | (~o25 & (~o2 & p2)),
  z21 = ~l21 | v2,
  z22 = (q3 & (~k2 & ~j2)) | (q3 & x1),
  z24 = x1 & ~a2,
  \[6]  = ~s13 & ~y1,
  \[7]  = ~u13 & ~y1,
  \[8]  = ~w13 & ~y1,
  \[9]  = ~y13 & ~y1,
  k12 = (i2 & q2) | (i2 & r2),
  k14 = (r & (~m & i)) | ((~c1 & ~r) | ((~c1 & ~m) | (~c1 & ~i))),
  k15 = (~b0 & (~a0 & s)) | ((~o1 & b0) | ((~o1 & ~a0) | (~o1 & ~s))),
  k17 = ~e4 & (~f4 & ~g4),
  k18 = k0 | (~l0 | ~d2),
  k21 = ~l21 | s2,
  k22 = (n3 & (~k2 & ~j2)) | (n3 & x1),
  k24 = (a4 & (z3 & y3)) | (l0 | n0),
  l12 = y1 | a2,
  l16 = ~j2 & ~k2,
  l19 = (~c16 & (~c & ~d)) | ~n19,
  l20 = (~y2 & (~h & f)) | ((~x2 & ~f) | y1),
  l21 = c & (~d & ~e),
  l23 = (~o23 & ~n16) | ((~o23 & x1) | (~o23 & ~u3)),
  l24 = a4 & b4,
  l25 = (~e0 & (~f0 & ~o2)) | (~m25 | ~n2),
  m13 = (~r & (~j & i)) | ((~r0 & r) | ((~r0 & ~j) | (~r0 & ~i))),
  m14 = (r & (~n & i)) | ((~d1 & ~r) | ((~d1 & ~n) | (~d1 & ~i))),
  m15 = (b0 & (~t & s)) | ((~p1 & ~b0) | ((~p1 & ~t) | (~p1 & ~s))),
  m16 = ~r2 & ~i3,
  m21 = (i3 & (~k2 & ~j2)) | (i3 & x1),
  m22 = (~p22 & ~n16) | ((~p22 & x1) | (~p22 & ~p3)),
  m23 = (~c1 & (~e & d)) | ((~s1 & e) | ~n23),
  m24 = a4 & (b4 & c4),
  m25 = (~m2 & (l2 & ~o2)) | (~m2 & (l2 & j2)),
  n12 = (~r12 & ~p12) | ((~r12 & ~o12) | ((~r12 & ~m0) | ((~q12 & ~p12) | ((~q12 & ~o12) | ((~q12 & ~m0) | ((~x1 & ~p12) | ((~x1 & ~o12) | (~x1 & ~m0)))))))),
  n16 = j2 | k2,
  n19 = l2 & m2,
  n20 = (~z2 & (~h & f)) | ((~y2 & ~f) | y1),
  n21 = (~q21 & ~n16) | ((~q21 & x1) | (~q21 & ~k3)),
  n22 = (~x0 & (~e & d)) | ((~n1 & e) | ~o22),
  n23 = ~l21 | d3,
  n24 = ~l24 | (~y3 | ~z3),
  n25 = e0 | (f0 | ~g0),
  a5 = \[18] ,
  a6 = \[44] ,
  a7 = \[70] ,
  a8 = \[96] ,
  b5 = \[19] ,
  b6 = \[45] ,
  b7 = \[71] ,
  b8 = \[97] ,
  c5 = \[20] ,
  c6 = \[46] ,
  c7 = \[72] ,
  c8 = \[98] ,
  d5 = \[21] ,
  d6 = \[47] ,
  d7 = \[73] ,
  e5 = \[22] ,
  e6 = \[48] ,
  e7 = \[74] ,
  f5 = \[23] ,
  f6 = \[49] ,
  f7 = \[75] ,
  g5 = \[24] ,
  g6 = \[50] ,
  g7 = \[76] ,
  h5 = \[25] ,
  h6 = \[51] ,
  h7 = \[77] ,
  i4 = \[0] ,
  i5 = \[26] ,
  i6 = \[52] ,
  i7 = \[78] ,
  j4 = \[1] ,
  j5 = \[27] ,
  j6 = \[53] ,
  j7 = \[79] ,
  k4 = \[2] ,
  k5 = \[28] ,
  k6 = \[54] ,
  k7 = \[80] ,
  l4 = \[3] ,
  l5 = \[29] ,
  l6 = \[55] ,
  l7 = \[81] ,
  m4 = \[4] ,
  m5 = \[30] ,
  m6 = \[56] ,
  m7 = \[82] ,
  n4 = \[5] ,
  n5 = \[31] ,
  n6 = \[57] ,
  n7 = \[83] ,
  o4 = \[6] ,
  o5 = \[32] ,
  o6 = \[58] ,
  o7 = \[84] ,
  o12 = ~y1 & a2,
  o14 = (r & (~o & i)) | ((~e1 & ~r) | ((~e1 & ~o) | (~e1 & ~i))),
  o15 = (b0 & (~u & s)) | ((~q1 & ~b0) | ((~q1 & ~u) | (~q1 & ~s))),
  o16 = (~l16 & (~i2 & ~i3)) | ~p16,
  o18 = a2 | ~f2,
  o19 = m2 & (n2 & o2),
  p4 = \[7] ,
  p5 = \[33] ,
  p6 = \[59] ,
  o21 = (~s0 & (~e & d)) | ((~i1 & e) | ~p21),
  p7 = \[85] ,
  o22 = ~l21 | y2,
  o23 = (t3 & (~k2 & ~j2)) | (t3 & x1),
  o24 = z3 & a4,
  o25 = ~l2 | (m2 | ~n2),
  q4 = \[8] ,
  q5 = \[34] ,
  q6 = \[60] ,
  q7 = \[86] ,
  r4 = \[9] ,
  r5 = \[35] ,
  r6 = \[61] ,
  r7 = \[87] ,
  s4 = \[10] ,
  s5 = \[36] ,
  s6 = \[62] ,
  s7 = \[88] ,
  t4 = \[11] ,
  t5 = \[37] ,
  t6 = \[63] ,
  t7 = \[89] ,
  u4 = \[12] ,
  u5 = \[38] ,
  u6 = \[64] ,
  u7 = \[90] ,
  v4 = \[13] ,
  v5 = \[39] ,
  v6 = \[65] ,
  v7 = \[91] ,
  w4 = \[14] ,
  w5 = \[40] ,
  w6 = \[66] ,
  w7 = \[92] ,
  x4 = \[15] ,
  x5 = \[41] ,
  x6 = \[67] ,
  x7 = \[93] ,
  y4 = \[16] ,
  y5 = \[42] ,
  y6 = \[68] ,
  y7 = \[94] ,
  z4 = \[17] ,
  z5 = \[43] ,
  z6 = \[69] ,
  z7 = \[95] ,
  p12 = (~f2 & (e2 & ~d0)) | (f2 & (~e2 & d0)),
  p16 = (d0 & (~q2 & ~x1)) | ((d0 & (~x1 & ~c0)) | ((~r2 & (~q2 & ~x1)) | ((~r2 & (~x1 & ~c0)) | (~i2 & ~x1)))),
  p18 = ~e2 | f2,
  p20 = (~h & (~g & f)) | ((~z2 & ~f) | y1),
  p21 = ~l21 | t2,
  p22 = (o3 & (~k2 & ~j2)) | (o3 & x1),
  p24 = ~m24 | (~y3 | ~z3),
  a13 = (~r2 & c0) | ((r2 & z1) | (z1 & c0)),
  a14 = (~r & (~p & i)) | ((~x0 & r) | ((~x0 & ~p) | (~x0 & ~i))),
  a15 = (~b0 & (~v & s)) | ((~j1 & b0) | ((~j1 & ~v) | (~j1 & ~s))),
  a16 = (b0 & (~a0 & s)) | ((~w1 & ~b0) | ((~w1 & ~a0) | (~w1 & ~s))),
  a18 = ~z3 | (~a4 | ~b4),
  a19 = ~e19 | (c | d),
  a20 = (~t2 & (~h & f)) | ((~s2 & ~f) | y1),
  a21 = (h & (~f3 & f)) | ((~e3 & ~f) | y1),
  a22 = (l3 & (~k2 & ~j2)) | (l3 & x1),
  a24 = (~d24 & ~n16) | ((~d24 & x1) | (~d24 & ~x3)),
  a25 = ~b25 & (b4 & a4),
  \[10]  = ~a14 & ~y1,
  \[11]  = ~c14 & ~y1,
  \[12]  = ~e14 & ~y1,
  \[13]  = ~g14 & ~y1,
  \[14]  = ~i14 & ~y1,
  q12 = (~h25 & (~g25 & ~f25)) | ((~h25 & (~g25 & m2)) | (~h25 & (~f25 & ~m2))),
  q13 = (~r & (~k & i)) | ((~s0 & r) | ((~s0 & ~k) | (~s0 & ~i))),
  q14 = (r & (~p & i)) | ((~f1 & ~r) | ((~f1 & ~p) | (~f1 & ~i))),
  q15 = (b0 & (~v & s)) | ((~r1 & ~b0) | ((~r1 & ~v) | (~r1 & ~s))),
  q16 = ~r2 & i3,
  q18 = (~s18 & ~w16) | ((~s18 & ~v16) | (~s18 & h0)),
  q19 = (~c16 & (~c & ~d)) | ~r19,
  \[15]  = ~k14 & ~y1,
  q21 = (j3 & (~k2 & ~j2)) | (j3 & x1),
  q23 = (~t23 & ~n16) | ((~t23 & x1) | (~t23 & ~v3)),
  q24 = c4 & (~d4 & e4),
  \[16]  = ~m14 & ~y1,
  \[17]  = ~o14 & ~y1,
  \[18]  = ~q14 & ~y1,
  \[19]  = ~s14 & ~y1,
  b13 = (~c13 & r2) | (~c13 & ~i3),
  b18 = ~c4 | (~d4 | e4),
  b19 = ~c19 & (x1 & ~l2),
  b23 = (~e23 & ~n16) | ((~e23 & x1) | (~e23 & ~s3)),
  b24 = (~f1 & (~e & d)) | ((~v1 & e) | ~c24),
  b25 = (~h0 & ~d4) | (~c25 | ~c4),
  \[20]  = ~u14 & ~y1,
  \[21]  = ~y14 & ~y1,
  \[22]  = ~a15 & ~y1,
  \[23]  = ~c15 & ~y1,
  \[24]  = ~e15 & ~y1,
  r12 = ~y1 & ~a2,
  r16 = (~l16 & (~i2 & i3)) | ~s16,
  r17 = f4 | g4,
  r18 = n0 | (e2 | ~f2),
  r19 = l2 & (m2 & n2),
  \[25]  = ~g15 & ~y1,
  r22 = (~u22 & ~n16) | ((~u22 & x1) | (~u22 & ~q3)),
  r23 = (~d1 & (~e & d)) | ((~t1 & e) | ~s23),
  r24 = ~s24 | (~o24 | ~y3),
  \[26]  = ~i15 & ~y1,
  \[27]  = ~k15 & ~y1,
  \[28]  = ~m15 & ~y1,
  \[29]  = ~o15 & ~y1,
  c12 = q2 & r2,
  c13 = (i3 & (r2 & d0)) | ((r2 & (i2 & d0)) | ((i3 & q2) | ((i3 & ~i2) | (q2 & i2)))),
  c14 = (~r & (~q & i)) | ((~y0 & r) | ((~y0 & ~q) | (~y0 & ~i))),
  c15 = (~b0 & (~w & s)) | ((~k1 & b0) | ((~k1 & ~w) | (~k1 & ~s))),
  c16 = e | ~x1,
  c17 = ~r17 & (b2 & y3),
  c19 = c | (d | e),
  c21 = (h & (~g3 & f)) | ((~f3 & ~f) | y1),
  c22 = (~f22 & ~n16) | ((~f22 & x1) | (~f22 & ~n3)),
  c23 = (~a1 & (~e & d)) | ((~q1 & e) | ~d23),
  c24 = ~l21 | g3,
  c25 = (~d25 & (i0 & ~h0)) | ((~d25 & (i0 & ~d4)) | ((~d25 & (~e4 & ~h0)) | (~d25 & (~e4 & ~d4)))),
  \[30]  = ~q15 & ~y1,
  \[31]  = ~s15 & ~y1,
  \[32]  = ~u15 & ~y1,
  \[33]  = ~w15 & ~y1,
  \[34]  = ~y15 & ~y1,
  s13 = (~r & (~l & i)) | ((~t0 & r) | ((~t0 & ~l) | (~t0 & ~i))),
  s14 = (r & (~q & i)) | ((~g1 & ~r) | ((~g1 & ~q) | (~g1 & ~i))),
  s15 = (b0 & (~w & s)) | ((~s1 & ~b0) | ((~s1 & ~w) | (~s1 & ~s))),
  s16 = (c0 & ~r2) | ((c0 & ~d0) | ((~r2 & ~q2) | ((~q2 & ~d0) | ~i2))),
  s18 = (h4 & ~y16) | a2,
  s19 = n2 & (o2 & p2),
  \[35]  = ~a16 & ~y1,
  s20 = (h & (~b3 & f)) | ((~a3 & ~f) | y1),
  s21 = (~v21 & ~n16) | ((~v21 & x1) | (~v21 & ~l3)),
  s22 = (~y0 & (~e & d)) | ((~o1 & e) | ~t22),
  s23 = ~l21 | e3,
  s24 = b4 & (c4 & ~d4),
  \[36]  = (~c16 & (~c & ~d)) | y1,
  \[37]  = (~d16 & (~x1 & i2)) | n0,
  \[38]  = (~h16 & (~y1 & z1)) | ((~g16 & (~f16 & ~x1)) | ~i16),
  \[39]  = ~t16 & ~y1,
  d16 = ~q2 | ~r2,
  d17 = z3 & (a4 & b4),
  d18 = ~f4 & ~g4,
  d20 = (~u2 & (~h & f)) | ((~t2 & ~f) | y1),
  d22 = (~v0 & (~e & d)) | ((~l1 & e) | ~e22),
  d23 = ~l21 | b3,
  d24 = (w3 & (~k2 & ~j2)) | (w3 & x1),
  d25 = (~j0 & f4) | ((i0 & ~e4) | ~e25),
  \[40]  = (~h17 & (~g17 & ~e17)) | ((~h17 & (~g17 & ~d17)) | ((~h17 & (~g17 & ~c17)) | ((~h17 & (b2 & ~e17)) | ((~h17 & (b2 & ~d17)) | (~h17 & (b2 & ~c17)))))),
  \[41]  = (~y17 & (~x17 & ~l0)) | (~w17 & (~v17 & ~u17)),
  \[42]  = (~e18 & ~g2) | (~e18 & ~h2),
  \[43]  = (~h18 & (~e2 & ~n0)) | (~g18 & (~f18 & ~n0)),
  \[44]  = (~q18 & (~p18 & ~n0)) | ((~o18 & (~g18 & ~n0)) | ~r18),
  t16 = (~x16 & ~w16) | ((~x16 & ~v16) | (~x16 & h0)),
  \[45]  = ~n0 & h2,
  t21 = (~t0 & (~e & d)) | ((~j1 & e) | ~u21),
  t22 = ~l21 | z2,
  t23 = (u3 & (~k2 & ~j2)) | (u3 & x1),
  t24 = y3 & z3,
  \[46]  = l0 & ~n0,
  \[47]  = (x19 & (~y1 & ~x1)) | (i2 & ~y1),
  \[48]  = (~u18 & ~x1) | (~u18 & j2),
  \[49]  = (~x18 & ~x1) | (~x18 & k2),
  e14 = (r & (~j & i)) | ((~z0 & ~r) | ((~z0 & ~j) | (~z0 & ~i))),
  e15 = (~b0 & (~\xx  & s)) | ((~l1 & b0) | ((~l1 & ~\xx ) | (~l1 & ~s))),
  e17 = c4 & (d4 & ~e4),
  e18 = (~d2 & ~l0) | (~b | n0),
  e19 = ~e & x1,
  e21 = (h & (~h3 & f)) | ((~g3 & ~f) | y1),
  e22 = ~l21 | w2,
  e23 = (r3 & (~k2 & ~j2)) | (r3 & x1),
  e25 = (~g4 & (f4 & ~k0)) | ((~g4 & (~k0 & ~j0)) | ((g4 & (f4 & k0)) | (g4 & (k0 & ~j0)))),
  \[50]  = (~b19 & (~y1 & ~a19)) | (~b19 & (~y1 & ~l2)),
  \[51]  = (~h19 & (~a19 & m2)) | ((~h19 & (~a19 & l2)) | ((~h19 & (~m2 & l2)) | (~h19 & (m2 & ~l2)))),
  \[52]  = (~y1 & (~l19 & ~a19)) | ((~y1 & (~l19 & ~j19)) | ((~y1 & (~l19 & ~l2)) | ((~y1 & (n2 & ~a19)) | ((~y1 & (n2 & ~j19)) | (~y1 & (n2 & ~l2)))))),
  \[53]  = (~y1 & (~q19 & ~a19)) | ((~y1 & (~q19 & ~o19)) | ((~y1 & (~q19 & ~l2)) | ((~y1 & (o2 & ~a19)) | ((~y1 & (o2 & ~o19)) | (~y1 & (o2 & ~l2)))))),
  \[54]  = (~y1 & (~u19 & ~a19)) | ((~y1 & (~u19 & ~s19)) | ((~y1 & (~u19 & ~n19)) | ((~y1 & (p2 & ~a19)) | ((~y1 & (p2 & ~s19)) | (~y1 & (p2 & ~n19)))))),
  u13 = (~r & (~m & i)) | ((~u0 & r) | ((~u0 & ~m) | (~u0 & ~i))),
  u14 = (~b0 & (~t & s)) | ((~h1 & b0) | ((~h1 & ~t) | (~h1 & ~s))),
  u15 = (b0 & (~\xx  & s)) | ((~t1 & ~b0) | ((~t1 & ~\xx ) | (~t1 & ~s))),
  u17 = ~k17 | (~j17 | l0),
  u18 = (w18 & (j2 & ~x1)) | ((~w18 & ~j2) | y1),
  u19 = (~c16 & (~c & ~d)) | (~o19 | ~l2),
  \[55]  = (~w19 & ~v19) | ((~w19 & x1) | (~w19 & ~q2)),
  u20 = (h & (~c3 & f)) | ((~b3 & ~f) | y1),
  u21 = ~l21 | u2,
  u22 = (p3 & (~k2 & ~j2)) | (p3 & x1),
  u24 = ~d4 & (e4 & f4),
  \[56]  = (~y1 & (~y19 & ~v19)) | ((~y1 & (~y19 & ~c12)) | ((~y1 & (~y19 & x1)) | ((~y1 & (r2 & ~v19)) | ((~y1 & (r2 & ~c12)) | (~y1 & (r2 & x1)))))),
  \[57]  = (~a20 & ~h) | (~a20 & s2),
  \[58]  = (~d20 & ~h) | (~d20 & t2),
  \[59]  = (~f20 & ~h) | (~f20 & u2),
  f16 = y1 | z1,
  f18 = a2 | ~e2,
  f20 = (~v2 & (~h & f)) | ((~u2 & ~f) | y1),
  f22 = (m3 & (~k2 & ~j2)) | (m3 & x1),
  f24 = (j2 & ~x1) | ((k2 & ~x1) | ~x3),
  f25 = (~l2 & ~i0) | ((l2 & ~h0) | ((~i0 & ~h0) | ~n2)),
  \[60]  = (~h20 & ~h) | (~h20 & v2),
  \[61]  = (~j20 & ~h) | (~j20 & w2),
  \[62]  = (~l20 & ~h) | (~l20 & x2),
  \[63]  = (~n20 & ~h) | (~n20 & y2),
  \[64]  = (~p20 & ~h) | (~p20 & z2),
  v16 = ~i0 & ~j0,
  v17 = n0 | (~b2 | c2),
  v19 = x19 | i2,
  \[65]  = (~s20 & h) | (~s20 & a3),
  v21 = (k3 & (~k2 & ~j2)) | (k3 & x1),
  v23 = (~y23 & ~n16) | ((~y23 & x1) | (~y23 & ~w3)),
  v24 = ~q24 | (~d17 | ~y3),
  \[66]  = (~u20 & h) | (~u20 & b3),
  \[67]  = (~w20 & h) | (~w20 & c3),
  \[68]  = (~y20 & h) | (~y20 & d3),
  \[69]  = (~a21 & h) | (~a21 & e3),
  g14 = (r & (~k & i)) | ((~a1 & ~r) | ((~a1 & ~k) | (~a1 & ~i))),
  g15 = (~b0 & (~y & s)) | ((~m1 & b0) | ((~m1 & ~y) | (~m1 & ~s))),
  g16 = (~r16 & (~n16 & ~z12)) | ((~r16 & (~n16 & ~l16)) | ((~r16 & (~n16 & ~q12)) | ((~r16 & (~q16 & ~z12)) | ((~r16 & (~q16 & ~l16)) | ((~r16 & (~q16 & ~q12)) | ((~r16 & (q2 & ~z12)) | ((~r16 & (q2 & ~l16)) | (~r16 & (q2 & ~q12))))))))),
  g17 = ~k17 | (~j17 | ~i17),
  g18 = (~k18 & (~j18 & ~h0)) | (~y16 & h4),
  g21 = (h & (~g & f)) | ((~h3 & ~f) | y1),
  g23 = (~j23 & ~n16) | ((~j23 & x1) | (~j23 & ~t3)),
  g24 = (~g1 & (~e & d)) | ((~w1 & e) | ~h24),
  g25 = (~l2 & ~k0) | ((l2 & ~j0) | ((~k0 & ~j0) | n2)),
  \[70]  = (~c21 & h) | (~c21 & f3),
  \[71]  = (~e21 & h) | (~e21 & g3),
  \[72]  = (~g21 & h) | (~g21 & h3),
  \[73]  = (~j21 & (~y1 & ~i21)) | ((~j21 & (~y1 & ~h21)) | (~j21 & (~y1 & c))),
  \[74]  = (~o21 & (~y1 & ~n21)) | ((~o21 & (~y1 & ~h21)) | (~o21 & (~y1 & c))),
  w12 = (~b13 & (~a13 & ~z12)) | ((~b13 & (~a13 & j2)) | ((~b13 & (~a13 & k2)) | ((~b13 & (~i2 & ~z12)) | ((~b13 & (~i2 & j2)) | ((~b13 & (~i2 & k2)) | ((~b13 & (~q2 & ~z12)) | ((~b13 & (~q2 & j2)) | (~b13 & (~q2 & k2))))))))),
  w13 = (~r & (~n & i)) | ((~v0 & r) | ((~v0 & ~n) | (~v0 & ~i))),
  w15 = (b0 & (~y & s)) | ((~u1 & ~b0) | ((~u1 & ~y) | (~u1 & ~s))),
  w16 = ~k0 & (l0 & d2),
  w17 = ~y3 | (~z3 | ~a4),
  w18 = (~l25 & (~p2 & g0)) | (~l25 & (~p2 & o2)),
  w19 = (~x19 & (~q2 & ~i2)) | ((x1 & ~q2) | y1),
  \[75]  = (~t21 & (~y1 & ~s21)) | ((~t21 & (~y1 & ~h21)) | (~t21 & (~y1 & c))),
  w20 = (h & (~d3 & f)) | ((~c3 & ~f) | y1),
  w22 = (~z22 & ~n16) | ((~z22 & x1) | (~z22 & ~r3)),
  w23 = (~e1 & (~e & d)) | ((~u1 & e) | ~x23),
  w24 = e4 & (f4 & g4),
  \[76]  = (~y21 & (~y1 & ~x21)) | ((~y21 & (~y1 & ~h21)) | (~y21 & (~y1 & c)));
endmodule

