module s713 (
  CK,
  G1,
  G10,
  G11,
  G12,
  G13,
  G14,
  G15,
  G16,
  G17,
  G18,
  G19,
  G2,
  G20,
  G21,
  G22,
  G23,
  G24,
  G25,
  G26,
  G27,
  G28,
  G29,
  G3,
  G30,
  G31,
  G32,
  G33,
  G34,
  G35,
  G36,
  G4,
  G5,
  G6,
  G8,
  G9,
  G83,
  G89BF,
  G87BF,
  G91,
  G90,
  G95BF,
  G105BF,
  G88BF,
  G98BF,
  G92,
  G101BF,
  G104BF,
  G84,
  G103BF,
  G99BF,
  G96BF,
  G86BF,
  G85,
  G100BF,
  G107,
  G97BF,
  G94,
  G106BF
);
  input CK;
  wire CK;
  input G1;
  wire G1;
  input G10;
  wire G10;
  input G11;
  wire G11;
  input G12;
  wire G12;
  input G13;
  wire G13;
  input G14;
  wire G14;
  input G15;
  wire G15;
  input G16;
  wire G16;
  input G17;
  wire G17;
  input G18;
  wire G18;
  input G19;
  wire G19;
  input G2;
  wire G2;
  input G20;
  wire G20;
  input G21;
  wire G21;
  input G22;
  wire G22;
  input G23;
  wire G23;
  input G24;
  wire G24;
  input G25;
  wire G25;
  input G26;
  wire G26;
  input G27;
  wire G27;
  input G28;
  wire G28;
  input G29;
  wire G29;
  input G3;
  wire G3;
  input G30;
  wire G30;
  input G31;
  wire G31;
  input G32;
  wire G32;
  input G33;
  wire G33;
  input G34;
  wire G34;
  input G35;
  wire G35;
  input G36;
  wire G36;
  input G4;
  wire G4;
  input G5;
  wire G5;
  input G6;
  wire G6;
  input G8;
  wire G8;
  input G9;
  wire G9;
  output G83;
  wire G83;
  output G89BF;
  wire G89BF;
  output G87BF;
  wire G87BF;
  output G91;
  wire G91;
  output G90;
  wire G90;
  output G95BF;
  wire G95BF;
  output G105BF;
  wire G105BF;
  output G88BF;
  wire G88BF;
  output G98BF;
  wire G98BF;
  output G92;
  wire G92;
  output G101BF;
  wire G101BF;
  output G104BF;
  wire G104BF;
  output G84;
  wire G84;
  output G103BF;
  wire G103BF;
  output G99BF;
  wire G99BF;
  output G96BF;
  wire G96BF;
  output G86BF;
  wire G86BF;
  output G85;
  wire G85;
  output G100BF;
  wire G100BF;
  output G107;
  wire G107;
  output G97BF;
  wire G97BF;
  output G94;
  wire G94;
  output G106BF;
  wire G106BF;
  wire __0__;
  wire __1__;
  wire __2__;
  wire __3__;
  wire __4__;
  wire __5__;
  wire __6__;
  wire __7__;
  wire __8__;
  wire __9__;
  wire __10__;
  wire __11__;
  wire __12__;
  wire __13__;
  wire __14__;
  wire __15__;
  wire __16__;
  wire __18__;
  wire __19__;
  wire __20__;
  wire __21__;
  wire __22__;
  wire __23__;
  wire __24__;
  wire __25__;
  wire __26__;
  wire __27__;
  wire __28__;
  wire __29__;
  wire __30__;
  wire __31__;
  wire __32__;
  wire __33__;
  wire __34__;
  wire __35__;
  wire __36__;
  wire __37__;
  wire __39__;
  wire __40__;
  wire __41__;
  wire __42__;
  wire __43__;
  wire __44__;
  wire __45__;
  wire __46__;
  wire __47__;
  wire __48__;
  wire __49__;
  wire __50__;
  wire __51__;
  wire __52__;
  wire __53__;
  wire __54__;
  wire __55__;
  wire __56__;
  wire __57__;
  wire __58__;
  wire __59__;
  wire __60__;
  wire __61__;
  wire __62__;
  wire __63__;
  wire __64__;
  wire __65__;
  wire __66__;
  wire __67__;
  wire __68__;
  wire __69__;
  wire __70__;
  wire __71__;
  wire __72__;
  wire __73__;
  wire __74__;
  wire __75__;
  wire __76__;
  wire __77__;
  wire __78__;
  wire __79__;
  FDRE #(
    .INIT(1'bx)
  ) __80__ (
    .D(__41__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__0__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __81__ (
    .D(__20__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __82__ (
    .D(__63__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__2__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __83__ (
    .D(__37__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__3__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __84__ (
    .D(__58__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__4__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __85__ (
    .D(__66__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__5__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __86__ (
    .D(__69__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__6__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __87__ (
    .D(__51__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__7__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __88__ (
    .D(__50__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__8__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __89__ (
    .D(__52__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__9__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __90__ (
    .D(__56__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__10__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __91__ (
    .D(__34__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__11__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __92__ (
    .D(__23__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__12__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __93__ (
    .D(__77__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__13__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __94__ (
    .D(__45__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__14__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __95__ (
    .D(__59__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__15__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __96__ (
    .D(__54__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__16__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __98__ (
    .I1(G23),
    .I0(__4__),
    .O(__18__)
  );
  LUT6 #(
    .INIT(64'h555555555575ffff)
  ) __99__ (
    .I5(G3),
    .I4(G11),
    .I3(G9),
    .I2(G10),
    .I1(G13),
    .I0(__18__),
    .O(__19__)
  );
  LUT4 #(
    .INIT(16'h0cac)
  ) __100__ (
    .I3(G4),
    .I2(__19__),
    .I1(__0__),
    .I0(__1__),
    .O(__20__)
  );
  LUT3 #(
    .INIT(8'hf7)
  ) __101__ (
    .I2(G4),
    .I1(__2__),
    .I0(G35),
    .O(__21__)
  );
  LUT4 #(
    .INIT(16'h0e00)
  ) __102__ (
    .I3(G25),
    .I2(__9__),
    .I1(G3),
    .I0(G11),
    .O(__22__)
  );
  LUT6 #(
    .INIT(64'hff00bf0000000000)
  ) __103__ (
    .I5(__12__),
    .I4(G3),
    .I3(__22__),
    .I2(G9),
    .I1(G10),
    .I0(G13),
    .O(__23__)
  );
  LUT4 #(
    .INIT(16'h0040)
  ) __104__ (
    .I3(G3),
    .I2(G9),
    .I1(G10),
    .I0(G13),
    .O(__24__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __105__ (
    .I1(__15__),
    .I0(G2),
    .O(__25__)
  );
  LUT6 #(
    .INIT(64'hffff0000ef000000)
  ) __106__ (
    .I5(G3),
    .I4(G24),
    .I3(G11),
    .I2(G9),
    .I1(G10),
    .I0(G13),
    .O(__26__)
  );
  LUT6 #(
    .INIT(64'h0000bf000000ffff)
  ) __107__ (
    .I5(__26__),
    .I4(G3),
    .I3(__25__),
    .I2(__22__),
    .I1(__3__),
    .I0(__24__),
    .O(__27__)
  );
  LUT6 #(
    .INIT(64'haaaaaaaaaaa80000)
  ) __108__ (
    .I5(G3),
    .I4(G11),
    .I3(G9),
    .I2(G10),
    .I1(G13),
    .I0(G22),
    .O(__28__)
  );
  LUT6 #(
    .INIT(64'haa00aa20aa00aa00)
  ) __109__ (
    .I5(G25),
    .I4(__9__),
    .I3(G3),
    .I2(G11),
    .I1(__24__),
    .I0(__3__),
    .O(__29__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __110__ (
    .I1(G10),
    .I0(G13),
    .O(__30__)
  );
  LUT6 #(
    .INIT(64'hfbf0f0f000000000)
  ) __111__ (
    .I5(__13__),
    .I4(G11),
    .I3(__18__),
    .I2(G3),
    .I1(__30__),
    .I0(G9),
    .O(__31__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __112__ (
    .I1(__11__),
    .I0(G2),
    .O(__32__)
  );
  LUT6 #(
    .INIT(64'h0f0f0fdf0f0f0f0f)
  ) __113__ (
    .I5(__32__),
    .I4(__31__),
    .I3(__29__),
    .I2(__28__),
    .I1(__27__),
    .I0(__5__),
    .O(__33__)
  );
  LUT3 #(
    .INIT(8'hb0)
  ) __114__ (
    .I2(__14__),
    .I1(__33__),
    .I0(G3),
    .O(__34__)
  );
  LUT5 #(
    .INIT(32'h00ff40ff)
  ) __115__ (
    .I4(G3),
    .I3(__22__),
    .I2(G9),
    .I1(G10),
    .I0(G13),
    .O(__35__)
  );
  LUT5 #(
    .INIT(32'h00008a00)
  ) __116__ (
    .I4(__35__),
    .I3(__12__),
    .I2(__5__),
    .I1(__27__),
    .I0(G1),
    .O(__36__)
  );
  LUT6 #(
    .INIT(64'hff10ffff10101010)
  ) __117__ (
    .I5(__29__),
    .I4(G2),
    .I3(G1),
    .I2(__36__),
    .I1(__31__),
    .I0(__34__),
    .O(__37__)
  );
  LUT2 #(
    .INIT(4'h7)
  ) __119__ (
    .I1(__29__),
    .I0(G17),
    .O(__39__)
  );
  LUT6 #(
    .INIT(64'hfbf0000000000000)
  ) __120__ (
    .I5(__18__),
    .I4(__0__),
    .I3(G11),
    .I2(G3),
    .I1(__30__),
    .I0(G9),
    .O(__40__)
  );
  LUT3 #(
    .INIT(8'hfd)
  ) __121__ (
    .I2(G4),
    .I1(__40__),
    .I0(__1__),
    .O(__41__)
  );
  LUT4 #(
    .INIT(16'h000b)
  ) __122__ (
    .I3(__31__),
    .I2(__29__),
    .I1(__5__),
    .I0(__27__),
    .O(__42__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __123__ (
    .I1(__16__),
    .I0(G4),
    .O(__43__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __124__ (
    .I1(__6__),
    .I0(__33__),
    .O(__44__)
  );
  LUT6 #(
    .INIT(64'hffff808000ff0000)
  ) __125__ (
    .I5(G8),
    .I4(__34__),
    .I3(G2),
    .I2(__44__),
    .I1(__43__),
    .I0(__42__),
    .O(__45__)
  );
  LUT3 #(
    .INIT(8'h40)
  ) __126__ (
    .I2(__9__),
    .I1(G21),
    .I0(G4),
    .O(__46__)
  );
  LUT2 #(
    .INIT(4'h7)
  ) __127__ (
    .I1(__31__),
    .I0(G15),
    .O(__47__)
  );
  LUT4 #(
    .INIT(16'h5fdf)
  ) __128__ (
    .I3(G3),
    .I2(__14__),
    .I1(__33__),
    .I0(G14),
    .O(__48__)
  );
  LUT6 #(
    .INIT(64'h0b00ff00ffffffff)
  ) __129__ (
    .I5(__26__),
    .I4(__3__),
    .I3(__25__),
    .I2(G3),
    .I1(__22__),
    .I0(__24__),
    .O(__49__)
  );
  LUT4 #(
    .INIT(16'hff5d)
  ) __130__ (
    .I3(G4),
    .I2(__49__),
    .I1(__8__),
    .I0(__2__),
    .O(__50__)
  );
  LUT5 #(
    .INIT(32'h00008a00)
  ) __131__ (
    .I4(G2),
    .I3(__14__),
    .I2(__33__),
    .I1(G3),
    .I0(__42__),
    .O(__51__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __132__ (
    .I1(__29__),
    .I0(G2),
    .O(__52__)
  );
  LUT3 #(
    .INIT(8'hf7)
  ) __133__ (
    .I2(__33__),
    .I1(__6__),
    .I0(G30),
    .O(__53__)
  );
  LUT4 #(
    .INIT(16'h0cac)
  ) __134__ (
    .I3(G4),
    .I2(__33__),
    .I1(__6__),
    .I0(__16__),
    .O(__54__)
  );
  LUT3 #(
    .INIT(8'hf7)
  ) __135__ (
    .I2(__27__),
    .I1(__5__),
    .I0(G16),
    .O(__55__)
  );
  LUT4 #(
    .INIT(16'h0004)
  ) __136__ (
    .I3(G2),
    .I2(__29__),
    .I1(__5__),
    .I0(__27__),
    .O(__56__)
  );
  LUT3 #(
    .INIT(8'hf7)
  ) __137__ (
    .I2(G4),
    .I1(__1__),
    .I0(G33),
    .O(__57__)
  );
  LUT5 #(
    .INIT(32'h000000b0)
  ) __138__ (
    .I4(G2),
    .I3(__29__),
    .I2(__31__),
    .I1(__5__),
    .I0(__27__),
    .O(__58__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __139__ (
    .I1(__5__),
    .I0(__27__),
    .O(__59__)
  );
  LUT4 #(
    .INIT(16'h8000)
  ) __140__ (
    .I3(G11),
    .I2(G13),
    .I1(G12),
    .I0(G28),
    .O(__60__)
  );
  LUT2 #(
    .INIT(4'h7)
  ) __141__ (
    .I1(__40__),
    .I0(G32),
    .O(__61__)
  );
  LUT3 #(
    .INIT(8'hf7)
  ) __142__ (
    .I2(__49__),
    .I1(__8__),
    .I0(G34),
    .O(__62__)
  );
  LUT4 #(
    .INIT(16'h0cac)
  ) __143__ (
    .I3(G4),
    .I2(__49__),
    .I1(__8__),
    .I0(__2__),
    .O(__63__)
  );
  LUT3 #(
    .INIT(8'h40)
  ) __144__ (
    .I2(__4__),
    .I1(G19),
    .I0(G4),
    .O(__64__)
  );
  LUT5 #(
    .INIT(32'h00000040)
  ) __145__ (
    .I4(G4),
    .I3(__29__),
    .I2(__8__),
    .I1(__2__),
    .I0(__49__),
    .O(__65__)
  );
  LUT6 #(
    .INIT(64'hffff101000ff0000)
  ) __146__ (
    .I5(G6),
    .I4(__59__),
    .I3(G2),
    .I2(__65__),
    .I1(__31__),
    .I0(__34__),
    .O(__66__)
  );
  LUT3 #(
    .INIT(8'h40)
  ) __147__ (
    .I2(G20),
    .I1(__10__),
    .I0(G4),
    .O(__67__)
  );
  LUT3 #(
    .INIT(8'hf7)
  ) __148__ (
    .I2(G4),
    .I1(__16__),
    .I0(G31),
    .O(__68__)
  );
  LUT4 #(
    .INIT(16'hff5d)
  ) __149__ (
    .I3(G4),
    .I2(__33__),
    .I1(__6__),
    .I0(__16__),
    .O(__69__)
  );
  LUT4 #(
    .INIT(16'h0040)
  ) __150__ (
    .I3(G4),
    .I2(__8__),
    .I1(__2__),
    .I0(__49__),
    .O(__70__)
  );
  LUT3 #(
    .INIT(8'h40)
  ) __151__ (
    .I2(__1__),
    .I1(__40__),
    .I0(G4),
    .O(__71__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __152__ (
    .I1(G10),
    .I0(G13),
    .O(__72__)
  );
  LUT6 #(
    .INIT(64'hbfff0000bfffbfff)
  ) __153__ (
    .I5(__72__),
    .I4(G9),
    .I3(__23__),
    .I2(__71__),
    .I1(__70__),
    .I0(G11),
    .O(__73__)
  );
  LUT6 #(
    .INIT(64'hff0fff55ff33ffff)
  ) __154__ (
    .I5(G9),
    .I4(G10),
    .I3(G13),
    .I2(__23__),
    .I1(__71__),
    .I0(__70__),
    .O(__74__)
  );
  LUT6 #(
    .INIT(64'hdf00000000000000)
  ) __155__ (
    .I5(G26),
    .I4(G12),
    .I3(__74__),
    .I2(__44__),
    .I1(__73__),
    .I0(__43__),
    .O(__75__)
  );
  LUT3 #(
    .INIT(8'h0b)
  ) __156__ (
    .I2(__29__),
    .I1(__5__),
    .I0(__27__),
    .O(__76__)
  );
  LUT6 #(
    .INIT(64'hffff404000ff0000)
  ) __157__ (
    .I5(G5),
    .I4(__31__),
    .I3(G2),
    .I2(__76__),
    .I1(__71__),
    .I0(__34__),
    .O(__77__)
  );
  LUT2 #(
    .INIT(4'h7)
  ) __158__ (
    .I1(G36),
    .I0(__23__),
    .O(__78__)
  );
  LUT3 #(
    .INIT(8'h40)
  ) __159__ (
    .I2(G18),
    .I1(__7__),
    .I0(G4),
    .O(__79__)
  );
  assign G83 = __64__;
  assign G89BF = __35__;
  assign G87BF = __19__;
  assign G91 = G27;
  assign G90 = __75__;
  assign G95BF = __53__;
  assign G105BF = __55__;
  assign G88BF = __49__;
  assign G98BF = __57__;
  assign G92 = __60__;
  assign G101BF = __78__;
  assign G104BF = __47__;
  assign G84 = __67__;
  assign G103BF = __48__;
  assign G99BF = __62__;
  assign G96BF = __68__;
  assign G86BF = __33__;
  assign G85 = __46__;
  assign G100BF = __21__;
  assign G107 = __79__;
  assign G97BF = __61__;
  assign G94 = G29;
  assign G106BF = __39__;
endmodule
