module alu_256(
  input wire a0, input wire b0,
  input wire a1, input wire b1,
  input wire a2, input wire b2,
  input wire a3, input wire b3,
  input wire a4, input wire b4,
  input wire a5, input wire b5,
  input wire a6, input wire b6,
  input wire a7, input wire b7,
  input wire a8, input wire b8,
  input wire a9, input wire b9,
  input wire a10, input wire b10,
  input wire a11, input wire b11,
  input wire a12, input wire b12,
  input wire a13, input wire b13,
  input wire a14, input wire b14,
  input wire a15, input wire b15,
  input wire a16, input wire b16,
  input wire a17, input wire b17,
  input wire a18, input wire b18,
  input wire a19, input wire b19,
  input wire a20, input wire b20,
  input wire a21, input wire b21,
  input wire a22, input wire b22,
  input wire a23, input wire b23,
  input wire a24, input wire b24,
  input wire a25, input wire b25,
  input wire a26, input wire b26,
  input wire a27, input wire b27,
  input wire a28, input wire b28,
  input wire a29, input wire b29,
  input wire a30, input wire b30,
  input wire a31, input wire b31,
  input wire a32, input wire b32,
  input wire a33, input wire b33,
  input wire a34, input wire b34,
  input wire a35, input wire b35,
  input wire a36, input wire b36,
  input wire a37, input wire b37,
  input wire a38, input wire b38,
  input wire a39, input wire b39,
  input wire a40, input wire b40,
  input wire a41, input wire b41,
  input wire a42, input wire b42,
  input wire a43, input wire b43,
  input wire a44, input wire b44,
  input wire a45, input wire b45,
  input wire a46, input wire b46,
  input wire a47, input wire b47,
  input wire a48, input wire b48,
  input wire a49, input wire b49,
  input wire a50, input wire b50,
  input wire a51, input wire b51,
  input wire a52, input wire b52,
  input wire a53, input wire b53,
  input wire a54, input wire b54,
  input wire a55, input wire b55,
  input wire a56, input wire b56,
  input wire a57, input wire b57,
  input wire a58, input wire b58,
  input wire a59, input wire b59,
  input wire a60, input wire b60,
  input wire a61, input wire b61,
  input wire a62, input wire b62,
  input wire a63, input wire b63,
  input wire a64, input wire b64,
  input wire a65, input wire b65,
  input wire a66, input wire b66,
  input wire a67, input wire b67,
  input wire a68, input wire b68,
  input wire a69, input wire b69,
  input wire a70, input wire b70,
  input wire a71, input wire b71,
  input wire a72, input wire b72,
  input wire a73, input wire b73,
  input wire a74, input wire b74,
  input wire a75, input wire b75,
  input wire a76, input wire b76,
  input wire a77, input wire b77,
  input wire a78, input wire b78,
  input wire a79, input wire b79,
  input wire a80, input wire b80,
  input wire a81, input wire b81,
  input wire a82, input wire b82,
  input wire a83, input wire b83,
  input wire a84, input wire b84,
  input wire a85, input wire b85,
  input wire a86, input wire b86,
  input wire a87, input wire b87,
  input wire a88, input wire b88,
  input wire a89, input wire b89,
  input wire a90, input wire b90,
  input wire a91, input wire b91,
  input wire a92, input wire b92,
  input wire a93, input wire b93,
  input wire a94, input wire b94,
  input wire a95, input wire b95,
  input wire a96, input wire b96,
  input wire a97, input wire b97,
  input wire a98, input wire b98,
  input wire a99, input wire b99,
  input wire a100, input wire b100,
  input wire a101, input wire b101,
  input wire a102, input wire b102,
  input wire a103, input wire b103,
  input wire a104, input wire b104,
  input wire a105, input wire b105,
  input wire a106, input wire b106,
  input wire a107, input wire b107,
  input wire a108, input wire b108,
  input wire a109, input wire b109,
  input wire a110, input wire b110,
  input wire a111, input wire b111,
  input wire a112, input wire b112,
  input wire a113, input wire b113,
  input wire a114, input wire b114,
  input wire a115, input wire b115,
  input wire a116, input wire b116,
  input wire a117, input wire b117,
  input wire a118, input wire b118,
  input wire a119, input wire b119,
  input wire a120, input wire b120,
  input wire a121, input wire b121,
  input wire a122, input wire b122,
  input wire a123, input wire b123,
  input wire a124, input wire b124,
  input wire a125, input wire b125,
  input wire a126, input wire b126,
  input wire a127, input wire b127,
  input wire a128, input wire b128,
  input wire a129, input wire b129,
  input wire a130, input wire b130,
  input wire a131, input wire b131,
  input wire a132, input wire b132,
  input wire a133, input wire b133,
  input wire a134, input wire b134,
  input wire a135, input wire b135,
  input wire a136, input wire b136,
  input wire a137, input wire b137,
  input wire a138, input wire b138,
  input wire a139, input wire b139,
  input wire a140, input wire b140,
  input wire a141, input wire b141,
  input wire a142, input wire b142,
  input wire a143, input wire b143,
  input wire a144, input wire b144,
  input wire a145, input wire b145,
  input wire a146, input wire b146,
  input wire a147, input wire b147,
  input wire a148, input wire b148,
  input wire a149, input wire b149,
  input wire a150, input wire b150,
  input wire a151, input wire b151,
  input wire a152, input wire b152,
  input wire a153, input wire b153,
  input wire a154, input wire b154,
  input wire a155, input wire b155,
  input wire a156, input wire b156,
  input wire a157, input wire b157,
  input wire a158, input wire b158,
  input wire a159, input wire b159,
  input wire a160, input wire b160,
  input wire a161, input wire b161,
  input wire a162, input wire b162,
  input wire a163, input wire b163,
  input wire a164, input wire b164,
  input wire a165, input wire b165,
  input wire a166, input wire b166,
  input wire a167, input wire b167,
  input wire a168, input wire b168,
  input wire a169, input wire b169,
  input wire a170, input wire b170,
  input wire a171, input wire b171,
  input wire a172, input wire b172,
  input wire a173, input wire b173,
  input wire a174, input wire b174,
  input wire a175, input wire b175,
  input wire a176, input wire b176,
  input wire a177, input wire b177,
  input wire a178, input wire b178,
  input wire a179, input wire b179,
  input wire a180, input wire b180,
  input wire a181, input wire b181,
  input wire a182, input wire b182,
  input wire a183, input wire b183,
  input wire a184, input wire b184,
  input wire a185, input wire b185,
  input wire a186, input wire b186,
  input wire a187, input wire b187,
  input wire a188, input wire b188,
  input wire a189, input wire b189,
  input wire a190, input wire b190,
  input wire a191, input wire b191,
  input wire a192, input wire b192,
  input wire a193, input wire b193,
  input wire a194, input wire b194,
  input wire a195, input wire b195,
  input wire a196, input wire b196,
  input wire a197, input wire b197,
  input wire a198, input wire b198,
  input wire a199, input wire b199,
  input wire a200, input wire b200,
  input wire a201, input wire b201,
  input wire a202, input wire b202,
  input wire a203, input wire b203,
  input wire a204, input wire b204,
  input wire a205, input wire b205,
  input wire a206, input wire b206,
  input wire a207, input wire b207,
  input wire a208, input wire b208,
  input wire a209, input wire b209,
  input wire a210, input wire b210,
  input wire a211, input wire b211,
  input wire a212, input wire b212,
  input wire a213, input wire b213,
  input wire a214, input wire b214,
  input wire a215, input wire b215,
  input wire a216, input wire b216,
  input wire a217, input wire b217,
  input wire a218, input wire b218,
  input wire a219, input wire b219,
  input wire a220, input wire b220,
  input wire a221, input wire b221,
  input wire a222, input wire b222,
  input wire a223, input wire b223,
  input wire a224, input wire b224,
  input wire a225, input wire b225,
  input wire a226, input wire b226,
  input wire a227, input wire b227,
  input wire a228, input wire b228,
  input wire a229, input wire b229,
  input wire a230, input wire b230,
  input wire a231, input wire b231,
  input wire a232, input wire b232,
  input wire a233, input wire b233,
  input wire a234, input wire b234,
  input wire a235, input wire b235,
  input wire a236, input wire b236,
  input wire a237, input wire b237,
  input wire a238, input wire b238,
  input wire a239, input wire b239,
  input wire a240, input wire b240,
  input wire a241, input wire b241,
  input wire a242, input wire b242,
  input wire a243, input wire b243,
  input wire a244, input wire b244,
  input wire a245, input wire b245,
  input wire a246, input wire b246,
  input wire a247, input wire b247,
  input wire a248, input wire b248,
  input wire a249, input wire b249,
  input wire a250, input wire b250,
  input wire a251, input wire b251,
  input wire a252, input wire b252,
  input wire a253, input wire b253,
  input wire a254, input wire b254,
  input wire a255, input wire b255,
  input wire op0,
  input wire op1,
  output wire y0,
  output wire y1,
  output wire y2,
  output wire y3,
  output wire y4,
  output wire y5,
  output wire y6,
  output wire y7,
  output wire y8,
  output wire y9,
  output wire y10,
  output wire y11,
  output wire y12,
  output wire y13,
  output wire y14,
  output wire y15,
  output wire y16,
  output wire y17,
  output wire y18,
  output wire y19,
  output wire y20,
  output wire y21,
  output wire y22,
  output wire y23,
  output wire y24,
  output wire y25,
  output wire y26,
  output wire y27,
  output wire y28,
  output wire y29,
  output wire y30,
  output wire y31,
  output wire y32,
  output wire y33,
  output wire y34,
  output wire y35,
  output wire y36,
  output wire y37,
  output wire y38,
  output wire y39,
  output wire y40,
  output wire y41,
  output wire y42,
  output wire y43,
  output wire y44,
  output wire y45,
  output wire y46,
  output wire y47,
  output wire y48,
  output wire y49,
  output wire y50,
  output wire y51,
  output wire y52,
  output wire y53,
  output wire y54,
  output wire y55,
  output wire y56,
  output wire y57,
  output wire y58,
  output wire y59,
  output wire y60,
  output wire y61,
  output wire y62,
  output wire y63,
  output wire y64,
  output wire y65,
  output wire y66,
  output wire y67,
  output wire y68,
  output wire y69,
  output wire y70,
  output wire y71,
  output wire y72,
  output wire y73,
  output wire y74,
  output wire y75,
  output wire y76,
  output wire y77,
  output wire y78,
  output wire y79,
  output wire y80,
  output wire y81,
  output wire y82,
  output wire y83,
  output wire y84,
  output wire y85,
  output wire y86,
  output wire y87,
  output wire y88,
  output wire y89,
  output wire y90,
  output wire y91,
  output wire y92,
  output wire y93,
  output wire y94,
  output wire y95,
  output wire y96,
  output wire y97,
  output wire y98,
  output wire y99,
  output wire y100,
  output wire y101,
  output wire y102,
  output wire y103,
  output wire y104,
  output wire y105,
  output wire y106,
  output wire y107,
  output wire y108,
  output wire y109,
  output wire y110,
  output wire y111,
  output wire y112,
  output wire y113,
  output wire y114,
  output wire y115,
  output wire y116,
  output wire y117,
  output wire y118,
  output wire y119,
  output wire y120,
  output wire y121,
  output wire y122,
  output wire y123,
  output wire y124,
  output wire y125,
  output wire y126,
  output wire y127,
  output wire y128,
  output wire y129,
  output wire y130,
  output wire y131,
  output wire y132,
  output wire y133,
  output wire y134,
  output wire y135,
  output wire y136,
  output wire y137,
  output wire y138,
  output wire y139,
  output wire y140,
  output wire y141,
  output wire y142,
  output wire y143,
  output wire y144,
  output wire y145,
  output wire y146,
  output wire y147,
  output wire y148,
  output wire y149,
  output wire y150,
  output wire y151,
  output wire y152,
  output wire y153,
  output wire y154,
  output wire y155,
  output wire y156,
  output wire y157,
  output wire y158,
  output wire y159,
  output wire y160,
  output wire y161,
  output wire y162,
  output wire y163,
  output wire y164,
  output wire y165,
  output wire y166,
  output wire y167,
  output wire y168,
  output wire y169,
  output wire y170,
  output wire y171,
  output wire y172,
  output wire y173,
  output wire y174,
  output wire y175,
  output wire y176,
  output wire y177,
  output wire y178,
  output wire y179,
  output wire y180,
  output wire y181,
  output wire y182,
  output wire y183,
  output wire y184,
  output wire y185,
  output wire y186,
  output wire y187,
  output wire y188,
  output wire y189,
  output wire y190,
  output wire y191,
  output wire y192,
  output wire y193,
  output wire y194,
  output wire y195,
  output wire y196,
  output wire y197,
  output wire y198,
  output wire y199,
  output wire y200,
  output wire y201,
  output wire y202,
  output wire y203,
  output wire y204,
  output wire y205,
  output wire y206,
  output wire y207,
  output wire y208,
  output wire y209,
  output wire y210,
  output wire y211,
  output wire y212,
  output wire y213,
  output wire y214,
  output wire y215,
  output wire y216,
  output wire y217,
  output wire y218,
  output wire y219,
  output wire y220,
  output wire y221,
  output wire y222,
  output wire y223,
  output wire y224,
  output wire y225,
  output wire y226,
  output wire y227,
  output wire y228,
  output wire y229,
  output wire y230,
  output wire y231,
  output wire y232,
  output wire y233,
  output wire y234,
  output wire y235,
  output wire y236,
  output wire y237,
  output wire y238,
  output wire y239,
  output wire y240,
  output wire y241,
  output wire y242,
  output wire y243,
  output wire y244,
  output wire y245,
  output wire y246,
  output wire y247,
  output wire y248,
  output wire y249,
  output wire y250,
  output wire y251,
  output wire y252,
  output wire y253,
  output wire y254,
  output wire y255
);
  wire add_sel, sub_sel, and_sel, or_sel;
  assign add_sel = ~op1 & ~op0;
  assign sub_sel = ~op1 & op0;
  assign and_sel = op1 & ~op0;
  assign or_sel  = op1 & op0;
  wire c0;
  wire c1;
  wire c2;
  wire c3;
  wire c4;
  wire c5;
  wire c6;
  wire c7;
  wire c8;
  wire c9;
  wire c10;
  wire c11;
  wire c12;
  wire c13;
  wire c14;
  wire c15;
  wire c16;
  wire c17;
  wire c18;
  wire c19;
  wire c20;
  wire c21;
  wire c22;
  wire c23;
  wire c24;
  wire c25;
  wire c26;
  wire c27;
  wire c28;
  wire c29;
  wire c30;
  wire c31;
  wire c32;
  wire c33;
  wire c34;
  wire c35;
  wire c36;
  wire c37;
  wire c38;
  wire c39;
  wire c40;
  wire c41;
  wire c42;
  wire c43;
  wire c44;
  wire c45;
  wire c46;
  wire c47;
  wire c48;
  wire c49;
  wire c50;
  wire c51;
  wire c52;
  wire c53;
  wire c54;
  wire c55;
  wire c56;
  wire c57;
  wire c58;
  wire c59;
  wire c60;
  wire c61;
  wire c62;
  wire c63;
  wire c64;
  wire c65;
  wire c66;
  wire c67;
  wire c68;
  wire c69;
  wire c70;
  wire c71;
  wire c72;
  wire c73;
  wire c74;
  wire c75;
  wire c76;
  wire c77;
  wire c78;
  wire c79;
  wire c80;
  wire c81;
  wire c82;
  wire c83;
  wire c84;
  wire c85;
  wire c86;
  wire c87;
  wire c88;
  wire c89;
  wire c90;
  wire c91;
  wire c92;
  wire c93;
  wire c94;
  wire c95;
  wire c96;
  wire c97;
  wire c98;
  wire c99;
  wire c100;
  wire c101;
  wire c102;
  wire c103;
  wire c104;
  wire c105;
  wire c106;
  wire c107;
  wire c108;
  wire c109;
  wire c110;
  wire c111;
  wire c112;
  wire c113;
  wire c114;
  wire c115;
  wire c116;
  wire c117;
  wire c118;
  wire c119;
  wire c120;
  wire c121;
  wire c122;
  wire c123;
  wire c124;
  wire c125;
  wire c126;
  wire c127;
  wire c128;
  wire c129;
  wire c130;
  wire c131;
  wire c132;
  wire c133;
  wire c134;
  wire c135;
  wire c136;
  wire c137;
  wire c138;
  wire c139;
  wire c140;
  wire c141;
  wire c142;
  wire c143;
  wire c144;
  wire c145;
  wire c146;
  wire c147;
  wire c148;
  wire c149;
  wire c150;
  wire c151;
  wire c152;
  wire c153;
  wire c154;
  wire c155;
  wire c156;
  wire c157;
  wire c158;
  wire c159;
  wire c160;
  wire c161;
  wire c162;
  wire c163;
  wire c164;
  wire c165;
  wire c166;
  wire c167;
  wire c168;
  wire c169;
  wire c170;
  wire c171;
  wire c172;
  wire c173;
  wire c174;
  wire c175;
  wire c176;
  wire c177;
  wire c178;
  wire c179;
  wire c180;
  wire c181;
  wire c182;
  wire c183;
  wire c184;
  wire c185;
  wire c186;
  wire c187;
  wire c188;
  wire c189;
  wire c190;
  wire c191;
  wire c192;
  wire c193;
  wire c194;
  wire c195;
  wire c196;
  wire c197;
  wire c198;
  wire c199;
  wire c200;
  wire c201;
  wire c202;
  wire c203;
  wire c204;
  wire c205;
  wire c206;
  wire c207;
  wire c208;
  wire c209;
  wire c210;
  wire c211;
  wire c212;
  wire c213;
  wire c214;
  wire c215;
  wire c216;
  wire c217;
  wire c218;
  wire c219;
  wire c220;
  wire c221;
  wire c222;
  wire c223;
  wire c224;
  wire c225;
  wire c226;
  wire c227;
  wire c228;
  wire c229;
  wire c230;
  wire c231;
  wire c232;
  wire c233;
  wire c234;
  wire c235;
  wire c236;
  wire c237;
  wire c238;
  wire c239;
  wire c240;
  wire c241;
  wire c242;
  wire c243;
  wire c244;
  wire c245;
  wire c246;
  wire c247;
  wire c248;
  wire c249;
  wire c250;
  wire c251;
  wire c252;
  wire c253;
  wire c254;
  wire c255;
  wire c256;
  assign c0 = 1'b0;
  wire s0, sub0, and0, or0;
  wire b_inv0;
  assign b_inv0 = ~b0;
  assign s0  = a0 ^ b0 ^ c0;
  assign sub0 = a0 ^ b_inv0 ^ c0;
  assign and0 = a0 & b0;
  assign or0  = a0 | b0;
  assign c1 = (a0 & b0) | (a0 & c0) | (b0 & c0);
  wire c_sub1;
  assign c_sub1 = (a0 & b_inv0) | (a0 & c0) | (b_inv0 & c0);
  wire s1, sub1, and1, or1;
  wire b_inv1;
  assign b_inv1 = ~b1;
  assign s1  = a1 ^ b1 ^ c1;
  assign sub1 = a1 ^ b_inv1 ^ c1;
  assign and1 = a1 & b1;
  assign or1  = a1 | b1;
  assign c2 = (a1 & b1) | (a1 & c1) | (b1 & c1);
  wire c_sub2;
  assign c_sub2 = (a1 & b_inv1) | (a1 & c1) | (b_inv1 & c1);
  wire s2, sub2, and2, or2;
  wire b_inv2;
  assign b_inv2 = ~b2;
  assign s2  = a2 ^ b2 ^ c2;
  assign sub2 = a2 ^ b_inv2 ^ c2;
  assign and2 = a2 & b2;
  assign or2  = a2 | b2;
  assign c3 = (a2 & b2) | (a2 & c2) | (b2 & c2);
  wire c_sub3;
  assign c_sub3 = (a2 & b_inv2) | (a2 & c2) | (b_inv2 & c2);
  wire s3, sub3, and3, or3;
  wire b_inv3;
  assign b_inv3 = ~b3;
  assign s3  = a3 ^ b3 ^ c3;
  assign sub3 = a3 ^ b_inv3 ^ c3;
  assign and3 = a3 & b3;
  assign or3  = a3 | b3;
  assign c4 = (a3 & b3) | (a3 & c3) | (b3 & c3);
  wire c_sub4;
  assign c_sub4 = (a3 & b_inv3) | (a3 & c3) | (b_inv3 & c3);
  wire s4, sub4, and4, or4;
  wire b_inv4;
  assign b_inv4 = ~b4;
  assign s4  = a4 ^ b4 ^ c4;
  assign sub4 = a4 ^ b_inv4 ^ c4;
  assign and4 = a4 & b4;
  assign or4  = a4 | b4;
  assign c5 = (a4 & b4) | (a4 & c4) | (b4 & c4);
  wire c_sub5;
  assign c_sub5 = (a4 & b_inv4) | (a4 & c4) | (b_inv4 & c4);
  wire s5, sub5, and5, or5;
  wire b_inv5;
  assign b_inv5 = ~b5;
  assign s5  = a5 ^ b5 ^ c5;
  assign sub5 = a5 ^ b_inv5 ^ c5;
  assign and5 = a5 & b5;
  assign or5  = a5 | b5;
  assign c6 = (a5 & b5) | (a5 & c5) | (b5 & c5);
  wire c_sub6;
  assign c_sub6 = (a5 & b_inv5) | (a5 & c5) | (b_inv5 & c5);
  wire s6, sub6, and6, or6;
  wire b_inv6;
  assign b_inv6 = ~b6;
  assign s6  = a6 ^ b6 ^ c6;
  assign sub6 = a6 ^ b_inv6 ^ c6;
  assign and6 = a6 & b6;
  assign or6  = a6 | b6;
  assign c7 = (a6 & b6) | (a6 & c6) | (b6 & c6);
  wire c_sub7;
  assign c_sub7 = (a6 & b_inv6) | (a6 & c6) | (b_inv6 & c6);
  wire s7, sub7, and7, or7;
  wire b_inv7;
  assign b_inv7 = ~b7;
  assign s7  = a7 ^ b7 ^ c7;
  assign sub7 = a7 ^ b_inv7 ^ c7;
  assign and7 = a7 & b7;
  assign or7  = a7 | b7;
  assign c8 = (a7 & b7) | (a7 & c7) | (b7 & c7);
  wire c_sub8;
  assign c_sub8 = (a7 & b_inv7) | (a7 & c7) | (b_inv7 & c7);
  wire s8, sub8, and8, or8;
  wire b_inv8;
  assign b_inv8 = ~b8;
  assign s8  = a8 ^ b8 ^ c8;
  assign sub8 = a8 ^ b_inv8 ^ c8;
  assign and8 = a8 & b8;
  assign or8  = a8 | b8;
  assign c9 = (a8 & b8) | (a8 & c8) | (b8 & c8);
  wire c_sub9;
  assign c_sub9 = (a8 & b_inv8) | (a8 & c8) | (b_inv8 & c8);
  wire s9, sub9, and9, or9;
  wire b_inv9;
  assign b_inv9 = ~b9;
  assign s9  = a9 ^ b9 ^ c9;
  assign sub9 = a9 ^ b_inv9 ^ c9;
  assign and9 = a9 & b9;
  assign or9  = a9 | b9;
  assign c10 = (a9 & b9) | (a9 & c9) | (b9 & c9);
  wire c_sub10;
  assign c_sub10 = (a9 & b_inv9) | (a9 & c9) | (b_inv9 & c9);
  wire s10, sub10, and10, or10;
  wire b_inv10;
  assign b_inv10 = ~b10;
  assign s10  = a10 ^ b10 ^ c10;
  assign sub10 = a10 ^ b_inv10 ^ c10;
  assign and10 = a10 & b10;
  assign or10  = a10 | b10;
  assign c11 = (a10 & b10) | (a10 & c10) | (b10 & c10);
  wire c_sub11;
  assign c_sub11 = (a10 & b_inv10) | (a10 & c10) | (b_inv10 & c10);
  wire s11, sub11, and11, or11;
  wire b_inv11;
  assign b_inv11 = ~b11;
  assign s11  = a11 ^ b11 ^ c11;
  assign sub11 = a11 ^ b_inv11 ^ c11;
  assign and11 = a11 & b11;
  assign or11  = a11 | b11;
  assign c12 = (a11 & b11) | (a11 & c11) | (b11 & c11);
  wire c_sub12;
  assign c_sub12 = (a11 & b_inv11) | (a11 & c11) | (b_inv11 & c11);
  wire s12, sub12, and12, or12;
  wire b_inv12;
  assign b_inv12 = ~b12;
  assign s12  = a12 ^ b12 ^ c12;
  assign sub12 = a12 ^ b_inv12 ^ c12;
  assign and12 = a12 & b12;
  assign or12  = a12 | b12;
  assign c13 = (a12 & b12) | (a12 & c12) | (b12 & c12);
  wire c_sub13;
  assign c_sub13 = (a12 & b_inv12) | (a12 & c12) | (b_inv12 & c12);
  wire s13, sub13, and13, or13;
  wire b_inv13;
  assign b_inv13 = ~b13;
  assign s13  = a13 ^ b13 ^ c13;
  assign sub13 = a13 ^ b_inv13 ^ c13;
  assign and13 = a13 & b13;
  assign or13  = a13 | b13;
  assign c14 = (a13 & b13) | (a13 & c13) | (b13 & c13);
  wire c_sub14;
  assign c_sub14 = (a13 & b_inv13) | (a13 & c13) | (b_inv13 & c13);
  wire s14, sub14, and14, or14;
  wire b_inv14;
  assign b_inv14 = ~b14;
  assign s14  = a14 ^ b14 ^ c14;
  assign sub14 = a14 ^ b_inv14 ^ c14;
  assign and14 = a14 & b14;
  assign or14  = a14 | b14;
  assign c15 = (a14 & b14) | (a14 & c14) | (b14 & c14);
  wire c_sub15;
  assign c_sub15 = (a14 & b_inv14) | (a14 & c14) | (b_inv14 & c14);
  wire s15, sub15, and15, or15;
  wire b_inv15;
  assign b_inv15 = ~b15;
  assign s15  = a15 ^ b15 ^ c15;
  assign sub15 = a15 ^ b_inv15 ^ c15;
  assign and15 = a15 & b15;
  assign or15  = a15 | b15;
  assign c16 = (a15 & b15) | (a15 & c15) | (b15 & c15);
  wire c_sub16;
  assign c_sub16 = (a15 & b_inv15) | (a15 & c15) | (b_inv15 & c15);
  wire s16, sub16, and16, or16;
  wire b_inv16;
  assign b_inv16 = ~b16;
  assign s16  = a16 ^ b16 ^ c16;
  assign sub16 = a16 ^ b_inv16 ^ c16;
  assign and16 = a16 & b16;
  assign or16  = a16 | b16;
  assign c17 = (a16 & b16) | (a16 & c16) | (b16 & c16);
  wire c_sub17;
  assign c_sub17 = (a16 & b_inv16) | (a16 & c16) | (b_inv16 & c16);
  wire s17, sub17, and17, or17;
  wire b_inv17;
  assign b_inv17 = ~b17;
  assign s17  = a17 ^ b17 ^ c17;
  assign sub17 = a17 ^ b_inv17 ^ c17;
  assign and17 = a17 & b17;
  assign or17  = a17 | b17;
  assign c18 = (a17 & b17) | (a17 & c17) | (b17 & c17);
  wire c_sub18;
  assign c_sub18 = (a17 & b_inv17) | (a17 & c17) | (b_inv17 & c17);
  wire s18, sub18, and18, or18;
  wire b_inv18;
  assign b_inv18 = ~b18;
  assign s18  = a18 ^ b18 ^ c18;
  assign sub18 = a18 ^ b_inv18 ^ c18;
  assign and18 = a18 & b18;
  assign or18  = a18 | b18;
  assign c19 = (a18 & b18) | (a18 & c18) | (b18 & c18);
  wire c_sub19;
  assign c_sub19 = (a18 & b_inv18) | (a18 & c18) | (b_inv18 & c18);
  wire s19, sub19, and19, or19;
  wire b_inv19;
  assign b_inv19 = ~b19;
  assign s19  = a19 ^ b19 ^ c19;
  assign sub19 = a19 ^ b_inv19 ^ c19;
  assign and19 = a19 & b19;
  assign or19  = a19 | b19;
  assign c20 = (a19 & b19) | (a19 & c19) | (b19 & c19);
  wire c_sub20;
  assign c_sub20 = (a19 & b_inv19) | (a19 & c19) | (b_inv19 & c19);
  wire s20, sub20, and20, or20;
  wire b_inv20;
  assign b_inv20 = ~b20;
  assign s20  = a20 ^ b20 ^ c20;
  assign sub20 = a20 ^ b_inv20 ^ c20;
  assign and20 = a20 & b20;
  assign or20  = a20 | b20;
  assign c21 = (a20 & b20) | (a20 & c20) | (b20 & c20);
  wire c_sub21;
  assign c_sub21 = (a20 & b_inv20) | (a20 & c20) | (b_inv20 & c20);
  wire s21, sub21, and21, or21;
  wire b_inv21;
  assign b_inv21 = ~b21;
  assign s21  = a21 ^ b21 ^ c21;
  assign sub21 = a21 ^ b_inv21 ^ c21;
  assign and21 = a21 & b21;
  assign or21  = a21 | b21;
  assign c22 = (a21 & b21) | (a21 & c21) | (b21 & c21);
  wire c_sub22;
  assign c_sub22 = (a21 & b_inv21) | (a21 & c21) | (b_inv21 & c21);
  wire s22, sub22, and22, or22;
  wire b_inv22;
  assign b_inv22 = ~b22;
  assign s22  = a22 ^ b22 ^ c22;
  assign sub22 = a22 ^ b_inv22 ^ c22;
  assign and22 = a22 & b22;
  assign or22  = a22 | b22;
  assign c23 = (a22 & b22) | (a22 & c22) | (b22 & c22);
  wire c_sub23;
  assign c_sub23 = (a22 & b_inv22) | (a22 & c22) | (b_inv22 & c22);
  wire s23, sub23, and23, or23;
  wire b_inv23;
  assign b_inv23 = ~b23;
  assign s23  = a23 ^ b23 ^ c23;
  assign sub23 = a23 ^ b_inv23 ^ c23;
  assign and23 = a23 & b23;
  assign or23  = a23 | b23;
  assign c24 = (a23 & b23) | (a23 & c23) | (b23 & c23);
  wire c_sub24;
  assign c_sub24 = (a23 & b_inv23) | (a23 & c23) | (b_inv23 & c23);
  wire s24, sub24, and24, or24;
  wire b_inv24;
  assign b_inv24 = ~b24;
  assign s24  = a24 ^ b24 ^ c24;
  assign sub24 = a24 ^ b_inv24 ^ c24;
  assign and24 = a24 & b24;
  assign or24  = a24 | b24;
  assign c25 = (a24 & b24) | (a24 & c24) | (b24 & c24);
  wire c_sub25;
  assign c_sub25 = (a24 & b_inv24) | (a24 & c24) | (b_inv24 & c24);
  wire s25, sub25, and25, or25;
  wire b_inv25;
  assign b_inv25 = ~b25;
  assign s25  = a25 ^ b25 ^ c25;
  assign sub25 = a25 ^ b_inv25 ^ c25;
  assign and25 = a25 & b25;
  assign or25  = a25 | b25;
  assign c26 = (a25 & b25) | (a25 & c25) | (b25 & c25);
  wire c_sub26;
  assign c_sub26 = (a25 & b_inv25) | (a25 & c25) | (b_inv25 & c25);
  wire s26, sub26, and26, or26;
  wire b_inv26;
  assign b_inv26 = ~b26;
  assign s26  = a26 ^ b26 ^ c26;
  assign sub26 = a26 ^ b_inv26 ^ c26;
  assign and26 = a26 & b26;
  assign or26  = a26 | b26;
  assign c27 = (a26 & b26) | (a26 & c26) | (b26 & c26);
  wire c_sub27;
  assign c_sub27 = (a26 & b_inv26) | (a26 & c26) | (b_inv26 & c26);
  wire s27, sub27, and27, or27;
  wire b_inv27;
  assign b_inv27 = ~b27;
  assign s27  = a27 ^ b27 ^ c27;
  assign sub27 = a27 ^ b_inv27 ^ c27;
  assign and27 = a27 & b27;
  assign or27  = a27 | b27;
  assign c28 = (a27 & b27) | (a27 & c27) | (b27 & c27);
  wire c_sub28;
  assign c_sub28 = (a27 & b_inv27) | (a27 & c27) | (b_inv27 & c27);
  wire s28, sub28, and28, or28;
  wire b_inv28;
  assign b_inv28 = ~b28;
  assign s28  = a28 ^ b28 ^ c28;
  assign sub28 = a28 ^ b_inv28 ^ c28;
  assign and28 = a28 & b28;
  assign or28  = a28 | b28;
  assign c29 = (a28 & b28) | (a28 & c28) | (b28 & c28);
  wire c_sub29;
  assign c_sub29 = (a28 & b_inv28) | (a28 & c28) | (b_inv28 & c28);
  wire s29, sub29, and29, or29;
  wire b_inv29;
  assign b_inv29 = ~b29;
  assign s29  = a29 ^ b29 ^ c29;
  assign sub29 = a29 ^ b_inv29 ^ c29;
  assign and29 = a29 & b29;
  assign or29  = a29 | b29;
  assign c30 = (a29 & b29) | (a29 & c29) | (b29 & c29);
  wire c_sub30;
  assign c_sub30 = (a29 & b_inv29) | (a29 & c29) | (b_inv29 & c29);
  wire s30, sub30, and30, or30;
  wire b_inv30;
  assign b_inv30 = ~b30;
  assign s30  = a30 ^ b30 ^ c30;
  assign sub30 = a30 ^ b_inv30 ^ c30;
  assign and30 = a30 & b30;
  assign or30  = a30 | b30;
  assign c31 = (a30 & b30) | (a30 & c30) | (b30 & c30);
  wire c_sub31;
  assign c_sub31 = (a30 & b_inv30) | (a30 & c30) | (b_inv30 & c30);
  wire s31, sub31, and31, or31;
  wire b_inv31;
  assign b_inv31 = ~b31;
  assign s31  = a31 ^ b31 ^ c31;
  assign sub31 = a31 ^ b_inv31 ^ c31;
  assign and31 = a31 & b31;
  assign or31  = a31 | b31;
  assign c32 = (a31 & b31) | (a31 & c31) | (b31 & c31);
  wire c_sub32;
  assign c_sub32 = (a31 & b_inv31) | (a31 & c31) | (b_inv31 & c31);
  wire s32, sub32, and32, or32;
  wire b_inv32;
  assign b_inv32 = ~b32;
  assign s32  = a32 ^ b32 ^ c32;
  assign sub32 = a32 ^ b_inv32 ^ c32;
  assign and32 = a32 & b32;
  assign or32  = a32 | b32;
  assign c33 = (a32 & b32) | (a32 & c32) | (b32 & c32);
  wire c_sub33;
  assign c_sub33 = (a32 & b_inv32) | (a32 & c32) | (b_inv32 & c32);
  wire s33, sub33, and33, or33;
  wire b_inv33;
  assign b_inv33 = ~b33;
  assign s33  = a33 ^ b33 ^ c33;
  assign sub33 = a33 ^ b_inv33 ^ c33;
  assign and33 = a33 & b33;
  assign or33  = a33 | b33;
  assign c34 = (a33 & b33) | (a33 & c33) | (b33 & c33);
  wire c_sub34;
  assign c_sub34 = (a33 & b_inv33) | (a33 & c33) | (b_inv33 & c33);
  wire s34, sub34, and34, or34;
  wire b_inv34;
  assign b_inv34 = ~b34;
  assign s34  = a34 ^ b34 ^ c34;
  assign sub34 = a34 ^ b_inv34 ^ c34;
  assign and34 = a34 & b34;
  assign or34  = a34 | b34;
  assign c35 = (a34 & b34) | (a34 & c34) | (b34 & c34);
  wire c_sub35;
  assign c_sub35 = (a34 & b_inv34) | (a34 & c34) | (b_inv34 & c34);
  wire s35, sub35, and35, or35;
  wire b_inv35;
  assign b_inv35 = ~b35;
  assign s35  = a35 ^ b35 ^ c35;
  assign sub35 = a35 ^ b_inv35 ^ c35;
  assign and35 = a35 & b35;
  assign or35  = a35 | b35;
  assign c36 = (a35 & b35) | (a35 & c35) | (b35 & c35);
  wire c_sub36;
  assign c_sub36 = (a35 & b_inv35) | (a35 & c35) | (b_inv35 & c35);
  wire s36, sub36, and36, or36;
  wire b_inv36;
  assign b_inv36 = ~b36;
  assign s36  = a36 ^ b36 ^ c36;
  assign sub36 = a36 ^ b_inv36 ^ c36;
  assign and36 = a36 & b36;
  assign or36  = a36 | b36;
  assign c37 = (a36 & b36) | (a36 & c36) | (b36 & c36);
  wire c_sub37;
  assign c_sub37 = (a36 & b_inv36) | (a36 & c36) | (b_inv36 & c36);
  wire s37, sub37, and37, or37;
  wire b_inv37;
  assign b_inv37 = ~b37;
  assign s37  = a37 ^ b37 ^ c37;
  assign sub37 = a37 ^ b_inv37 ^ c37;
  assign and37 = a37 & b37;
  assign or37  = a37 | b37;
  assign c38 = (a37 & b37) | (a37 & c37) | (b37 & c37);
  wire c_sub38;
  assign c_sub38 = (a37 & b_inv37) | (a37 & c37) | (b_inv37 & c37);
  wire s38, sub38, and38, or38;
  wire b_inv38;
  assign b_inv38 = ~b38;
  assign s38  = a38 ^ b38 ^ c38;
  assign sub38 = a38 ^ b_inv38 ^ c38;
  assign and38 = a38 & b38;
  assign or38  = a38 | b38;
  assign c39 = (a38 & b38) | (a38 & c38) | (b38 & c38);
  wire c_sub39;
  assign c_sub39 = (a38 & b_inv38) | (a38 & c38) | (b_inv38 & c38);
  wire s39, sub39, and39, or39;
  wire b_inv39;
  assign b_inv39 = ~b39;
  assign s39  = a39 ^ b39 ^ c39;
  assign sub39 = a39 ^ b_inv39 ^ c39;
  assign and39 = a39 & b39;
  assign or39  = a39 | b39;
  assign c40 = (a39 & b39) | (a39 & c39) | (b39 & c39);
  wire c_sub40;
  assign c_sub40 = (a39 & b_inv39) | (a39 & c39) | (b_inv39 & c39);
  wire s40, sub40, and40, or40;
  wire b_inv40;
  assign b_inv40 = ~b40;
  assign s40  = a40 ^ b40 ^ c40;
  assign sub40 = a40 ^ b_inv40 ^ c40;
  assign and40 = a40 & b40;
  assign or40  = a40 | b40;
  assign c41 = (a40 & b40) | (a40 & c40) | (b40 & c40);
  wire c_sub41;
  assign c_sub41 = (a40 & b_inv40) | (a40 & c40) | (b_inv40 & c40);
  wire s41, sub41, and41, or41;
  wire b_inv41;
  assign b_inv41 = ~b41;
  assign s41  = a41 ^ b41 ^ c41;
  assign sub41 = a41 ^ b_inv41 ^ c41;
  assign and41 = a41 & b41;
  assign or41  = a41 | b41;
  assign c42 = (a41 & b41) | (a41 & c41) | (b41 & c41);
  wire c_sub42;
  assign c_sub42 = (a41 & b_inv41) | (a41 & c41) | (b_inv41 & c41);
  wire s42, sub42, and42, or42;
  wire b_inv42;
  assign b_inv42 = ~b42;
  assign s42  = a42 ^ b42 ^ c42;
  assign sub42 = a42 ^ b_inv42 ^ c42;
  assign and42 = a42 & b42;
  assign or42  = a42 | b42;
  assign c43 = (a42 & b42) | (a42 & c42) | (b42 & c42);
  wire c_sub43;
  assign c_sub43 = (a42 & b_inv42) | (a42 & c42) | (b_inv42 & c42);
  wire s43, sub43, and43, or43;
  wire b_inv43;
  assign b_inv43 = ~b43;
  assign s43  = a43 ^ b43 ^ c43;
  assign sub43 = a43 ^ b_inv43 ^ c43;
  assign and43 = a43 & b43;
  assign or43  = a43 | b43;
  assign c44 = (a43 & b43) | (a43 & c43) | (b43 & c43);
  wire c_sub44;
  assign c_sub44 = (a43 & b_inv43) | (a43 & c43) | (b_inv43 & c43);
  wire s44, sub44, and44, or44;
  wire b_inv44;
  assign b_inv44 = ~b44;
  assign s44  = a44 ^ b44 ^ c44;
  assign sub44 = a44 ^ b_inv44 ^ c44;
  assign and44 = a44 & b44;
  assign or44  = a44 | b44;
  assign c45 = (a44 & b44) | (a44 & c44) | (b44 & c44);
  wire c_sub45;
  assign c_sub45 = (a44 & b_inv44) | (a44 & c44) | (b_inv44 & c44);
  wire s45, sub45, and45, or45;
  wire b_inv45;
  assign b_inv45 = ~b45;
  assign s45  = a45 ^ b45 ^ c45;
  assign sub45 = a45 ^ b_inv45 ^ c45;
  assign and45 = a45 & b45;
  assign or45  = a45 | b45;
  assign c46 = (a45 & b45) | (a45 & c45) | (b45 & c45);
  wire c_sub46;
  assign c_sub46 = (a45 & b_inv45) | (a45 & c45) | (b_inv45 & c45);
  wire s46, sub46, and46, or46;
  wire b_inv46;
  assign b_inv46 = ~b46;
  assign s46  = a46 ^ b46 ^ c46;
  assign sub46 = a46 ^ b_inv46 ^ c46;
  assign and46 = a46 & b46;
  assign or46  = a46 | b46;
  assign c47 = (a46 & b46) | (a46 & c46) | (b46 & c46);
  wire c_sub47;
  assign c_sub47 = (a46 & b_inv46) | (a46 & c46) | (b_inv46 & c46);
  wire s47, sub47, and47, or47;
  wire b_inv47;
  assign b_inv47 = ~b47;
  assign s47  = a47 ^ b47 ^ c47;
  assign sub47 = a47 ^ b_inv47 ^ c47;
  assign and47 = a47 & b47;
  assign or47  = a47 | b47;
  assign c48 = (a47 & b47) | (a47 & c47) | (b47 & c47);
  wire c_sub48;
  assign c_sub48 = (a47 & b_inv47) | (a47 & c47) | (b_inv47 & c47);
  wire s48, sub48, and48, or48;
  wire b_inv48;
  assign b_inv48 = ~b48;
  assign s48  = a48 ^ b48 ^ c48;
  assign sub48 = a48 ^ b_inv48 ^ c48;
  assign and48 = a48 & b48;
  assign or48  = a48 | b48;
  assign c49 = (a48 & b48) | (a48 & c48) | (b48 & c48);
  wire c_sub49;
  assign c_sub49 = (a48 & b_inv48) | (a48 & c48) | (b_inv48 & c48);
  wire s49, sub49, and49, or49;
  wire b_inv49;
  assign b_inv49 = ~b49;
  assign s49  = a49 ^ b49 ^ c49;
  assign sub49 = a49 ^ b_inv49 ^ c49;
  assign and49 = a49 & b49;
  assign or49  = a49 | b49;
  assign c50 = (a49 & b49) | (a49 & c49) | (b49 & c49);
  wire c_sub50;
  assign c_sub50 = (a49 & b_inv49) | (a49 & c49) | (b_inv49 & c49);
  wire s50, sub50, and50, or50;
  wire b_inv50;
  assign b_inv50 = ~b50;
  assign s50  = a50 ^ b50 ^ c50;
  assign sub50 = a50 ^ b_inv50 ^ c50;
  assign and50 = a50 & b50;
  assign or50  = a50 | b50;
  assign c51 = (a50 & b50) | (a50 & c50) | (b50 & c50);
  wire c_sub51;
  assign c_sub51 = (a50 & b_inv50) | (a50 & c50) | (b_inv50 & c50);
  wire s51, sub51, and51, or51;
  wire b_inv51;
  assign b_inv51 = ~b51;
  assign s51  = a51 ^ b51 ^ c51;
  assign sub51 = a51 ^ b_inv51 ^ c51;
  assign and51 = a51 & b51;
  assign or51  = a51 | b51;
  assign c52 = (a51 & b51) | (a51 & c51) | (b51 & c51);
  wire c_sub52;
  assign c_sub52 = (a51 & b_inv51) | (a51 & c51) | (b_inv51 & c51);
  wire s52, sub52, and52, or52;
  wire b_inv52;
  assign b_inv52 = ~b52;
  assign s52  = a52 ^ b52 ^ c52;
  assign sub52 = a52 ^ b_inv52 ^ c52;
  assign and52 = a52 & b52;
  assign or52  = a52 | b52;
  assign c53 = (a52 & b52) | (a52 & c52) | (b52 & c52);
  wire c_sub53;
  assign c_sub53 = (a52 & b_inv52) | (a52 & c52) | (b_inv52 & c52);
  wire s53, sub53, and53, or53;
  wire b_inv53;
  assign b_inv53 = ~b53;
  assign s53  = a53 ^ b53 ^ c53;
  assign sub53 = a53 ^ b_inv53 ^ c53;
  assign and53 = a53 & b53;
  assign or53  = a53 | b53;
  assign c54 = (a53 & b53) | (a53 & c53) | (b53 & c53);
  wire c_sub54;
  assign c_sub54 = (a53 & b_inv53) | (a53 & c53) | (b_inv53 & c53);
  wire s54, sub54, and54, or54;
  wire b_inv54;
  assign b_inv54 = ~b54;
  assign s54  = a54 ^ b54 ^ c54;
  assign sub54 = a54 ^ b_inv54 ^ c54;
  assign and54 = a54 & b54;
  assign or54  = a54 | b54;
  assign c55 = (a54 & b54) | (a54 & c54) | (b54 & c54);
  wire c_sub55;
  assign c_sub55 = (a54 & b_inv54) | (a54 & c54) | (b_inv54 & c54);
  wire s55, sub55, and55, or55;
  wire b_inv55;
  assign b_inv55 = ~b55;
  assign s55  = a55 ^ b55 ^ c55;
  assign sub55 = a55 ^ b_inv55 ^ c55;
  assign and55 = a55 & b55;
  assign or55  = a55 | b55;
  assign c56 = (a55 & b55) | (a55 & c55) | (b55 & c55);
  wire c_sub56;
  assign c_sub56 = (a55 & b_inv55) | (a55 & c55) | (b_inv55 & c55);
  wire s56, sub56, and56, or56;
  wire b_inv56;
  assign b_inv56 = ~b56;
  assign s56  = a56 ^ b56 ^ c56;
  assign sub56 = a56 ^ b_inv56 ^ c56;
  assign and56 = a56 & b56;
  assign or56  = a56 | b56;
  assign c57 = (a56 & b56) | (a56 & c56) | (b56 & c56);
  wire c_sub57;
  assign c_sub57 = (a56 & b_inv56) | (a56 & c56) | (b_inv56 & c56);
  wire s57, sub57, and57, or57;
  wire b_inv57;
  assign b_inv57 = ~b57;
  assign s57  = a57 ^ b57 ^ c57;
  assign sub57 = a57 ^ b_inv57 ^ c57;
  assign and57 = a57 & b57;
  assign or57  = a57 | b57;
  assign c58 = (a57 & b57) | (a57 & c57) | (b57 & c57);
  wire c_sub58;
  assign c_sub58 = (a57 & b_inv57) | (a57 & c57) | (b_inv57 & c57);
  wire s58, sub58, and58, or58;
  wire b_inv58;
  assign b_inv58 = ~b58;
  assign s58  = a58 ^ b58 ^ c58;
  assign sub58 = a58 ^ b_inv58 ^ c58;
  assign and58 = a58 & b58;
  assign or58  = a58 | b58;
  assign c59 = (a58 & b58) | (a58 & c58) | (b58 & c58);
  wire c_sub59;
  assign c_sub59 = (a58 & b_inv58) | (a58 & c58) | (b_inv58 & c58);
  wire s59, sub59, and59, or59;
  wire b_inv59;
  assign b_inv59 = ~b59;
  assign s59  = a59 ^ b59 ^ c59;
  assign sub59 = a59 ^ b_inv59 ^ c59;
  assign and59 = a59 & b59;
  assign or59  = a59 | b59;
  assign c60 = (a59 & b59) | (a59 & c59) | (b59 & c59);
  wire c_sub60;
  assign c_sub60 = (a59 & b_inv59) | (a59 & c59) | (b_inv59 & c59);
  wire s60, sub60, and60, or60;
  wire b_inv60;
  assign b_inv60 = ~b60;
  assign s60  = a60 ^ b60 ^ c60;
  assign sub60 = a60 ^ b_inv60 ^ c60;
  assign and60 = a60 & b60;
  assign or60  = a60 | b60;
  assign c61 = (a60 & b60) | (a60 & c60) | (b60 & c60);
  wire c_sub61;
  assign c_sub61 = (a60 & b_inv60) | (a60 & c60) | (b_inv60 & c60);
  wire s61, sub61, and61, or61;
  wire b_inv61;
  assign b_inv61 = ~b61;
  assign s61  = a61 ^ b61 ^ c61;
  assign sub61 = a61 ^ b_inv61 ^ c61;
  assign and61 = a61 & b61;
  assign or61  = a61 | b61;
  assign c62 = (a61 & b61) | (a61 & c61) | (b61 & c61);
  wire c_sub62;
  assign c_sub62 = (a61 & b_inv61) | (a61 & c61) | (b_inv61 & c61);
  wire s62, sub62, and62, or62;
  wire b_inv62;
  assign b_inv62 = ~b62;
  assign s62  = a62 ^ b62 ^ c62;
  assign sub62 = a62 ^ b_inv62 ^ c62;
  assign and62 = a62 & b62;
  assign or62  = a62 | b62;
  assign c63 = (a62 & b62) | (a62 & c62) | (b62 & c62);
  wire c_sub63;
  assign c_sub63 = (a62 & b_inv62) | (a62 & c62) | (b_inv62 & c62);
  wire s63, sub63, and63, or63;
  wire b_inv63;
  assign b_inv63 = ~b63;
  assign s63  = a63 ^ b63 ^ c63;
  assign sub63 = a63 ^ b_inv63 ^ c63;
  assign and63 = a63 & b63;
  assign or63  = a63 | b63;
  assign c64 = (a63 & b63) | (a63 & c63) | (b63 & c63);
  wire c_sub64;
  assign c_sub64 = (a63 & b_inv63) | (a63 & c63) | (b_inv63 & c63);
  wire s64, sub64, and64, or64;
  wire b_inv64;
  assign b_inv64 = ~b64;
  assign s64  = a64 ^ b64 ^ c64;
  assign sub64 = a64 ^ b_inv64 ^ c64;
  assign and64 = a64 & b64;
  assign or64  = a64 | b64;
  assign c65 = (a64 & b64) | (a64 & c64) | (b64 & c64);
  wire c_sub65;
  assign c_sub65 = (a64 & b_inv64) | (a64 & c64) | (b_inv64 & c64);
  wire s65, sub65, and65, or65;
  wire b_inv65;
  assign b_inv65 = ~b65;
  assign s65  = a65 ^ b65 ^ c65;
  assign sub65 = a65 ^ b_inv65 ^ c65;
  assign and65 = a65 & b65;
  assign or65  = a65 | b65;
  assign c66 = (a65 & b65) | (a65 & c65) | (b65 & c65);
  wire c_sub66;
  assign c_sub66 = (a65 & b_inv65) | (a65 & c65) | (b_inv65 & c65);
  wire s66, sub66, and66, or66;
  wire b_inv66;
  assign b_inv66 = ~b66;
  assign s66  = a66 ^ b66 ^ c66;
  assign sub66 = a66 ^ b_inv66 ^ c66;
  assign and66 = a66 & b66;
  assign or66  = a66 | b66;
  assign c67 = (a66 & b66) | (a66 & c66) | (b66 & c66);
  wire c_sub67;
  assign c_sub67 = (a66 & b_inv66) | (a66 & c66) | (b_inv66 & c66);
  wire s67, sub67, and67, or67;
  wire b_inv67;
  assign b_inv67 = ~b67;
  assign s67  = a67 ^ b67 ^ c67;
  assign sub67 = a67 ^ b_inv67 ^ c67;
  assign and67 = a67 & b67;
  assign or67  = a67 | b67;
  assign c68 = (a67 & b67) | (a67 & c67) | (b67 & c67);
  wire c_sub68;
  assign c_sub68 = (a67 & b_inv67) | (a67 & c67) | (b_inv67 & c67);
  wire s68, sub68, and68, or68;
  wire b_inv68;
  assign b_inv68 = ~b68;
  assign s68  = a68 ^ b68 ^ c68;
  assign sub68 = a68 ^ b_inv68 ^ c68;
  assign and68 = a68 & b68;
  assign or68  = a68 | b68;
  assign c69 = (a68 & b68) | (a68 & c68) | (b68 & c68);
  wire c_sub69;
  assign c_sub69 = (a68 & b_inv68) | (a68 & c68) | (b_inv68 & c68);
  wire s69, sub69, and69, or69;
  wire b_inv69;
  assign b_inv69 = ~b69;
  assign s69  = a69 ^ b69 ^ c69;
  assign sub69 = a69 ^ b_inv69 ^ c69;
  assign and69 = a69 & b69;
  assign or69  = a69 | b69;
  assign c70 = (a69 & b69) | (a69 & c69) | (b69 & c69);
  wire c_sub70;
  assign c_sub70 = (a69 & b_inv69) | (a69 & c69) | (b_inv69 & c69);
  wire s70, sub70, and70, or70;
  wire b_inv70;
  assign b_inv70 = ~b70;
  assign s70  = a70 ^ b70 ^ c70;
  assign sub70 = a70 ^ b_inv70 ^ c70;
  assign and70 = a70 & b70;
  assign or70  = a70 | b70;
  assign c71 = (a70 & b70) | (a70 & c70) | (b70 & c70);
  wire c_sub71;
  assign c_sub71 = (a70 & b_inv70) | (a70 & c70) | (b_inv70 & c70);
  wire s71, sub71, and71, or71;
  wire b_inv71;
  assign b_inv71 = ~b71;
  assign s71  = a71 ^ b71 ^ c71;
  assign sub71 = a71 ^ b_inv71 ^ c71;
  assign and71 = a71 & b71;
  assign or71  = a71 | b71;
  assign c72 = (a71 & b71) | (a71 & c71) | (b71 & c71);
  wire c_sub72;
  assign c_sub72 = (a71 & b_inv71) | (a71 & c71) | (b_inv71 & c71);
  wire s72, sub72, and72, or72;
  wire b_inv72;
  assign b_inv72 = ~b72;
  assign s72  = a72 ^ b72 ^ c72;
  assign sub72 = a72 ^ b_inv72 ^ c72;
  assign and72 = a72 & b72;
  assign or72  = a72 | b72;
  assign c73 = (a72 & b72) | (a72 & c72) | (b72 & c72);
  wire c_sub73;
  assign c_sub73 = (a72 & b_inv72) | (a72 & c72) | (b_inv72 & c72);
  wire s73, sub73, and73, or73;
  wire b_inv73;
  assign b_inv73 = ~b73;
  assign s73  = a73 ^ b73 ^ c73;
  assign sub73 = a73 ^ b_inv73 ^ c73;
  assign and73 = a73 & b73;
  assign or73  = a73 | b73;
  assign c74 = (a73 & b73) | (a73 & c73) | (b73 & c73);
  wire c_sub74;
  assign c_sub74 = (a73 & b_inv73) | (a73 & c73) | (b_inv73 & c73);
  wire s74, sub74, and74, or74;
  wire b_inv74;
  assign b_inv74 = ~b74;
  assign s74  = a74 ^ b74 ^ c74;
  assign sub74 = a74 ^ b_inv74 ^ c74;
  assign and74 = a74 & b74;
  assign or74  = a74 | b74;
  assign c75 = (a74 & b74) | (a74 & c74) | (b74 & c74);
  wire c_sub75;
  assign c_sub75 = (a74 & b_inv74) | (a74 & c74) | (b_inv74 & c74);
  wire s75, sub75, and75, or75;
  wire b_inv75;
  assign b_inv75 = ~b75;
  assign s75  = a75 ^ b75 ^ c75;
  assign sub75 = a75 ^ b_inv75 ^ c75;
  assign and75 = a75 & b75;
  assign or75  = a75 | b75;
  assign c76 = (a75 & b75) | (a75 & c75) | (b75 & c75);
  wire c_sub76;
  assign c_sub76 = (a75 & b_inv75) | (a75 & c75) | (b_inv75 & c75);
  wire s76, sub76, and76, or76;
  wire b_inv76;
  assign b_inv76 = ~b76;
  assign s76  = a76 ^ b76 ^ c76;
  assign sub76 = a76 ^ b_inv76 ^ c76;
  assign and76 = a76 & b76;
  assign or76  = a76 | b76;
  assign c77 = (a76 & b76) | (a76 & c76) | (b76 & c76);
  wire c_sub77;
  assign c_sub77 = (a76 & b_inv76) | (a76 & c76) | (b_inv76 & c76);
  wire s77, sub77, and77, or77;
  wire b_inv77;
  assign b_inv77 = ~b77;
  assign s77  = a77 ^ b77 ^ c77;
  assign sub77 = a77 ^ b_inv77 ^ c77;
  assign and77 = a77 & b77;
  assign or77  = a77 | b77;
  assign c78 = (a77 & b77) | (a77 & c77) | (b77 & c77);
  wire c_sub78;
  assign c_sub78 = (a77 & b_inv77) | (a77 & c77) | (b_inv77 & c77);
  wire s78, sub78, and78, or78;
  wire b_inv78;
  assign b_inv78 = ~b78;
  assign s78  = a78 ^ b78 ^ c78;
  assign sub78 = a78 ^ b_inv78 ^ c78;
  assign and78 = a78 & b78;
  assign or78  = a78 | b78;
  assign c79 = (a78 & b78) | (a78 & c78) | (b78 & c78);
  wire c_sub79;
  assign c_sub79 = (a78 & b_inv78) | (a78 & c78) | (b_inv78 & c78);
  wire s79, sub79, and79, or79;
  wire b_inv79;
  assign b_inv79 = ~b79;
  assign s79  = a79 ^ b79 ^ c79;
  assign sub79 = a79 ^ b_inv79 ^ c79;
  assign and79 = a79 & b79;
  assign or79  = a79 | b79;
  assign c80 = (a79 & b79) | (a79 & c79) | (b79 & c79);
  wire c_sub80;
  assign c_sub80 = (a79 & b_inv79) | (a79 & c79) | (b_inv79 & c79);
  wire s80, sub80, and80, or80;
  wire b_inv80;
  assign b_inv80 = ~b80;
  assign s80  = a80 ^ b80 ^ c80;
  assign sub80 = a80 ^ b_inv80 ^ c80;
  assign and80 = a80 & b80;
  assign or80  = a80 | b80;
  assign c81 = (a80 & b80) | (a80 & c80) | (b80 & c80);
  wire c_sub81;
  assign c_sub81 = (a80 & b_inv80) | (a80 & c80) | (b_inv80 & c80);
  wire s81, sub81, and81, or81;
  wire b_inv81;
  assign b_inv81 = ~b81;
  assign s81  = a81 ^ b81 ^ c81;
  assign sub81 = a81 ^ b_inv81 ^ c81;
  assign and81 = a81 & b81;
  assign or81  = a81 | b81;
  assign c82 = (a81 & b81) | (a81 & c81) | (b81 & c81);
  wire c_sub82;
  assign c_sub82 = (a81 & b_inv81) | (a81 & c81) | (b_inv81 & c81);
  wire s82, sub82, and82, or82;
  wire b_inv82;
  assign b_inv82 = ~b82;
  assign s82  = a82 ^ b82 ^ c82;
  assign sub82 = a82 ^ b_inv82 ^ c82;
  assign and82 = a82 & b82;
  assign or82  = a82 | b82;
  assign c83 = (a82 & b82) | (a82 & c82) | (b82 & c82);
  wire c_sub83;
  assign c_sub83 = (a82 & b_inv82) | (a82 & c82) | (b_inv82 & c82);
  wire s83, sub83, and83, or83;
  wire b_inv83;
  assign b_inv83 = ~b83;
  assign s83  = a83 ^ b83 ^ c83;
  assign sub83 = a83 ^ b_inv83 ^ c83;
  assign and83 = a83 & b83;
  assign or83  = a83 | b83;
  assign c84 = (a83 & b83) | (a83 & c83) | (b83 & c83);
  wire c_sub84;
  assign c_sub84 = (a83 & b_inv83) | (a83 & c83) | (b_inv83 & c83);
  wire s84, sub84, and84, or84;
  wire b_inv84;
  assign b_inv84 = ~b84;
  assign s84  = a84 ^ b84 ^ c84;
  assign sub84 = a84 ^ b_inv84 ^ c84;
  assign and84 = a84 & b84;
  assign or84  = a84 | b84;
  assign c85 = (a84 & b84) | (a84 & c84) | (b84 & c84);
  wire c_sub85;
  assign c_sub85 = (a84 & b_inv84) | (a84 & c84) | (b_inv84 & c84);
  wire s85, sub85, and85, or85;
  wire b_inv85;
  assign b_inv85 = ~b85;
  assign s85  = a85 ^ b85 ^ c85;
  assign sub85 = a85 ^ b_inv85 ^ c85;
  assign and85 = a85 & b85;
  assign or85  = a85 | b85;
  assign c86 = (a85 & b85) | (a85 & c85) | (b85 & c85);
  wire c_sub86;
  assign c_sub86 = (a85 & b_inv85) | (a85 & c85) | (b_inv85 & c85);
  wire s86, sub86, and86, or86;
  wire b_inv86;
  assign b_inv86 = ~b86;
  assign s86  = a86 ^ b86 ^ c86;
  assign sub86 = a86 ^ b_inv86 ^ c86;
  assign and86 = a86 & b86;
  assign or86  = a86 | b86;
  assign c87 = (a86 & b86) | (a86 & c86) | (b86 & c86);
  wire c_sub87;
  assign c_sub87 = (a86 & b_inv86) | (a86 & c86) | (b_inv86 & c86);
  wire s87, sub87, and87, or87;
  wire b_inv87;
  assign b_inv87 = ~b87;
  assign s87  = a87 ^ b87 ^ c87;
  assign sub87 = a87 ^ b_inv87 ^ c87;
  assign and87 = a87 & b87;
  assign or87  = a87 | b87;
  assign c88 = (a87 & b87) | (a87 & c87) | (b87 & c87);
  wire c_sub88;
  assign c_sub88 = (a87 & b_inv87) | (a87 & c87) | (b_inv87 & c87);
  wire s88, sub88, and88, or88;
  wire b_inv88;
  assign b_inv88 = ~b88;
  assign s88  = a88 ^ b88 ^ c88;
  assign sub88 = a88 ^ b_inv88 ^ c88;
  assign and88 = a88 & b88;
  assign or88  = a88 | b88;
  assign c89 = (a88 & b88) | (a88 & c88) | (b88 & c88);
  wire c_sub89;
  assign c_sub89 = (a88 & b_inv88) | (a88 & c88) | (b_inv88 & c88);
  wire s89, sub89, and89, or89;
  wire b_inv89;
  assign b_inv89 = ~b89;
  assign s89  = a89 ^ b89 ^ c89;
  assign sub89 = a89 ^ b_inv89 ^ c89;
  assign and89 = a89 & b89;
  assign or89  = a89 | b89;
  assign c90 = (a89 & b89) | (a89 & c89) | (b89 & c89);
  wire c_sub90;
  assign c_sub90 = (a89 & b_inv89) | (a89 & c89) | (b_inv89 & c89);
  wire s90, sub90, and90, or90;
  wire b_inv90;
  assign b_inv90 = ~b90;
  assign s90  = a90 ^ b90 ^ c90;
  assign sub90 = a90 ^ b_inv90 ^ c90;
  assign and90 = a90 & b90;
  assign or90  = a90 | b90;
  assign c91 = (a90 & b90) | (a90 & c90) | (b90 & c90);
  wire c_sub91;
  assign c_sub91 = (a90 & b_inv90) | (a90 & c90) | (b_inv90 & c90);
  wire s91, sub91, and91, or91;
  wire b_inv91;
  assign b_inv91 = ~b91;
  assign s91  = a91 ^ b91 ^ c91;
  assign sub91 = a91 ^ b_inv91 ^ c91;
  assign and91 = a91 & b91;
  assign or91  = a91 | b91;
  assign c92 = (a91 & b91) | (a91 & c91) | (b91 & c91);
  wire c_sub92;
  assign c_sub92 = (a91 & b_inv91) | (a91 & c91) | (b_inv91 & c91);
  wire s92, sub92, and92, or92;
  wire b_inv92;
  assign b_inv92 = ~b92;
  assign s92  = a92 ^ b92 ^ c92;
  assign sub92 = a92 ^ b_inv92 ^ c92;
  assign and92 = a92 & b92;
  assign or92  = a92 | b92;
  assign c93 = (a92 & b92) | (a92 & c92) | (b92 & c92);
  wire c_sub93;
  assign c_sub93 = (a92 & b_inv92) | (a92 & c92) | (b_inv92 & c92);
  wire s93, sub93, and93, or93;
  wire b_inv93;
  assign b_inv93 = ~b93;
  assign s93  = a93 ^ b93 ^ c93;
  assign sub93 = a93 ^ b_inv93 ^ c93;
  assign and93 = a93 & b93;
  assign or93  = a93 | b93;
  assign c94 = (a93 & b93) | (a93 & c93) | (b93 & c93);
  wire c_sub94;
  assign c_sub94 = (a93 & b_inv93) | (a93 & c93) | (b_inv93 & c93);
  wire s94, sub94, and94, or94;
  wire b_inv94;
  assign b_inv94 = ~b94;
  assign s94  = a94 ^ b94 ^ c94;
  assign sub94 = a94 ^ b_inv94 ^ c94;
  assign and94 = a94 & b94;
  assign or94  = a94 | b94;
  assign c95 = (a94 & b94) | (a94 & c94) | (b94 & c94);
  wire c_sub95;
  assign c_sub95 = (a94 & b_inv94) | (a94 & c94) | (b_inv94 & c94);
  wire s95, sub95, and95, or95;
  wire b_inv95;
  assign b_inv95 = ~b95;
  assign s95  = a95 ^ b95 ^ c95;
  assign sub95 = a95 ^ b_inv95 ^ c95;
  assign and95 = a95 & b95;
  assign or95  = a95 | b95;
  assign c96 = (a95 & b95) | (a95 & c95) | (b95 & c95);
  wire c_sub96;
  assign c_sub96 = (a95 & b_inv95) | (a95 & c95) | (b_inv95 & c95);
  wire s96, sub96, and96, or96;
  wire b_inv96;
  assign b_inv96 = ~b96;
  assign s96  = a96 ^ b96 ^ c96;
  assign sub96 = a96 ^ b_inv96 ^ c96;
  assign and96 = a96 & b96;
  assign or96  = a96 | b96;
  assign c97 = (a96 & b96) | (a96 & c96) | (b96 & c96);
  wire c_sub97;
  assign c_sub97 = (a96 & b_inv96) | (a96 & c96) | (b_inv96 & c96);
  wire s97, sub97, and97, or97;
  wire b_inv97;
  assign b_inv97 = ~b97;
  assign s97  = a97 ^ b97 ^ c97;
  assign sub97 = a97 ^ b_inv97 ^ c97;
  assign and97 = a97 & b97;
  assign or97  = a97 | b97;
  assign c98 = (a97 & b97) | (a97 & c97) | (b97 & c97);
  wire c_sub98;
  assign c_sub98 = (a97 & b_inv97) | (a97 & c97) | (b_inv97 & c97);
  wire s98, sub98, and98, or98;
  wire b_inv98;
  assign b_inv98 = ~b98;
  assign s98  = a98 ^ b98 ^ c98;
  assign sub98 = a98 ^ b_inv98 ^ c98;
  assign and98 = a98 & b98;
  assign or98  = a98 | b98;
  assign c99 = (a98 & b98) | (a98 & c98) | (b98 & c98);
  wire c_sub99;
  assign c_sub99 = (a98 & b_inv98) | (a98 & c98) | (b_inv98 & c98);
  wire s99, sub99, and99, or99;
  wire b_inv99;
  assign b_inv99 = ~b99;
  assign s99  = a99 ^ b99 ^ c99;
  assign sub99 = a99 ^ b_inv99 ^ c99;
  assign and99 = a99 & b99;
  assign or99  = a99 | b99;
  assign c100 = (a99 & b99) | (a99 & c99) | (b99 & c99);
  wire c_sub100;
  assign c_sub100 = (a99 & b_inv99) | (a99 & c99) | (b_inv99 & c99);
  wire s100, sub100, and100, or100;
  wire b_inv100;
  assign b_inv100 = ~b100;
  assign s100  = a100 ^ b100 ^ c100;
  assign sub100 = a100 ^ b_inv100 ^ c100;
  assign and100 = a100 & b100;
  assign or100  = a100 | b100;
  assign c101 = (a100 & b100) | (a100 & c100) | (b100 & c100);
  wire c_sub101;
  assign c_sub101 = (a100 & b_inv100) | (a100 & c100) | (b_inv100 & c100);
  wire s101, sub101, and101, or101;
  wire b_inv101;
  assign b_inv101 = ~b101;
  assign s101  = a101 ^ b101 ^ c101;
  assign sub101 = a101 ^ b_inv101 ^ c101;
  assign and101 = a101 & b101;
  assign or101  = a101 | b101;
  assign c102 = (a101 & b101) | (a101 & c101) | (b101 & c101);
  wire c_sub102;
  assign c_sub102 = (a101 & b_inv101) | (a101 & c101) | (b_inv101 & c101);
  wire s102, sub102, and102, or102;
  wire b_inv102;
  assign b_inv102 = ~b102;
  assign s102  = a102 ^ b102 ^ c102;
  assign sub102 = a102 ^ b_inv102 ^ c102;
  assign and102 = a102 & b102;
  assign or102  = a102 | b102;
  assign c103 = (a102 & b102) | (a102 & c102) | (b102 & c102);
  wire c_sub103;
  assign c_sub103 = (a102 & b_inv102) | (a102 & c102) | (b_inv102 & c102);
  wire s103, sub103, and103, or103;
  wire b_inv103;
  assign b_inv103 = ~b103;
  assign s103  = a103 ^ b103 ^ c103;
  assign sub103 = a103 ^ b_inv103 ^ c103;
  assign and103 = a103 & b103;
  assign or103  = a103 | b103;
  assign c104 = (a103 & b103) | (a103 & c103) | (b103 & c103);
  wire c_sub104;
  assign c_sub104 = (a103 & b_inv103) | (a103 & c103) | (b_inv103 & c103);
  wire s104, sub104, and104, or104;
  wire b_inv104;
  assign b_inv104 = ~b104;
  assign s104  = a104 ^ b104 ^ c104;
  assign sub104 = a104 ^ b_inv104 ^ c104;
  assign and104 = a104 & b104;
  assign or104  = a104 | b104;
  assign c105 = (a104 & b104) | (a104 & c104) | (b104 & c104);
  wire c_sub105;
  assign c_sub105 = (a104 & b_inv104) | (a104 & c104) | (b_inv104 & c104);
  wire s105, sub105, and105, or105;
  wire b_inv105;
  assign b_inv105 = ~b105;
  assign s105  = a105 ^ b105 ^ c105;
  assign sub105 = a105 ^ b_inv105 ^ c105;
  assign and105 = a105 & b105;
  assign or105  = a105 | b105;
  assign c106 = (a105 & b105) | (a105 & c105) | (b105 & c105);
  wire c_sub106;
  assign c_sub106 = (a105 & b_inv105) | (a105 & c105) | (b_inv105 & c105);
  wire s106, sub106, and106, or106;
  wire b_inv106;
  assign b_inv106 = ~b106;
  assign s106  = a106 ^ b106 ^ c106;
  assign sub106 = a106 ^ b_inv106 ^ c106;
  assign and106 = a106 & b106;
  assign or106  = a106 | b106;
  assign c107 = (a106 & b106) | (a106 & c106) | (b106 & c106);
  wire c_sub107;
  assign c_sub107 = (a106 & b_inv106) | (a106 & c106) | (b_inv106 & c106);
  wire s107, sub107, and107, or107;
  wire b_inv107;
  assign b_inv107 = ~b107;
  assign s107  = a107 ^ b107 ^ c107;
  assign sub107 = a107 ^ b_inv107 ^ c107;
  assign and107 = a107 & b107;
  assign or107  = a107 | b107;
  assign c108 = (a107 & b107) | (a107 & c107) | (b107 & c107);
  wire c_sub108;
  assign c_sub108 = (a107 & b_inv107) | (a107 & c107) | (b_inv107 & c107);
  wire s108, sub108, and108, or108;
  wire b_inv108;
  assign b_inv108 = ~b108;
  assign s108  = a108 ^ b108 ^ c108;
  assign sub108 = a108 ^ b_inv108 ^ c108;
  assign and108 = a108 & b108;
  assign or108  = a108 | b108;
  assign c109 = (a108 & b108) | (a108 & c108) | (b108 & c108);
  wire c_sub109;
  assign c_sub109 = (a108 & b_inv108) | (a108 & c108) | (b_inv108 & c108);
  wire s109, sub109, and109, or109;
  wire b_inv109;
  assign b_inv109 = ~b109;
  assign s109  = a109 ^ b109 ^ c109;
  assign sub109 = a109 ^ b_inv109 ^ c109;
  assign and109 = a109 & b109;
  assign or109  = a109 | b109;
  assign c110 = (a109 & b109) | (a109 & c109) | (b109 & c109);
  wire c_sub110;
  assign c_sub110 = (a109 & b_inv109) | (a109 & c109) | (b_inv109 & c109);
  wire s110, sub110, and110, or110;
  wire b_inv110;
  assign b_inv110 = ~b110;
  assign s110  = a110 ^ b110 ^ c110;
  assign sub110 = a110 ^ b_inv110 ^ c110;
  assign and110 = a110 & b110;
  assign or110  = a110 | b110;
  assign c111 = (a110 & b110) | (a110 & c110) | (b110 & c110);
  wire c_sub111;
  assign c_sub111 = (a110 & b_inv110) | (a110 & c110) | (b_inv110 & c110);
  wire s111, sub111, and111, or111;
  wire b_inv111;
  assign b_inv111 = ~b111;
  assign s111  = a111 ^ b111 ^ c111;
  assign sub111 = a111 ^ b_inv111 ^ c111;
  assign and111 = a111 & b111;
  assign or111  = a111 | b111;
  assign c112 = (a111 & b111) | (a111 & c111) | (b111 & c111);
  wire c_sub112;
  assign c_sub112 = (a111 & b_inv111) | (a111 & c111) | (b_inv111 & c111);
  wire s112, sub112, and112, or112;
  wire b_inv112;
  assign b_inv112 = ~b112;
  assign s112  = a112 ^ b112 ^ c112;
  assign sub112 = a112 ^ b_inv112 ^ c112;
  assign and112 = a112 & b112;
  assign or112  = a112 | b112;
  assign c113 = (a112 & b112) | (a112 & c112) | (b112 & c112);
  wire c_sub113;
  assign c_sub113 = (a112 & b_inv112) | (a112 & c112) | (b_inv112 & c112);
  wire s113, sub113, and113, or113;
  wire b_inv113;
  assign b_inv113 = ~b113;
  assign s113  = a113 ^ b113 ^ c113;
  assign sub113 = a113 ^ b_inv113 ^ c113;
  assign and113 = a113 & b113;
  assign or113  = a113 | b113;
  assign c114 = (a113 & b113) | (a113 & c113) | (b113 & c113);
  wire c_sub114;
  assign c_sub114 = (a113 & b_inv113) | (a113 & c113) | (b_inv113 & c113);
  wire s114, sub114, and114, or114;
  wire b_inv114;
  assign b_inv114 = ~b114;
  assign s114  = a114 ^ b114 ^ c114;
  assign sub114 = a114 ^ b_inv114 ^ c114;
  assign and114 = a114 & b114;
  assign or114  = a114 | b114;
  assign c115 = (a114 & b114) | (a114 & c114) | (b114 & c114);
  wire c_sub115;
  assign c_sub115 = (a114 & b_inv114) | (a114 & c114) | (b_inv114 & c114);
  wire s115, sub115, and115, or115;
  wire b_inv115;
  assign b_inv115 = ~b115;
  assign s115  = a115 ^ b115 ^ c115;
  assign sub115 = a115 ^ b_inv115 ^ c115;
  assign and115 = a115 & b115;
  assign or115  = a115 | b115;
  assign c116 = (a115 & b115) | (a115 & c115) | (b115 & c115);
  wire c_sub116;
  assign c_sub116 = (a115 & b_inv115) | (a115 & c115) | (b_inv115 & c115);
  wire s116, sub116, and116, or116;
  wire b_inv116;
  assign b_inv116 = ~b116;
  assign s116  = a116 ^ b116 ^ c116;
  assign sub116 = a116 ^ b_inv116 ^ c116;
  assign and116 = a116 & b116;
  assign or116  = a116 | b116;
  assign c117 = (a116 & b116) | (a116 & c116) | (b116 & c116);
  wire c_sub117;
  assign c_sub117 = (a116 & b_inv116) | (a116 & c116) | (b_inv116 & c116);
  wire s117, sub117, and117, or117;
  wire b_inv117;
  assign b_inv117 = ~b117;
  assign s117  = a117 ^ b117 ^ c117;
  assign sub117 = a117 ^ b_inv117 ^ c117;
  assign and117 = a117 & b117;
  assign or117  = a117 | b117;
  assign c118 = (a117 & b117) | (a117 & c117) | (b117 & c117);
  wire c_sub118;
  assign c_sub118 = (a117 & b_inv117) | (a117 & c117) | (b_inv117 & c117);
  wire s118, sub118, and118, or118;
  wire b_inv118;
  assign b_inv118 = ~b118;
  assign s118  = a118 ^ b118 ^ c118;
  assign sub118 = a118 ^ b_inv118 ^ c118;
  assign and118 = a118 & b118;
  assign or118  = a118 | b118;
  assign c119 = (a118 & b118) | (a118 & c118) | (b118 & c118);
  wire c_sub119;
  assign c_sub119 = (a118 & b_inv118) | (a118 & c118) | (b_inv118 & c118);
  wire s119, sub119, and119, or119;
  wire b_inv119;
  assign b_inv119 = ~b119;
  assign s119  = a119 ^ b119 ^ c119;
  assign sub119 = a119 ^ b_inv119 ^ c119;
  assign and119 = a119 & b119;
  assign or119  = a119 | b119;
  assign c120 = (a119 & b119) | (a119 & c119) | (b119 & c119);
  wire c_sub120;
  assign c_sub120 = (a119 & b_inv119) | (a119 & c119) | (b_inv119 & c119);
  wire s120, sub120, and120, or120;
  wire b_inv120;
  assign b_inv120 = ~b120;
  assign s120  = a120 ^ b120 ^ c120;
  assign sub120 = a120 ^ b_inv120 ^ c120;
  assign and120 = a120 & b120;
  assign or120  = a120 | b120;
  assign c121 = (a120 & b120) | (a120 & c120) | (b120 & c120);
  wire c_sub121;
  assign c_sub121 = (a120 & b_inv120) | (a120 & c120) | (b_inv120 & c120);
  wire s121, sub121, and121, or121;
  wire b_inv121;
  assign b_inv121 = ~b121;
  assign s121  = a121 ^ b121 ^ c121;
  assign sub121 = a121 ^ b_inv121 ^ c121;
  assign and121 = a121 & b121;
  assign or121  = a121 | b121;
  assign c122 = (a121 & b121) | (a121 & c121) | (b121 & c121);
  wire c_sub122;
  assign c_sub122 = (a121 & b_inv121) | (a121 & c121) | (b_inv121 & c121);
  wire s122, sub122, and122, or122;
  wire b_inv122;
  assign b_inv122 = ~b122;
  assign s122  = a122 ^ b122 ^ c122;
  assign sub122 = a122 ^ b_inv122 ^ c122;
  assign and122 = a122 & b122;
  assign or122  = a122 | b122;
  assign c123 = (a122 & b122) | (a122 & c122) | (b122 & c122);
  wire c_sub123;
  assign c_sub123 = (a122 & b_inv122) | (a122 & c122) | (b_inv122 & c122);
  wire s123, sub123, and123, or123;
  wire b_inv123;
  assign b_inv123 = ~b123;
  assign s123  = a123 ^ b123 ^ c123;
  assign sub123 = a123 ^ b_inv123 ^ c123;
  assign and123 = a123 & b123;
  assign or123  = a123 | b123;
  assign c124 = (a123 & b123) | (a123 & c123) | (b123 & c123);
  wire c_sub124;
  assign c_sub124 = (a123 & b_inv123) | (a123 & c123) | (b_inv123 & c123);
  wire s124, sub124, and124, or124;
  wire b_inv124;
  assign b_inv124 = ~b124;
  assign s124  = a124 ^ b124 ^ c124;
  assign sub124 = a124 ^ b_inv124 ^ c124;
  assign and124 = a124 & b124;
  assign or124  = a124 | b124;
  assign c125 = (a124 & b124) | (a124 & c124) | (b124 & c124);
  wire c_sub125;
  assign c_sub125 = (a124 & b_inv124) | (a124 & c124) | (b_inv124 & c124);
  wire s125, sub125, and125, or125;
  wire b_inv125;
  assign b_inv125 = ~b125;
  assign s125  = a125 ^ b125 ^ c125;
  assign sub125 = a125 ^ b_inv125 ^ c125;
  assign and125 = a125 & b125;
  assign or125  = a125 | b125;
  assign c126 = (a125 & b125) | (a125 & c125) | (b125 & c125);
  wire c_sub126;
  assign c_sub126 = (a125 & b_inv125) | (a125 & c125) | (b_inv125 & c125);
  wire s126, sub126, and126, or126;
  wire b_inv126;
  assign b_inv126 = ~b126;
  assign s126  = a126 ^ b126 ^ c126;
  assign sub126 = a126 ^ b_inv126 ^ c126;
  assign and126 = a126 & b126;
  assign or126  = a126 | b126;
  assign c127 = (a126 & b126) | (a126 & c126) | (b126 & c126);
  wire c_sub127;
  assign c_sub127 = (a126 & b_inv126) | (a126 & c126) | (b_inv126 & c126);
  wire s127, sub127, and127, or127;
  wire b_inv127;
  assign b_inv127 = ~b127;
  assign s127  = a127 ^ b127 ^ c127;
  assign sub127 = a127 ^ b_inv127 ^ c127;
  assign and127 = a127 & b127;
  assign or127  = a127 | b127;
  assign c128 = (a127 & b127) | (a127 & c127) | (b127 & c127);
  wire c_sub128;
  assign c_sub128 = (a127 & b_inv127) | (a127 & c127) | (b_inv127 & c127);
  wire s128, sub128, and128, or128;
  wire b_inv128;
  assign b_inv128 = ~b128;
  assign s128  = a128 ^ b128 ^ c128;
  assign sub128 = a128 ^ b_inv128 ^ c128;
  assign and128 = a128 & b128;
  assign or128  = a128 | b128;
  assign c129 = (a128 & b128) | (a128 & c128) | (b128 & c128);
  wire c_sub129;
  assign c_sub129 = (a128 & b_inv128) | (a128 & c128) | (b_inv128 & c128);
  wire s129, sub129, and129, or129;
  wire b_inv129;
  assign b_inv129 = ~b129;
  assign s129  = a129 ^ b129 ^ c129;
  assign sub129 = a129 ^ b_inv129 ^ c129;
  assign and129 = a129 & b129;
  assign or129  = a129 | b129;
  assign c130 = (a129 & b129) | (a129 & c129) | (b129 & c129);
  wire c_sub130;
  assign c_sub130 = (a129 & b_inv129) | (a129 & c129) | (b_inv129 & c129);
  wire s130, sub130, and130, or130;
  wire b_inv130;
  assign b_inv130 = ~b130;
  assign s130  = a130 ^ b130 ^ c130;
  assign sub130 = a130 ^ b_inv130 ^ c130;
  assign and130 = a130 & b130;
  assign or130  = a130 | b130;
  assign c131 = (a130 & b130) | (a130 & c130) | (b130 & c130);
  wire c_sub131;
  assign c_sub131 = (a130 & b_inv130) | (a130 & c130) | (b_inv130 & c130);
  wire s131, sub131, and131, or131;
  wire b_inv131;
  assign b_inv131 = ~b131;
  assign s131  = a131 ^ b131 ^ c131;
  assign sub131 = a131 ^ b_inv131 ^ c131;
  assign and131 = a131 & b131;
  assign or131  = a131 | b131;
  assign c132 = (a131 & b131) | (a131 & c131) | (b131 & c131);
  wire c_sub132;
  assign c_sub132 = (a131 & b_inv131) | (a131 & c131) | (b_inv131 & c131);
  wire s132, sub132, and132, or132;
  wire b_inv132;
  assign b_inv132 = ~b132;
  assign s132  = a132 ^ b132 ^ c132;
  assign sub132 = a132 ^ b_inv132 ^ c132;
  assign and132 = a132 & b132;
  assign or132  = a132 | b132;
  assign c133 = (a132 & b132) | (a132 & c132) | (b132 & c132);
  wire c_sub133;
  assign c_sub133 = (a132 & b_inv132) | (a132 & c132) | (b_inv132 & c132);
  wire s133, sub133, and133, or133;
  wire b_inv133;
  assign b_inv133 = ~b133;
  assign s133  = a133 ^ b133 ^ c133;
  assign sub133 = a133 ^ b_inv133 ^ c133;
  assign and133 = a133 & b133;
  assign or133  = a133 | b133;
  assign c134 = (a133 & b133) | (a133 & c133) | (b133 & c133);
  wire c_sub134;
  assign c_sub134 = (a133 & b_inv133) | (a133 & c133) | (b_inv133 & c133);
  wire s134, sub134, and134, or134;
  wire b_inv134;
  assign b_inv134 = ~b134;
  assign s134  = a134 ^ b134 ^ c134;
  assign sub134 = a134 ^ b_inv134 ^ c134;
  assign and134 = a134 & b134;
  assign or134  = a134 | b134;
  assign c135 = (a134 & b134) | (a134 & c134) | (b134 & c134);
  wire c_sub135;
  assign c_sub135 = (a134 & b_inv134) | (a134 & c134) | (b_inv134 & c134);
  wire s135, sub135, and135, or135;
  wire b_inv135;
  assign b_inv135 = ~b135;
  assign s135  = a135 ^ b135 ^ c135;
  assign sub135 = a135 ^ b_inv135 ^ c135;
  assign and135 = a135 & b135;
  assign or135  = a135 | b135;
  assign c136 = (a135 & b135) | (a135 & c135) | (b135 & c135);
  wire c_sub136;
  assign c_sub136 = (a135 & b_inv135) | (a135 & c135) | (b_inv135 & c135);
  wire s136, sub136, and136, or136;
  wire b_inv136;
  assign b_inv136 = ~b136;
  assign s136  = a136 ^ b136 ^ c136;
  assign sub136 = a136 ^ b_inv136 ^ c136;
  assign and136 = a136 & b136;
  assign or136  = a136 | b136;
  assign c137 = (a136 & b136) | (a136 & c136) | (b136 & c136);
  wire c_sub137;
  assign c_sub137 = (a136 & b_inv136) | (a136 & c136) | (b_inv136 & c136);
  wire s137, sub137, and137, or137;
  wire b_inv137;
  assign b_inv137 = ~b137;
  assign s137  = a137 ^ b137 ^ c137;
  assign sub137 = a137 ^ b_inv137 ^ c137;
  assign and137 = a137 & b137;
  assign or137  = a137 | b137;
  assign c138 = (a137 & b137) | (a137 & c137) | (b137 & c137);
  wire c_sub138;
  assign c_sub138 = (a137 & b_inv137) | (a137 & c137) | (b_inv137 & c137);
  wire s138, sub138, and138, or138;
  wire b_inv138;
  assign b_inv138 = ~b138;
  assign s138  = a138 ^ b138 ^ c138;
  assign sub138 = a138 ^ b_inv138 ^ c138;
  assign and138 = a138 & b138;
  assign or138  = a138 | b138;
  assign c139 = (a138 & b138) | (a138 & c138) | (b138 & c138);
  wire c_sub139;
  assign c_sub139 = (a138 & b_inv138) | (a138 & c138) | (b_inv138 & c138);
  wire s139, sub139, and139, or139;
  wire b_inv139;
  assign b_inv139 = ~b139;
  assign s139  = a139 ^ b139 ^ c139;
  assign sub139 = a139 ^ b_inv139 ^ c139;
  assign and139 = a139 & b139;
  assign or139  = a139 | b139;
  assign c140 = (a139 & b139) | (a139 & c139) | (b139 & c139);
  wire c_sub140;
  assign c_sub140 = (a139 & b_inv139) | (a139 & c139) | (b_inv139 & c139);
  wire s140, sub140, and140, or140;
  wire b_inv140;
  assign b_inv140 = ~b140;
  assign s140  = a140 ^ b140 ^ c140;
  assign sub140 = a140 ^ b_inv140 ^ c140;
  assign and140 = a140 & b140;
  assign or140  = a140 | b140;
  assign c141 = (a140 & b140) | (a140 & c140) | (b140 & c140);
  wire c_sub141;
  assign c_sub141 = (a140 & b_inv140) | (a140 & c140) | (b_inv140 & c140);
  wire s141, sub141, and141, or141;
  wire b_inv141;
  assign b_inv141 = ~b141;
  assign s141  = a141 ^ b141 ^ c141;
  assign sub141 = a141 ^ b_inv141 ^ c141;
  assign and141 = a141 & b141;
  assign or141  = a141 | b141;
  assign c142 = (a141 & b141) | (a141 & c141) | (b141 & c141);
  wire c_sub142;
  assign c_sub142 = (a141 & b_inv141) | (a141 & c141) | (b_inv141 & c141);
  wire s142, sub142, and142, or142;
  wire b_inv142;
  assign b_inv142 = ~b142;
  assign s142  = a142 ^ b142 ^ c142;
  assign sub142 = a142 ^ b_inv142 ^ c142;
  assign and142 = a142 & b142;
  assign or142  = a142 | b142;
  assign c143 = (a142 & b142) | (a142 & c142) | (b142 & c142);
  wire c_sub143;
  assign c_sub143 = (a142 & b_inv142) | (a142 & c142) | (b_inv142 & c142);
  wire s143, sub143, and143, or143;
  wire b_inv143;
  assign b_inv143 = ~b143;
  assign s143  = a143 ^ b143 ^ c143;
  assign sub143 = a143 ^ b_inv143 ^ c143;
  assign and143 = a143 & b143;
  assign or143  = a143 | b143;
  assign c144 = (a143 & b143) | (a143 & c143) | (b143 & c143);
  wire c_sub144;
  assign c_sub144 = (a143 & b_inv143) | (a143 & c143) | (b_inv143 & c143);
  wire s144, sub144, and144, or144;
  wire b_inv144;
  assign b_inv144 = ~b144;
  assign s144  = a144 ^ b144 ^ c144;
  assign sub144 = a144 ^ b_inv144 ^ c144;
  assign and144 = a144 & b144;
  assign or144  = a144 | b144;
  assign c145 = (a144 & b144) | (a144 & c144) | (b144 & c144);
  wire c_sub145;
  assign c_sub145 = (a144 & b_inv144) | (a144 & c144) | (b_inv144 & c144);
  wire s145, sub145, and145, or145;
  wire b_inv145;
  assign b_inv145 = ~b145;
  assign s145  = a145 ^ b145 ^ c145;
  assign sub145 = a145 ^ b_inv145 ^ c145;
  assign and145 = a145 & b145;
  assign or145  = a145 | b145;
  assign c146 = (a145 & b145) | (a145 & c145) | (b145 & c145);
  wire c_sub146;
  assign c_sub146 = (a145 & b_inv145) | (a145 & c145) | (b_inv145 & c145);
  wire s146, sub146, and146, or146;
  wire b_inv146;
  assign b_inv146 = ~b146;
  assign s146  = a146 ^ b146 ^ c146;
  assign sub146 = a146 ^ b_inv146 ^ c146;
  assign and146 = a146 & b146;
  assign or146  = a146 | b146;
  assign c147 = (a146 & b146) | (a146 & c146) | (b146 & c146);
  wire c_sub147;
  assign c_sub147 = (a146 & b_inv146) | (a146 & c146) | (b_inv146 & c146);
  wire s147, sub147, and147, or147;
  wire b_inv147;
  assign b_inv147 = ~b147;
  assign s147  = a147 ^ b147 ^ c147;
  assign sub147 = a147 ^ b_inv147 ^ c147;
  assign and147 = a147 & b147;
  assign or147  = a147 | b147;
  assign c148 = (a147 & b147) | (a147 & c147) | (b147 & c147);
  wire c_sub148;
  assign c_sub148 = (a147 & b_inv147) | (a147 & c147) | (b_inv147 & c147);
  wire s148, sub148, and148, or148;
  wire b_inv148;
  assign b_inv148 = ~b148;
  assign s148  = a148 ^ b148 ^ c148;
  assign sub148 = a148 ^ b_inv148 ^ c148;
  assign and148 = a148 & b148;
  assign or148  = a148 | b148;
  assign c149 = (a148 & b148) | (a148 & c148) | (b148 & c148);
  wire c_sub149;
  assign c_sub149 = (a148 & b_inv148) | (a148 & c148) | (b_inv148 & c148);
  wire s149, sub149, and149, or149;
  wire b_inv149;
  assign b_inv149 = ~b149;
  assign s149  = a149 ^ b149 ^ c149;
  assign sub149 = a149 ^ b_inv149 ^ c149;
  assign and149 = a149 & b149;
  assign or149  = a149 | b149;
  assign c150 = (a149 & b149) | (a149 & c149) | (b149 & c149);
  wire c_sub150;
  assign c_sub150 = (a149 & b_inv149) | (a149 & c149) | (b_inv149 & c149);
  wire s150, sub150, and150, or150;
  wire b_inv150;
  assign b_inv150 = ~b150;
  assign s150  = a150 ^ b150 ^ c150;
  assign sub150 = a150 ^ b_inv150 ^ c150;
  assign and150 = a150 & b150;
  assign or150  = a150 | b150;
  assign c151 = (a150 & b150) | (a150 & c150) | (b150 & c150);
  wire c_sub151;
  assign c_sub151 = (a150 & b_inv150) | (a150 & c150) | (b_inv150 & c150);
  wire s151, sub151, and151, or151;
  wire b_inv151;
  assign b_inv151 = ~b151;
  assign s151  = a151 ^ b151 ^ c151;
  assign sub151 = a151 ^ b_inv151 ^ c151;
  assign and151 = a151 & b151;
  assign or151  = a151 | b151;
  assign c152 = (a151 & b151) | (a151 & c151) | (b151 & c151);
  wire c_sub152;
  assign c_sub152 = (a151 & b_inv151) | (a151 & c151) | (b_inv151 & c151);
  wire s152, sub152, and152, or152;
  wire b_inv152;
  assign b_inv152 = ~b152;
  assign s152  = a152 ^ b152 ^ c152;
  assign sub152 = a152 ^ b_inv152 ^ c152;
  assign and152 = a152 & b152;
  assign or152  = a152 | b152;
  assign c153 = (a152 & b152) | (a152 & c152) | (b152 & c152);
  wire c_sub153;
  assign c_sub153 = (a152 & b_inv152) | (a152 & c152) | (b_inv152 & c152);
  wire s153, sub153, and153, or153;
  wire b_inv153;
  assign b_inv153 = ~b153;
  assign s153  = a153 ^ b153 ^ c153;
  assign sub153 = a153 ^ b_inv153 ^ c153;
  assign and153 = a153 & b153;
  assign or153  = a153 | b153;
  assign c154 = (a153 & b153) | (a153 & c153) | (b153 & c153);
  wire c_sub154;
  assign c_sub154 = (a153 & b_inv153) | (a153 & c153) | (b_inv153 & c153);
  wire s154, sub154, and154, or154;
  wire b_inv154;
  assign b_inv154 = ~b154;
  assign s154  = a154 ^ b154 ^ c154;
  assign sub154 = a154 ^ b_inv154 ^ c154;
  assign and154 = a154 & b154;
  assign or154  = a154 | b154;
  assign c155 = (a154 & b154) | (a154 & c154) | (b154 & c154);
  wire c_sub155;
  assign c_sub155 = (a154 & b_inv154) | (a154 & c154) | (b_inv154 & c154);
  wire s155, sub155, and155, or155;
  wire b_inv155;
  assign b_inv155 = ~b155;
  assign s155  = a155 ^ b155 ^ c155;
  assign sub155 = a155 ^ b_inv155 ^ c155;
  assign and155 = a155 & b155;
  assign or155  = a155 | b155;
  assign c156 = (a155 & b155) | (a155 & c155) | (b155 & c155);
  wire c_sub156;
  assign c_sub156 = (a155 & b_inv155) | (a155 & c155) | (b_inv155 & c155);
  wire s156, sub156, and156, or156;
  wire b_inv156;
  assign b_inv156 = ~b156;
  assign s156  = a156 ^ b156 ^ c156;
  assign sub156 = a156 ^ b_inv156 ^ c156;
  assign and156 = a156 & b156;
  assign or156  = a156 | b156;
  assign c157 = (a156 & b156) | (a156 & c156) | (b156 & c156);
  wire c_sub157;
  assign c_sub157 = (a156 & b_inv156) | (a156 & c156) | (b_inv156 & c156);
  wire s157, sub157, and157, or157;
  wire b_inv157;
  assign b_inv157 = ~b157;
  assign s157  = a157 ^ b157 ^ c157;
  assign sub157 = a157 ^ b_inv157 ^ c157;
  assign and157 = a157 & b157;
  assign or157  = a157 | b157;
  assign c158 = (a157 & b157) | (a157 & c157) | (b157 & c157);
  wire c_sub158;
  assign c_sub158 = (a157 & b_inv157) | (a157 & c157) | (b_inv157 & c157);
  wire s158, sub158, and158, or158;
  wire b_inv158;
  assign b_inv158 = ~b158;
  assign s158  = a158 ^ b158 ^ c158;
  assign sub158 = a158 ^ b_inv158 ^ c158;
  assign and158 = a158 & b158;
  assign or158  = a158 | b158;
  assign c159 = (a158 & b158) | (a158 & c158) | (b158 & c158);
  wire c_sub159;
  assign c_sub159 = (a158 & b_inv158) | (a158 & c158) | (b_inv158 & c158);
  wire s159, sub159, and159, or159;
  wire b_inv159;
  assign b_inv159 = ~b159;
  assign s159  = a159 ^ b159 ^ c159;
  assign sub159 = a159 ^ b_inv159 ^ c159;
  assign and159 = a159 & b159;
  assign or159  = a159 | b159;
  assign c160 = (a159 & b159) | (a159 & c159) | (b159 & c159);
  wire c_sub160;
  assign c_sub160 = (a159 & b_inv159) | (a159 & c159) | (b_inv159 & c159);
  wire s160, sub160, and160, or160;
  wire b_inv160;
  assign b_inv160 = ~b160;
  assign s160  = a160 ^ b160 ^ c160;
  assign sub160 = a160 ^ b_inv160 ^ c160;
  assign and160 = a160 & b160;
  assign or160  = a160 | b160;
  assign c161 = (a160 & b160) | (a160 & c160) | (b160 & c160);
  wire c_sub161;
  assign c_sub161 = (a160 & b_inv160) | (a160 & c160) | (b_inv160 & c160);
  wire s161, sub161, and161, or161;
  wire b_inv161;
  assign b_inv161 = ~b161;
  assign s161  = a161 ^ b161 ^ c161;
  assign sub161 = a161 ^ b_inv161 ^ c161;
  assign and161 = a161 & b161;
  assign or161  = a161 | b161;
  assign c162 = (a161 & b161) | (a161 & c161) | (b161 & c161);
  wire c_sub162;
  assign c_sub162 = (a161 & b_inv161) | (a161 & c161) | (b_inv161 & c161);
  wire s162, sub162, and162, or162;
  wire b_inv162;
  assign b_inv162 = ~b162;
  assign s162  = a162 ^ b162 ^ c162;
  assign sub162 = a162 ^ b_inv162 ^ c162;
  assign and162 = a162 & b162;
  assign or162  = a162 | b162;
  assign c163 = (a162 & b162) | (a162 & c162) | (b162 & c162);
  wire c_sub163;
  assign c_sub163 = (a162 & b_inv162) | (a162 & c162) | (b_inv162 & c162);
  wire s163, sub163, and163, or163;
  wire b_inv163;
  assign b_inv163 = ~b163;
  assign s163  = a163 ^ b163 ^ c163;
  assign sub163 = a163 ^ b_inv163 ^ c163;
  assign and163 = a163 & b163;
  assign or163  = a163 | b163;
  assign c164 = (a163 & b163) | (a163 & c163) | (b163 & c163);
  wire c_sub164;
  assign c_sub164 = (a163 & b_inv163) | (a163 & c163) | (b_inv163 & c163);
  wire s164, sub164, and164, or164;
  wire b_inv164;
  assign b_inv164 = ~b164;
  assign s164  = a164 ^ b164 ^ c164;
  assign sub164 = a164 ^ b_inv164 ^ c164;
  assign and164 = a164 & b164;
  assign or164  = a164 | b164;
  assign c165 = (a164 & b164) | (a164 & c164) | (b164 & c164);
  wire c_sub165;
  assign c_sub165 = (a164 & b_inv164) | (a164 & c164) | (b_inv164 & c164);
  wire s165, sub165, and165, or165;
  wire b_inv165;
  assign b_inv165 = ~b165;
  assign s165  = a165 ^ b165 ^ c165;
  assign sub165 = a165 ^ b_inv165 ^ c165;
  assign and165 = a165 & b165;
  assign or165  = a165 | b165;
  assign c166 = (a165 & b165) | (a165 & c165) | (b165 & c165);
  wire c_sub166;
  assign c_sub166 = (a165 & b_inv165) | (a165 & c165) | (b_inv165 & c165);
  wire s166, sub166, and166, or166;
  wire b_inv166;
  assign b_inv166 = ~b166;
  assign s166  = a166 ^ b166 ^ c166;
  assign sub166 = a166 ^ b_inv166 ^ c166;
  assign and166 = a166 & b166;
  assign or166  = a166 | b166;
  assign c167 = (a166 & b166) | (a166 & c166) | (b166 & c166);
  wire c_sub167;
  assign c_sub167 = (a166 & b_inv166) | (a166 & c166) | (b_inv166 & c166);
  wire s167, sub167, and167, or167;
  wire b_inv167;
  assign b_inv167 = ~b167;
  assign s167  = a167 ^ b167 ^ c167;
  assign sub167 = a167 ^ b_inv167 ^ c167;
  assign and167 = a167 & b167;
  assign or167  = a167 | b167;
  assign c168 = (a167 & b167) | (a167 & c167) | (b167 & c167);
  wire c_sub168;
  assign c_sub168 = (a167 & b_inv167) | (a167 & c167) | (b_inv167 & c167);
  wire s168, sub168, and168, or168;
  wire b_inv168;
  assign b_inv168 = ~b168;
  assign s168  = a168 ^ b168 ^ c168;
  assign sub168 = a168 ^ b_inv168 ^ c168;
  assign and168 = a168 & b168;
  assign or168  = a168 | b168;
  assign c169 = (a168 & b168) | (a168 & c168) | (b168 & c168);
  wire c_sub169;
  assign c_sub169 = (a168 & b_inv168) | (a168 & c168) | (b_inv168 & c168);
  wire s169, sub169, and169, or169;
  wire b_inv169;
  assign b_inv169 = ~b169;
  assign s169  = a169 ^ b169 ^ c169;
  assign sub169 = a169 ^ b_inv169 ^ c169;
  assign and169 = a169 & b169;
  assign or169  = a169 | b169;
  assign c170 = (a169 & b169) | (a169 & c169) | (b169 & c169);
  wire c_sub170;
  assign c_sub170 = (a169 & b_inv169) | (a169 & c169) | (b_inv169 & c169);
  wire s170, sub170, and170, or170;
  wire b_inv170;
  assign b_inv170 = ~b170;
  assign s170  = a170 ^ b170 ^ c170;
  assign sub170 = a170 ^ b_inv170 ^ c170;
  assign and170 = a170 & b170;
  assign or170  = a170 | b170;
  assign c171 = (a170 & b170) | (a170 & c170) | (b170 & c170);
  wire c_sub171;
  assign c_sub171 = (a170 & b_inv170) | (a170 & c170) | (b_inv170 & c170);
  wire s171, sub171, and171, or171;
  wire b_inv171;
  assign b_inv171 = ~b171;
  assign s171  = a171 ^ b171 ^ c171;
  assign sub171 = a171 ^ b_inv171 ^ c171;
  assign and171 = a171 & b171;
  assign or171  = a171 | b171;
  assign c172 = (a171 & b171) | (a171 & c171) | (b171 & c171);
  wire c_sub172;
  assign c_sub172 = (a171 & b_inv171) | (a171 & c171) | (b_inv171 & c171);
  wire s172, sub172, and172, or172;
  wire b_inv172;
  assign b_inv172 = ~b172;
  assign s172  = a172 ^ b172 ^ c172;
  assign sub172 = a172 ^ b_inv172 ^ c172;
  assign and172 = a172 & b172;
  assign or172  = a172 | b172;
  assign c173 = (a172 & b172) | (a172 & c172) | (b172 & c172);
  wire c_sub173;
  assign c_sub173 = (a172 & b_inv172) | (a172 & c172) | (b_inv172 & c172);
  wire s173, sub173, and173, or173;
  wire b_inv173;
  assign b_inv173 = ~b173;
  assign s173  = a173 ^ b173 ^ c173;
  assign sub173 = a173 ^ b_inv173 ^ c173;
  assign and173 = a173 & b173;
  assign or173  = a173 | b173;
  assign c174 = (a173 & b173) | (a173 & c173) | (b173 & c173);
  wire c_sub174;
  assign c_sub174 = (a173 & b_inv173) | (a173 & c173) | (b_inv173 & c173);
  wire s174, sub174, and174, or174;
  wire b_inv174;
  assign b_inv174 = ~b174;
  assign s174  = a174 ^ b174 ^ c174;
  assign sub174 = a174 ^ b_inv174 ^ c174;
  assign and174 = a174 & b174;
  assign or174  = a174 | b174;
  assign c175 = (a174 & b174) | (a174 & c174) | (b174 & c174);
  wire c_sub175;
  assign c_sub175 = (a174 & b_inv174) | (a174 & c174) | (b_inv174 & c174);
  wire s175, sub175, and175, or175;
  wire b_inv175;
  assign b_inv175 = ~b175;
  assign s175  = a175 ^ b175 ^ c175;
  assign sub175 = a175 ^ b_inv175 ^ c175;
  assign and175 = a175 & b175;
  assign or175  = a175 | b175;
  assign c176 = (a175 & b175) | (a175 & c175) | (b175 & c175);
  wire c_sub176;
  assign c_sub176 = (a175 & b_inv175) | (a175 & c175) | (b_inv175 & c175);
  wire s176, sub176, and176, or176;
  wire b_inv176;
  assign b_inv176 = ~b176;
  assign s176  = a176 ^ b176 ^ c176;
  assign sub176 = a176 ^ b_inv176 ^ c176;
  assign and176 = a176 & b176;
  assign or176  = a176 | b176;
  assign c177 = (a176 & b176) | (a176 & c176) | (b176 & c176);
  wire c_sub177;
  assign c_sub177 = (a176 & b_inv176) | (a176 & c176) | (b_inv176 & c176);
  wire s177, sub177, and177, or177;
  wire b_inv177;
  assign b_inv177 = ~b177;
  assign s177  = a177 ^ b177 ^ c177;
  assign sub177 = a177 ^ b_inv177 ^ c177;
  assign and177 = a177 & b177;
  assign or177  = a177 | b177;
  assign c178 = (a177 & b177) | (a177 & c177) | (b177 & c177);
  wire c_sub178;
  assign c_sub178 = (a177 & b_inv177) | (a177 & c177) | (b_inv177 & c177);
  wire s178, sub178, and178, or178;
  wire b_inv178;
  assign b_inv178 = ~b178;
  assign s178  = a178 ^ b178 ^ c178;
  assign sub178 = a178 ^ b_inv178 ^ c178;
  assign and178 = a178 & b178;
  assign or178  = a178 | b178;
  assign c179 = (a178 & b178) | (a178 & c178) | (b178 & c178);
  wire c_sub179;
  assign c_sub179 = (a178 & b_inv178) | (a178 & c178) | (b_inv178 & c178);
  wire s179, sub179, and179, or179;
  wire b_inv179;
  assign b_inv179 = ~b179;
  assign s179  = a179 ^ b179 ^ c179;
  assign sub179 = a179 ^ b_inv179 ^ c179;
  assign and179 = a179 & b179;
  assign or179  = a179 | b179;
  assign c180 = (a179 & b179) | (a179 & c179) | (b179 & c179);
  wire c_sub180;
  assign c_sub180 = (a179 & b_inv179) | (a179 & c179) | (b_inv179 & c179);
  wire s180, sub180, and180, or180;
  wire b_inv180;
  assign b_inv180 = ~b180;
  assign s180  = a180 ^ b180 ^ c180;
  assign sub180 = a180 ^ b_inv180 ^ c180;
  assign and180 = a180 & b180;
  assign or180  = a180 | b180;
  assign c181 = (a180 & b180) | (a180 & c180) | (b180 & c180);
  wire c_sub181;
  assign c_sub181 = (a180 & b_inv180) | (a180 & c180) | (b_inv180 & c180);
  wire s181, sub181, and181, or181;
  wire b_inv181;
  assign b_inv181 = ~b181;
  assign s181  = a181 ^ b181 ^ c181;
  assign sub181 = a181 ^ b_inv181 ^ c181;
  assign and181 = a181 & b181;
  assign or181  = a181 | b181;
  assign c182 = (a181 & b181) | (a181 & c181) | (b181 & c181);
  wire c_sub182;
  assign c_sub182 = (a181 & b_inv181) | (a181 & c181) | (b_inv181 & c181);
  wire s182, sub182, and182, or182;
  wire b_inv182;
  assign b_inv182 = ~b182;
  assign s182  = a182 ^ b182 ^ c182;
  assign sub182 = a182 ^ b_inv182 ^ c182;
  assign and182 = a182 & b182;
  assign or182  = a182 | b182;
  assign c183 = (a182 & b182) | (a182 & c182) | (b182 & c182);
  wire c_sub183;
  assign c_sub183 = (a182 & b_inv182) | (a182 & c182) | (b_inv182 & c182);
  wire s183, sub183, and183, or183;
  wire b_inv183;
  assign b_inv183 = ~b183;
  assign s183  = a183 ^ b183 ^ c183;
  assign sub183 = a183 ^ b_inv183 ^ c183;
  assign and183 = a183 & b183;
  assign or183  = a183 | b183;
  assign c184 = (a183 & b183) | (a183 & c183) | (b183 & c183);
  wire c_sub184;
  assign c_sub184 = (a183 & b_inv183) | (a183 & c183) | (b_inv183 & c183);
  wire s184, sub184, and184, or184;
  wire b_inv184;
  assign b_inv184 = ~b184;
  assign s184  = a184 ^ b184 ^ c184;
  assign sub184 = a184 ^ b_inv184 ^ c184;
  assign and184 = a184 & b184;
  assign or184  = a184 | b184;
  assign c185 = (a184 & b184) | (a184 & c184) | (b184 & c184);
  wire c_sub185;
  assign c_sub185 = (a184 & b_inv184) | (a184 & c184) | (b_inv184 & c184);
  wire s185, sub185, and185, or185;
  wire b_inv185;
  assign b_inv185 = ~b185;
  assign s185  = a185 ^ b185 ^ c185;
  assign sub185 = a185 ^ b_inv185 ^ c185;
  assign and185 = a185 & b185;
  assign or185  = a185 | b185;
  assign c186 = (a185 & b185) | (a185 & c185) | (b185 & c185);
  wire c_sub186;
  assign c_sub186 = (a185 & b_inv185) | (a185 & c185) | (b_inv185 & c185);
  wire s186, sub186, and186, or186;
  wire b_inv186;
  assign b_inv186 = ~b186;
  assign s186  = a186 ^ b186 ^ c186;
  assign sub186 = a186 ^ b_inv186 ^ c186;
  assign and186 = a186 & b186;
  assign or186  = a186 | b186;
  assign c187 = (a186 & b186) | (a186 & c186) | (b186 & c186);
  wire c_sub187;
  assign c_sub187 = (a186 & b_inv186) | (a186 & c186) | (b_inv186 & c186);
  wire s187, sub187, and187, or187;
  wire b_inv187;
  assign b_inv187 = ~b187;
  assign s187  = a187 ^ b187 ^ c187;
  assign sub187 = a187 ^ b_inv187 ^ c187;
  assign and187 = a187 & b187;
  assign or187  = a187 | b187;
  assign c188 = (a187 & b187) | (a187 & c187) | (b187 & c187);
  wire c_sub188;
  assign c_sub188 = (a187 & b_inv187) | (a187 & c187) | (b_inv187 & c187);
  wire s188, sub188, and188, or188;
  wire b_inv188;
  assign b_inv188 = ~b188;
  assign s188  = a188 ^ b188 ^ c188;
  assign sub188 = a188 ^ b_inv188 ^ c188;
  assign and188 = a188 & b188;
  assign or188  = a188 | b188;
  assign c189 = (a188 & b188) | (a188 & c188) | (b188 & c188);
  wire c_sub189;
  assign c_sub189 = (a188 & b_inv188) | (a188 & c188) | (b_inv188 & c188);
  wire s189, sub189, and189, or189;
  wire b_inv189;
  assign b_inv189 = ~b189;
  assign s189  = a189 ^ b189 ^ c189;
  assign sub189 = a189 ^ b_inv189 ^ c189;
  assign and189 = a189 & b189;
  assign or189  = a189 | b189;
  assign c190 = (a189 & b189) | (a189 & c189) | (b189 & c189);
  wire c_sub190;
  assign c_sub190 = (a189 & b_inv189) | (a189 & c189) | (b_inv189 & c189);
  wire s190, sub190, and190, or190;
  wire b_inv190;
  assign b_inv190 = ~b190;
  assign s190  = a190 ^ b190 ^ c190;
  assign sub190 = a190 ^ b_inv190 ^ c190;
  assign and190 = a190 & b190;
  assign or190  = a190 | b190;
  assign c191 = (a190 & b190) | (a190 & c190) | (b190 & c190);
  wire c_sub191;
  assign c_sub191 = (a190 & b_inv190) | (a190 & c190) | (b_inv190 & c190);
  wire s191, sub191, and191, or191;
  wire b_inv191;
  assign b_inv191 = ~b191;
  assign s191  = a191 ^ b191 ^ c191;
  assign sub191 = a191 ^ b_inv191 ^ c191;
  assign and191 = a191 & b191;
  assign or191  = a191 | b191;
  assign c192 = (a191 & b191) | (a191 & c191) | (b191 & c191);
  wire c_sub192;
  assign c_sub192 = (a191 & b_inv191) | (a191 & c191) | (b_inv191 & c191);
  wire s192, sub192, and192, or192;
  wire b_inv192;
  assign b_inv192 = ~b192;
  assign s192  = a192 ^ b192 ^ c192;
  assign sub192 = a192 ^ b_inv192 ^ c192;
  assign and192 = a192 & b192;
  assign or192  = a192 | b192;
  assign c193 = (a192 & b192) | (a192 & c192) | (b192 & c192);
  wire c_sub193;
  assign c_sub193 = (a192 & b_inv192) | (a192 & c192) | (b_inv192 & c192);
  wire s193, sub193, and193, or193;
  wire b_inv193;
  assign b_inv193 = ~b193;
  assign s193  = a193 ^ b193 ^ c193;
  assign sub193 = a193 ^ b_inv193 ^ c193;
  assign and193 = a193 & b193;
  assign or193  = a193 | b193;
  assign c194 = (a193 & b193) | (a193 & c193) | (b193 & c193);
  wire c_sub194;
  assign c_sub194 = (a193 & b_inv193) | (a193 & c193) | (b_inv193 & c193);
  wire s194, sub194, and194, or194;
  wire b_inv194;
  assign b_inv194 = ~b194;
  assign s194  = a194 ^ b194 ^ c194;
  assign sub194 = a194 ^ b_inv194 ^ c194;
  assign and194 = a194 & b194;
  assign or194  = a194 | b194;
  assign c195 = (a194 & b194) | (a194 & c194) | (b194 & c194);
  wire c_sub195;
  assign c_sub195 = (a194 & b_inv194) | (a194 & c194) | (b_inv194 & c194);
  wire s195, sub195, and195, or195;
  wire b_inv195;
  assign b_inv195 = ~b195;
  assign s195  = a195 ^ b195 ^ c195;
  assign sub195 = a195 ^ b_inv195 ^ c195;
  assign and195 = a195 & b195;
  assign or195  = a195 | b195;
  assign c196 = (a195 & b195) | (a195 & c195) | (b195 & c195);
  wire c_sub196;
  assign c_sub196 = (a195 & b_inv195) | (a195 & c195) | (b_inv195 & c195);
  wire s196, sub196, and196, or196;
  wire b_inv196;
  assign b_inv196 = ~b196;
  assign s196  = a196 ^ b196 ^ c196;
  assign sub196 = a196 ^ b_inv196 ^ c196;
  assign and196 = a196 & b196;
  assign or196  = a196 | b196;
  assign c197 = (a196 & b196) | (a196 & c196) | (b196 & c196);
  wire c_sub197;
  assign c_sub197 = (a196 & b_inv196) | (a196 & c196) | (b_inv196 & c196);
  wire s197, sub197, and197, or197;
  wire b_inv197;
  assign b_inv197 = ~b197;
  assign s197  = a197 ^ b197 ^ c197;
  assign sub197 = a197 ^ b_inv197 ^ c197;
  assign and197 = a197 & b197;
  assign or197  = a197 | b197;
  assign c198 = (a197 & b197) | (a197 & c197) | (b197 & c197);
  wire c_sub198;
  assign c_sub198 = (a197 & b_inv197) | (a197 & c197) | (b_inv197 & c197);
  wire s198, sub198, and198, or198;
  wire b_inv198;
  assign b_inv198 = ~b198;
  assign s198  = a198 ^ b198 ^ c198;
  assign sub198 = a198 ^ b_inv198 ^ c198;
  assign and198 = a198 & b198;
  assign or198  = a198 | b198;
  assign c199 = (a198 & b198) | (a198 & c198) | (b198 & c198);
  wire c_sub199;
  assign c_sub199 = (a198 & b_inv198) | (a198 & c198) | (b_inv198 & c198);
  wire s199, sub199, and199, or199;
  wire b_inv199;
  assign b_inv199 = ~b199;
  assign s199  = a199 ^ b199 ^ c199;
  assign sub199 = a199 ^ b_inv199 ^ c199;
  assign and199 = a199 & b199;
  assign or199  = a199 | b199;
  assign c200 = (a199 & b199) | (a199 & c199) | (b199 & c199);
  wire c_sub200;
  assign c_sub200 = (a199 & b_inv199) | (a199 & c199) | (b_inv199 & c199);
  wire s200, sub200, and200, or200;
  wire b_inv200;
  assign b_inv200 = ~b200;
  assign s200  = a200 ^ b200 ^ c200;
  assign sub200 = a200 ^ b_inv200 ^ c200;
  assign and200 = a200 & b200;
  assign or200  = a200 | b200;
  assign c201 = (a200 & b200) | (a200 & c200) | (b200 & c200);
  wire c_sub201;
  assign c_sub201 = (a200 & b_inv200) | (a200 & c200) | (b_inv200 & c200);
  wire s201, sub201, and201, or201;
  wire b_inv201;
  assign b_inv201 = ~b201;
  assign s201  = a201 ^ b201 ^ c201;
  assign sub201 = a201 ^ b_inv201 ^ c201;
  assign and201 = a201 & b201;
  assign or201  = a201 | b201;
  assign c202 = (a201 & b201) | (a201 & c201) | (b201 & c201);
  wire c_sub202;
  assign c_sub202 = (a201 & b_inv201) | (a201 & c201) | (b_inv201 & c201);
  wire s202, sub202, and202, or202;
  wire b_inv202;
  assign b_inv202 = ~b202;
  assign s202  = a202 ^ b202 ^ c202;
  assign sub202 = a202 ^ b_inv202 ^ c202;
  assign and202 = a202 & b202;
  assign or202  = a202 | b202;
  assign c203 = (a202 & b202) | (a202 & c202) | (b202 & c202);
  wire c_sub203;
  assign c_sub203 = (a202 & b_inv202) | (a202 & c202) | (b_inv202 & c202);
  wire s203, sub203, and203, or203;
  wire b_inv203;
  assign b_inv203 = ~b203;
  assign s203  = a203 ^ b203 ^ c203;
  assign sub203 = a203 ^ b_inv203 ^ c203;
  assign and203 = a203 & b203;
  assign or203  = a203 | b203;
  assign c204 = (a203 & b203) | (a203 & c203) | (b203 & c203);
  wire c_sub204;
  assign c_sub204 = (a203 & b_inv203) | (a203 & c203) | (b_inv203 & c203);
  wire s204, sub204, and204, or204;
  wire b_inv204;
  assign b_inv204 = ~b204;
  assign s204  = a204 ^ b204 ^ c204;
  assign sub204 = a204 ^ b_inv204 ^ c204;
  assign and204 = a204 & b204;
  assign or204  = a204 | b204;
  assign c205 = (a204 & b204) | (a204 & c204) | (b204 & c204);
  wire c_sub205;
  assign c_sub205 = (a204 & b_inv204) | (a204 & c204) | (b_inv204 & c204);
  wire s205, sub205, and205, or205;
  wire b_inv205;
  assign b_inv205 = ~b205;
  assign s205  = a205 ^ b205 ^ c205;
  assign sub205 = a205 ^ b_inv205 ^ c205;
  assign and205 = a205 & b205;
  assign or205  = a205 | b205;
  assign c206 = (a205 & b205) | (a205 & c205) | (b205 & c205);
  wire c_sub206;
  assign c_sub206 = (a205 & b_inv205) | (a205 & c205) | (b_inv205 & c205);
  wire s206, sub206, and206, or206;
  wire b_inv206;
  assign b_inv206 = ~b206;
  assign s206  = a206 ^ b206 ^ c206;
  assign sub206 = a206 ^ b_inv206 ^ c206;
  assign and206 = a206 & b206;
  assign or206  = a206 | b206;
  assign c207 = (a206 & b206) | (a206 & c206) | (b206 & c206);
  wire c_sub207;
  assign c_sub207 = (a206 & b_inv206) | (a206 & c206) | (b_inv206 & c206);
  wire s207, sub207, and207, or207;
  wire b_inv207;
  assign b_inv207 = ~b207;
  assign s207  = a207 ^ b207 ^ c207;
  assign sub207 = a207 ^ b_inv207 ^ c207;
  assign and207 = a207 & b207;
  assign or207  = a207 | b207;
  assign c208 = (a207 & b207) | (a207 & c207) | (b207 & c207);
  wire c_sub208;
  assign c_sub208 = (a207 & b_inv207) | (a207 & c207) | (b_inv207 & c207);
  wire s208, sub208, and208, or208;
  wire b_inv208;
  assign b_inv208 = ~b208;
  assign s208  = a208 ^ b208 ^ c208;
  assign sub208 = a208 ^ b_inv208 ^ c208;
  assign and208 = a208 & b208;
  assign or208  = a208 | b208;
  assign c209 = (a208 & b208) | (a208 & c208) | (b208 & c208);
  wire c_sub209;
  assign c_sub209 = (a208 & b_inv208) | (a208 & c208) | (b_inv208 & c208);
  wire s209, sub209, and209, or209;
  wire b_inv209;
  assign b_inv209 = ~b209;
  assign s209  = a209 ^ b209 ^ c209;
  assign sub209 = a209 ^ b_inv209 ^ c209;
  assign and209 = a209 & b209;
  assign or209  = a209 | b209;
  assign c210 = (a209 & b209) | (a209 & c209) | (b209 & c209);
  wire c_sub210;
  assign c_sub210 = (a209 & b_inv209) | (a209 & c209) | (b_inv209 & c209);
  wire s210, sub210, and210, or210;
  wire b_inv210;
  assign b_inv210 = ~b210;
  assign s210  = a210 ^ b210 ^ c210;
  assign sub210 = a210 ^ b_inv210 ^ c210;
  assign and210 = a210 & b210;
  assign or210  = a210 | b210;
  assign c211 = (a210 & b210) | (a210 & c210) | (b210 & c210);
  wire c_sub211;
  assign c_sub211 = (a210 & b_inv210) | (a210 & c210) | (b_inv210 & c210);
  wire s211, sub211, and211, or211;
  wire b_inv211;
  assign b_inv211 = ~b211;
  assign s211  = a211 ^ b211 ^ c211;
  assign sub211 = a211 ^ b_inv211 ^ c211;
  assign and211 = a211 & b211;
  assign or211  = a211 | b211;
  assign c212 = (a211 & b211) | (a211 & c211) | (b211 & c211);
  wire c_sub212;
  assign c_sub212 = (a211 & b_inv211) | (a211 & c211) | (b_inv211 & c211);
  wire s212, sub212, and212, or212;
  wire b_inv212;
  assign b_inv212 = ~b212;
  assign s212  = a212 ^ b212 ^ c212;
  assign sub212 = a212 ^ b_inv212 ^ c212;
  assign and212 = a212 & b212;
  assign or212  = a212 | b212;
  assign c213 = (a212 & b212) | (a212 & c212) | (b212 & c212);
  wire c_sub213;
  assign c_sub213 = (a212 & b_inv212) | (a212 & c212) | (b_inv212 & c212);
  wire s213, sub213, and213, or213;
  wire b_inv213;
  assign b_inv213 = ~b213;
  assign s213  = a213 ^ b213 ^ c213;
  assign sub213 = a213 ^ b_inv213 ^ c213;
  assign and213 = a213 & b213;
  assign or213  = a213 | b213;
  assign c214 = (a213 & b213) | (a213 & c213) | (b213 & c213);
  wire c_sub214;
  assign c_sub214 = (a213 & b_inv213) | (a213 & c213) | (b_inv213 & c213);
  wire s214, sub214, and214, or214;
  wire b_inv214;
  assign b_inv214 = ~b214;
  assign s214  = a214 ^ b214 ^ c214;
  assign sub214 = a214 ^ b_inv214 ^ c214;
  assign and214 = a214 & b214;
  assign or214  = a214 | b214;
  assign c215 = (a214 & b214) | (a214 & c214) | (b214 & c214);
  wire c_sub215;
  assign c_sub215 = (a214 & b_inv214) | (a214 & c214) | (b_inv214 & c214);
  wire s215, sub215, and215, or215;
  wire b_inv215;
  assign b_inv215 = ~b215;
  assign s215  = a215 ^ b215 ^ c215;
  assign sub215 = a215 ^ b_inv215 ^ c215;
  assign and215 = a215 & b215;
  assign or215  = a215 | b215;
  assign c216 = (a215 & b215) | (a215 & c215) | (b215 & c215);
  wire c_sub216;
  assign c_sub216 = (a215 & b_inv215) | (a215 & c215) | (b_inv215 & c215);
  wire s216, sub216, and216, or216;
  wire b_inv216;
  assign b_inv216 = ~b216;
  assign s216  = a216 ^ b216 ^ c216;
  assign sub216 = a216 ^ b_inv216 ^ c216;
  assign and216 = a216 & b216;
  assign or216  = a216 | b216;
  assign c217 = (a216 & b216) | (a216 & c216) | (b216 & c216);
  wire c_sub217;
  assign c_sub217 = (a216 & b_inv216) | (a216 & c216) | (b_inv216 & c216);
  wire s217, sub217, and217, or217;
  wire b_inv217;
  assign b_inv217 = ~b217;
  assign s217  = a217 ^ b217 ^ c217;
  assign sub217 = a217 ^ b_inv217 ^ c217;
  assign and217 = a217 & b217;
  assign or217  = a217 | b217;
  assign c218 = (a217 & b217) | (a217 & c217) | (b217 & c217);
  wire c_sub218;
  assign c_sub218 = (a217 & b_inv217) | (a217 & c217) | (b_inv217 & c217);
  wire s218, sub218, and218, or218;
  wire b_inv218;
  assign b_inv218 = ~b218;
  assign s218  = a218 ^ b218 ^ c218;
  assign sub218 = a218 ^ b_inv218 ^ c218;
  assign and218 = a218 & b218;
  assign or218  = a218 | b218;
  assign c219 = (a218 & b218) | (a218 & c218) | (b218 & c218);
  wire c_sub219;
  assign c_sub219 = (a218 & b_inv218) | (a218 & c218) | (b_inv218 & c218);
  wire s219, sub219, and219, or219;
  wire b_inv219;
  assign b_inv219 = ~b219;
  assign s219  = a219 ^ b219 ^ c219;
  assign sub219 = a219 ^ b_inv219 ^ c219;
  assign and219 = a219 & b219;
  assign or219  = a219 | b219;
  assign c220 = (a219 & b219) | (a219 & c219) | (b219 & c219);
  wire c_sub220;
  assign c_sub220 = (a219 & b_inv219) | (a219 & c219) | (b_inv219 & c219);
  wire s220, sub220, and220, or220;
  wire b_inv220;
  assign b_inv220 = ~b220;
  assign s220  = a220 ^ b220 ^ c220;
  assign sub220 = a220 ^ b_inv220 ^ c220;
  assign and220 = a220 & b220;
  assign or220  = a220 | b220;
  assign c221 = (a220 & b220) | (a220 & c220) | (b220 & c220);
  wire c_sub221;
  assign c_sub221 = (a220 & b_inv220) | (a220 & c220) | (b_inv220 & c220);
  wire s221, sub221, and221, or221;
  wire b_inv221;
  assign b_inv221 = ~b221;
  assign s221  = a221 ^ b221 ^ c221;
  assign sub221 = a221 ^ b_inv221 ^ c221;
  assign and221 = a221 & b221;
  assign or221  = a221 | b221;
  assign c222 = (a221 & b221) | (a221 & c221) | (b221 & c221);
  wire c_sub222;
  assign c_sub222 = (a221 & b_inv221) | (a221 & c221) | (b_inv221 & c221);
  wire s222, sub222, and222, or222;
  wire b_inv222;
  assign b_inv222 = ~b222;
  assign s222  = a222 ^ b222 ^ c222;
  assign sub222 = a222 ^ b_inv222 ^ c222;
  assign and222 = a222 & b222;
  assign or222  = a222 | b222;
  assign c223 = (a222 & b222) | (a222 & c222) | (b222 & c222);
  wire c_sub223;
  assign c_sub223 = (a222 & b_inv222) | (a222 & c222) | (b_inv222 & c222);
  wire s223, sub223, and223, or223;
  wire b_inv223;
  assign b_inv223 = ~b223;
  assign s223  = a223 ^ b223 ^ c223;
  assign sub223 = a223 ^ b_inv223 ^ c223;
  assign and223 = a223 & b223;
  assign or223  = a223 | b223;
  assign c224 = (a223 & b223) | (a223 & c223) | (b223 & c223);
  wire c_sub224;
  assign c_sub224 = (a223 & b_inv223) | (a223 & c223) | (b_inv223 & c223);
  wire s224, sub224, and224, or224;
  wire b_inv224;
  assign b_inv224 = ~b224;
  assign s224  = a224 ^ b224 ^ c224;
  assign sub224 = a224 ^ b_inv224 ^ c224;
  assign and224 = a224 & b224;
  assign or224  = a224 | b224;
  assign c225 = (a224 & b224) | (a224 & c224) | (b224 & c224);
  wire c_sub225;
  assign c_sub225 = (a224 & b_inv224) | (a224 & c224) | (b_inv224 & c224);
  wire s225, sub225, and225, or225;
  wire b_inv225;
  assign b_inv225 = ~b225;
  assign s225  = a225 ^ b225 ^ c225;
  assign sub225 = a225 ^ b_inv225 ^ c225;
  assign and225 = a225 & b225;
  assign or225  = a225 | b225;
  assign c226 = (a225 & b225) | (a225 & c225) | (b225 & c225);
  wire c_sub226;
  assign c_sub226 = (a225 & b_inv225) | (a225 & c225) | (b_inv225 & c225);
  wire s226, sub226, and226, or226;
  wire b_inv226;
  assign b_inv226 = ~b226;
  assign s226  = a226 ^ b226 ^ c226;
  assign sub226 = a226 ^ b_inv226 ^ c226;
  assign and226 = a226 & b226;
  assign or226  = a226 | b226;
  assign c227 = (a226 & b226) | (a226 & c226) | (b226 & c226);
  wire c_sub227;
  assign c_sub227 = (a226 & b_inv226) | (a226 & c226) | (b_inv226 & c226);
  wire s227, sub227, and227, or227;
  wire b_inv227;
  assign b_inv227 = ~b227;
  assign s227  = a227 ^ b227 ^ c227;
  assign sub227 = a227 ^ b_inv227 ^ c227;
  assign and227 = a227 & b227;
  assign or227  = a227 | b227;
  assign c228 = (a227 & b227) | (a227 & c227) | (b227 & c227);
  wire c_sub228;
  assign c_sub228 = (a227 & b_inv227) | (a227 & c227) | (b_inv227 & c227);
  wire s228, sub228, and228, or228;
  wire b_inv228;
  assign b_inv228 = ~b228;
  assign s228  = a228 ^ b228 ^ c228;
  assign sub228 = a228 ^ b_inv228 ^ c228;
  assign and228 = a228 & b228;
  assign or228  = a228 | b228;
  assign c229 = (a228 & b228) | (a228 & c228) | (b228 & c228);
  wire c_sub229;
  assign c_sub229 = (a228 & b_inv228) | (a228 & c228) | (b_inv228 & c228);
  wire s229, sub229, and229, or229;
  wire b_inv229;
  assign b_inv229 = ~b229;
  assign s229  = a229 ^ b229 ^ c229;
  assign sub229 = a229 ^ b_inv229 ^ c229;
  assign and229 = a229 & b229;
  assign or229  = a229 | b229;
  assign c230 = (a229 & b229) | (a229 & c229) | (b229 & c229);
  wire c_sub230;
  assign c_sub230 = (a229 & b_inv229) | (a229 & c229) | (b_inv229 & c229);
  wire s230, sub230, and230, or230;
  wire b_inv230;
  assign b_inv230 = ~b230;
  assign s230  = a230 ^ b230 ^ c230;
  assign sub230 = a230 ^ b_inv230 ^ c230;
  assign and230 = a230 & b230;
  assign or230  = a230 | b230;
  assign c231 = (a230 & b230) | (a230 & c230) | (b230 & c230);
  wire c_sub231;
  assign c_sub231 = (a230 & b_inv230) | (a230 & c230) | (b_inv230 & c230);
  wire s231, sub231, and231, or231;
  wire b_inv231;
  assign b_inv231 = ~b231;
  assign s231  = a231 ^ b231 ^ c231;
  assign sub231 = a231 ^ b_inv231 ^ c231;
  assign and231 = a231 & b231;
  assign or231  = a231 | b231;
  assign c232 = (a231 & b231) | (a231 & c231) | (b231 & c231);
  wire c_sub232;
  assign c_sub232 = (a231 & b_inv231) | (a231 & c231) | (b_inv231 & c231);
  wire s232, sub232, and232, or232;
  wire b_inv232;
  assign b_inv232 = ~b232;
  assign s232  = a232 ^ b232 ^ c232;
  assign sub232 = a232 ^ b_inv232 ^ c232;
  assign and232 = a232 & b232;
  assign or232  = a232 | b232;
  assign c233 = (a232 & b232) | (a232 & c232) | (b232 & c232);
  wire c_sub233;
  assign c_sub233 = (a232 & b_inv232) | (a232 & c232) | (b_inv232 & c232);
  wire s233, sub233, and233, or233;
  wire b_inv233;
  assign b_inv233 = ~b233;
  assign s233  = a233 ^ b233 ^ c233;
  assign sub233 = a233 ^ b_inv233 ^ c233;
  assign and233 = a233 & b233;
  assign or233  = a233 | b233;
  assign c234 = (a233 & b233) | (a233 & c233) | (b233 & c233);
  wire c_sub234;
  assign c_sub234 = (a233 & b_inv233) | (a233 & c233) | (b_inv233 & c233);
  wire s234, sub234, and234, or234;
  wire b_inv234;
  assign b_inv234 = ~b234;
  assign s234  = a234 ^ b234 ^ c234;
  assign sub234 = a234 ^ b_inv234 ^ c234;
  assign and234 = a234 & b234;
  assign or234  = a234 | b234;
  assign c235 = (a234 & b234) | (a234 & c234) | (b234 & c234);
  wire c_sub235;
  assign c_sub235 = (a234 & b_inv234) | (a234 & c234) | (b_inv234 & c234);
  wire s235, sub235, and235, or235;
  wire b_inv235;
  assign b_inv235 = ~b235;
  assign s235  = a235 ^ b235 ^ c235;
  assign sub235 = a235 ^ b_inv235 ^ c235;
  assign and235 = a235 & b235;
  assign or235  = a235 | b235;
  assign c236 = (a235 & b235) | (a235 & c235) | (b235 & c235);
  wire c_sub236;
  assign c_sub236 = (a235 & b_inv235) | (a235 & c235) | (b_inv235 & c235);
  wire s236, sub236, and236, or236;
  wire b_inv236;
  assign b_inv236 = ~b236;
  assign s236  = a236 ^ b236 ^ c236;
  assign sub236 = a236 ^ b_inv236 ^ c236;
  assign and236 = a236 & b236;
  assign or236  = a236 | b236;
  assign c237 = (a236 & b236) | (a236 & c236) | (b236 & c236);
  wire c_sub237;
  assign c_sub237 = (a236 & b_inv236) | (a236 & c236) | (b_inv236 & c236);
  wire s237, sub237, and237, or237;
  wire b_inv237;
  assign b_inv237 = ~b237;
  assign s237  = a237 ^ b237 ^ c237;
  assign sub237 = a237 ^ b_inv237 ^ c237;
  assign and237 = a237 & b237;
  assign or237  = a237 | b237;
  assign c238 = (a237 & b237) | (a237 & c237) | (b237 & c237);
  wire c_sub238;
  assign c_sub238 = (a237 & b_inv237) | (a237 & c237) | (b_inv237 & c237);
  wire s238, sub238, and238, or238;
  wire b_inv238;
  assign b_inv238 = ~b238;
  assign s238  = a238 ^ b238 ^ c238;
  assign sub238 = a238 ^ b_inv238 ^ c238;
  assign and238 = a238 & b238;
  assign or238  = a238 | b238;
  assign c239 = (a238 & b238) | (a238 & c238) | (b238 & c238);
  wire c_sub239;
  assign c_sub239 = (a238 & b_inv238) | (a238 & c238) | (b_inv238 & c238);
  wire s239, sub239, and239, or239;
  wire b_inv239;
  assign b_inv239 = ~b239;
  assign s239  = a239 ^ b239 ^ c239;
  assign sub239 = a239 ^ b_inv239 ^ c239;
  assign and239 = a239 & b239;
  assign or239  = a239 | b239;
  assign c240 = (a239 & b239) | (a239 & c239) | (b239 & c239);
  wire c_sub240;
  assign c_sub240 = (a239 & b_inv239) | (a239 & c239) | (b_inv239 & c239);
  wire s240, sub240, and240, or240;
  wire b_inv240;
  assign b_inv240 = ~b240;
  assign s240  = a240 ^ b240 ^ c240;
  assign sub240 = a240 ^ b_inv240 ^ c240;
  assign and240 = a240 & b240;
  assign or240  = a240 | b240;
  assign c241 = (a240 & b240) | (a240 & c240) | (b240 & c240);
  wire c_sub241;
  assign c_sub241 = (a240 & b_inv240) | (a240 & c240) | (b_inv240 & c240);
  wire s241, sub241, and241, or241;
  wire b_inv241;
  assign b_inv241 = ~b241;
  assign s241  = a241 ^ b241 ^ c241;
  assign sub241 = a241 ^ b_inv241 ^ c241;
  assign and241 = a241 & b241;
  assign or241  = a241 | b241;
  assign c242 = (a241 & b241) | (a241 & c241) | (b241 & c241);
  wire c_sub242;
  assign c_sub242 = (a241 & b_inv241) | (a241 & c241) | (b_inv241 & c241);
  wire s242, sub242, and242, or242;
  wire b_inv242;
  assign b_inv242 = ~b242;
  assign s242  = a242 ^ b242 ^ c242;
  assign sub242 = a242 ^ b_inv242 ^ c242;
  assign and242 = a242 & b242;
  assign or242  = a242 | b242;
  assign c243 = (a242 & b242) | (a242 & c242) | (b242 & c242);
  wire c_sub243;
  assign c_sub243 = (a242 & b_inv242) | (a242 & c242) | (b_inv242 & c242);
  wire s243, sub243, and243, or243;
  wire b_inv243;
  assign b_inv243 = ~b243;
  assign s243  = a243 ^ b243 ^ c243;
  assign sub243 = a243 ^ b_inv243 ^ c243;
  assign and243 = a243 & b243;
  assign or243  = a243 | b243;
  assign c244 = (a243 & b243) | (a243 & c243) | (b243 & c243);
  wire c_sub244;
  assign c_sub244 = (a243 & b_inv243) | (a243 & c243) | (b_inv243 & c243);
  wire s244, sub244, and244, or244;
  wire b_inv244;
  assign b_inv244 = ~b244;
  assign s244  = a244 ^ b244 ^ c244;
  assign sub244 = a244 ^ b_inv244 ^ c244;
  assign and244 = a244 & b244;
  assign or244  = a244 | b244;
  assign c245 = (a244 & b244) | (a244 & c244) | (b244 & c244);
  wire c_sub245;
  assign c_sub245 = (a244 & b_inv244) | (a244 & c244) | (b_inv244 & c244);
  wire s245, sub245, and245, or245;
  wire b_inv245;
  assign b_inv245 = ~b245;
  assign s245  = a245 ^ b245 ^ c245;
  assign sub245 = a245 ^ b_inv245 ^ c245;
  assign and245 = a245 & b245;
  assign or245  = a245 | b245;
  assign c246 = (a245 & b245) | (a245 & c245) | (b245 & c245);
  wire c_sub246;
  assign c_sub246 = (a245 & b_inv245) | (a245 & c245) | (b_inv245 & c245);
  wire s246, sub246, and246, or246;
  wire b_inv246;
  assign b_inv246 = ~b246;
  assign s246  = a246 ^ b246 ^ c246;
  assign sub246 = a246 ^ b_inv246 ^ c246;
  assign and246 = a246 & b246;
  assign or246  = a246 | b246;
  assign c247 = (a246 & b246) | (a246 & c246) | (b246 & c246);
  wire c_sub247;
  assign c_sub247 = (a246 & b_inv246) | (a246 & c246) | (b_inv246 & c246);
  wire s247, sub247, and247, or247;
  wire b_inv247;
  assign b_inv247 = ~b247;
  assign s247  = a247 ^ b247 ^ c247;
  assign sub247 = a247 ^ b_inv247 ^ c247;
  assign and247 = a247 & b247;
  assign or247  = a247 | b247;
  assign c248 = (a247 & b247) | (a247 & c247) | (b247 & c247);
  wire c_sub248;
  assign c_sub248 = (a247 & b_inv247) | (a247 & c247) | (b_inv247 & c247);
  wire s248, sub248, and248, or248;
  wire b_inv248;
  assign b_inv248 = ~b248;
  assign s248  = a248 ^ b248 ^ c248;
  assign sub248 = a248 ^ b_inv248 ^ c248;
  assign and248 = a248 & b248;
  assign or248  = a248 | b248;
  assign c249 = (a248 & b248) | (a248 & c248) | (b248 & c248);
  wire c_sub249;
  assign c_sub249 = (a248 & b_inv248) | (a248 & c248) | (b_inv248 & c248);
  wire s249, sub249, and249, or249;
  wire b_inv249;
  assign b_inv249 = ~b249;
  assign s249  = a249 ^ b249 ^ c249;
  assign sub249 = a249 ^ b_inv249 ^ c249;
  assign and249 = a249 & b249;
  assign or249  = a249 | b249;
  assign c250 = (a249 & b249) | (a249 & c249) | (b249 & c249);
  wire c_sub250;
  assign c_sub250 = (a249 & b_inv249) | (a249 & c249) | (b_inv249 & c249);
  wire s250, sub250, and250, or250;
  wire b_inv250;
  assign b_inv250 = ~b250;
  assign s250  = a250 ^ b250 ^ c250;
  assign sub250 = a250 ^ b_inv250 ^ c250;
  assign and250 = a250 & b250;
  assign or250  = a250 | b250;
  assign c251 = (a250 & b250) | (a250 & c250) | (b250 & c250);
  wire c_sub251;
  assign c_sub251 = (a250 & b_inv250) | (a250 & c250) | (b_inv250 & c250);
  wire s251, sub251, and251, or251;
  wire b_inv251;
  assign b_inv251 = ~b251;
  assign s251  = a251 ^ b251 ^ c251;
  assign sub251 = a251 ^ b_inv251 ^ c251;
  assign and251 = a251 & b251;
  assign or251  = a251 | b251;
  assign c252 = (a251 & b251) | (a251 & c251) | (b251 & c251);
  wire c_sub252;
  assign c_sub252 = (a251 & b_inv251) | (a251 & c251) | (b_inv251 & c251);
  wire s252, sub252, and252, or252;
  wire b_inv252;
  assign b_inv252 = ~b252;
  assign s252  = a252 ^ b252 ^ c252;
  assign sub252 = a252 ^ b_inv252 ^ c252;
  assign and252 = a252 & b252;
  assign or252  = a252 | b252;
  assign c253 = (a252 & b252) | (a252 & c252) | (b252 & c252);
  wire c_sub253;
  assign c_sub253 = (a252 & b_inv252) | (a252 & c252) | (b_inv252 & c252);
  wire s253, sub253, and253, or253;
  wire b_inv253;
  assign b_inv253 = ~b253;
  assign s253  = a253 ^ b253 ^ c253;
  assign sub253 = a253 ^ b_inv253 ^ c253;
  assign and253 = a253 & b253;
  assign or253  = a253 | b253;
  assign c254 = (a253 & b253) | (a253 & c253) | (b253 & c253);
  wire c_sub254;
  assign c_sub254 = (a253 & b_inv253) | (a253 & c253) | (b_inv253 & c253);
  wire s254, sub254, and254, or254;
  wire b_inv254;
  assign b_inv254 = ~b254;
  assign s254  = a254 ^ b254 ^ c254;
  assign sub254 = a254 ^ b_inv254 ^ c254;
  assign and254 = a254 & b254;
  assign or254  = a254 | b254;
  assign c255 = (a254 & b254) | (a254 & c254) | (b254 & c254);
  wire c_sub255;
  assign c_sub255 = (a254 & b_inv254) | (a254 & c254) | (b_inv254 & c254);
  wire s255, sub255, and255, or255;
  wire b_inv255;
  assign b_inv255 = ~b255;
  assign s255  = a255 ^ b255 ^ c255;
  assign sub255 = a255 ^ b_inv255 ^ c255;
  assign and255 = a255 & b255;
  assign or255  = a255 | b255;
  assign c256 = (a255 & b255) | (a255 & c255) | (b255 & c255);
  wire c_sub256;
  assign c_sub256 = (a255 & b_inv255) | (a255 & c255) | (b_inv255 & c255);
  assign y0 = (add_sel & s0) | (sub_sel & sub0) | (and_sel & and0) | (or_sel & or0);
  assign y1 = (add_sel & s1) | (sub_sel & sub1) | (and_sel & and1) | (or_sel & or1);
  assign y2 = (add_sel & s2) | (sub_sel & sub2) | (and_sel & and2) | (or_sel & or2);
  assign y3 = (add_sel & s3) | (sub_sel & sub3) | (and_sel & and3) | (or_sel & or3);
  assign y4 = (add_sel & s4) | (sub_sel & sub4) | (and_sel & and4) | (or_sel & or4);
  assign y5 = (add_sel & s5) | (sub_sel & sub5) | (and_sel & and5) | (or_sel & or5);
  assign y6 = (add_sel & s6) | (sub_sel & sub6) | (and_sel & and6) | (or_sel & or6);
  assign y7 = (add_sel & s7) | (sub_sel & sub7) | (and_sel & and7) | (or_sel & or7);
  assign y8 = (add_sel & s8) | (sub_sel & sub8) | (and_sel & and8) | (or_sel & or8);
  assign y9 = (add_sel & s9) | (sub_sel & sub9) | (and_sel & and9) | (or_sel & or9);
  assign y10 = (add_sel & s10) | (sub_sel & sub10) | (and_sel & and10) | (or_sel & or10);
  assign y11 = (add_sel & s11) | (sub_sel & sub11) | (and_sel & and11) | (or_sel & or11);
  assign y12 = (add_sel & s12) | (sub_sel & sub12) | (and_sel & and12) | (or_sel & or12);
  assign y13 = (add_sel & s13) | (sub_sel & sub13) | (and_sel & and13) | (or_sel & or13);
  assign y14 = (add_sel & s14) | (sub_sel & sub14) | (and_sel & and14) | (or_sel & or14);
  assign y15 = (add_sel & s15) | (sub_sel & sub15) | (and_sel & and15) | (or_sel & or15);
  assign y16 = (add_sel & s16) | (sub_sel & sub16) | (and_sel & and16) | (or_sel & or16);
  assign y17 = (add_sel & s17) | (sub_sel & sub17) | (and_sel & and17) | (or_sel & or17);
  assign y18 = (add_sel & s18) | (sub_sel & sub18) | (and_sel & and18) | (or_sel & or18);
  assign y19 = (add_sel & s19) | (sub_sel & sub19) | (and_sel & and19) | (or_sel & or19);
  assign y20 = (add_sel & s20) | (sub_sel & sub20) | (and_sel & and20) | (or_sel & or20);
  assign y21 = (add_sel & s21) | (sub_sel & sub21) | (and_sel & and21) | (or_sel & or21);
  assign y22 = (add_sel & s22) | (sub_sel & sub22) | (and_sel & and22) | (or_sel & or22);
  assign y23 = (add_sel & s23) | (sub_sel & sub23) | (and_sel & and23) | (or_sel & or23);
  assign y24 = (add_sel & s24) | (sub_sel & sub24) | (and_sel & and24) | (or_sel & or24);
  assign y25 = (add_sel & s25) | (sub_sel & sub25) | (and_sel & and25) | (or_sel & or25);
  assign y26 = (add_sel & s26) | (sub_sel & sub26) | (and_sel & and26) | (or_sel & or26);
  assign y27 = (add_sel & s27) | (sub_sel & sub27) | (and_sel & and27) | (or_sel & or27);
  assign y28 = (add_sel & s28) | (sub_sel & sub28) | (and_sel & and28) | (or_sel & or28);
  assign y29 = (add_sel & s29) | (sub_sel & sub29) | (and_sel & and29) | (or_sel & or29);
  assign y30 = (add_sel & s30) | (sub_sel & sub30) | (and_sel & and30) | (or_sel & or30);
  assign y31 = (add_sel & s31) | (sub_sel & sub31) | (and_sel & and31) | (or_sel & or31);
  assign y32 = (add_sel & s32) | (sub_sel & sub32) | (and_sel & and32) | (or_sel & or32);
  assign y33 = (add_sel & s33) | (sub_sel & sub33) | (and_sel & and33) | (or_sel & or33);
  assign y34 = (add_sel & s34) | (sub_sel & sub34) | (and_sel & and34) | (or_sel & or34);
  assign y35 = (add_sel & s35) | (sub_sel & sub35) | (and_sel & and35) | (or_sel & or35);
  assign y36 = (add_sel & s36) | (sub_sel & sub36) | (and_sel & and36) | (or_sel & or36);
  assign y37 = (add_sel & s37) | (sub_sel & sub37) | (and_sel & and37) | (or_sel & or37);
  assign y38 = (add_sel & s38) | (sub_sel & sub38) | (and_sel & and38) | (or_sel & or38);
  assign y39 = (add_sel & s39) | (sub_sel & sub39) | (and_sel & and39) | (or_sel & or39);
  assign y40 = (add_sel & s40) | (sub_sel & sub40) | (and_sel & and40) | (or_sel & or40);
  assign y41 = (add_sel & s41) | (sub_sel & sub41) | (and_sel & and41) | (or_sel & or41);
  assign y42 = (add_sel & s42) | (sub_sel & sub42) | (and_sel & and42) | (or_sel & or42);
  assign y43 = (add_sel & s43) | (sub_sel & sub43) | (and_sel & and43) | (or_sel & or43);
  assign y44 = (add_sel & s44) | (sub_sel & sub44) | (and_sel & and44) | (or_sel & or44);
  assign y45 = (add_sel & s45) | (sub_sel & sub45) | (and_sel & and45) | (or_sel & or45);
  assign y46 = (add_sel & s46) | (sub_sel & sub46) | (and_sel & and46) | (or_sel & or46);
  assign y47 = (add_sel & s47) | (sub_sel & sub47) | (and_sel & and47) | (or_sel & or47);
  assign y48 = (add_sel & s48) | (sub_sel & sub48) | (and_sel & and48) | (or_sel & or48);
  assign y49 = (add_sel & s49) | (sub_sel & sub49) | (and_sel & and49) | (or_sel & or49);
  assign y50 = (add_sel & s50) | (sub_sel & sub50) | (and_sel & and50) | (or_sel & or50);
  assign y51 = (add_sel & s51) | (sub_sel & sub51) | (and_sel & and51) | (or_sel & or51);
  assign y52 = (add_sel & s52) | (sub_sel & sub52) | (and_sel & and52) | (or_sel & or52);
  assign y53 = (add_sel & s53) | (sub_sel & sub53) | (and_sel & and53) | (or_sel & or53);
  assign y54 = (add_sel & s54) | (sub_sel & sub54) | (and_sel & and54) | (or_sel & or54);
  assign y55 = (add_sel & s55) | (sub_sel & sub55) | (and_sel & and55) | (or_sel & or55);
  assign y56 = (add_sel & s56) | (sub_sel & sub56) | (and_sel & and56) | (or_sel & or56);
  assign y57 = (add_sel & s57) | (sub_sel & sub57) | (and_sel & and57) | (or_sel & or57);
  assign y58 = (add_sel & s58) | (sub_sel & sub58) | (and_sel & and58) | (or_sel & or58);
  assign y59 = (add_sel & s59) | (sub_sel & sub59) | (and_sel & and59) | (or_sel & or59);
  assign y60 = (add_sel & s60) | (sub_sel & sub60) | (and_sel & and60) | (or_sel & or60);
  assign y61 = (add_sel & s61) | (sub_sel & sub61) | (and_sel & and61) | (or_sel & or61);
  assign y62 = (add_sel & s62) | (sub_sel & sub62) | (and_sel & and62) | (or_sel & or62);
  assign y63 = (add_sel & s63) | (sub_sel & sub63) | (and_sel & and63) | (or_sel & or63);
  assign y64 = (add_sel & s64) | (sub_sel & sub64) | (and_sel & and64) | (or_sel & or64);
  assign y65 = (add_sel & s65) | (sub_sel & sub65) | (and_sel & and65) | (or_sel & or65);
  assign y66 = (add_sel & s66) | (sub_sel & sub66) | (and_sel & and66) | (or_sel & or66);
  assign y67 = (add_sel & s67) | (sub_sel & sub67) | (and_sel & and67) | (or_sel & or67);
  assign y68 = (add_sel & s68) | (sub_sel & sub68) | (and_sel & and68) | (or_sel & or68);
  assign y69 = (add_sel & s69) | (sub_sel & sub69) | (and_sel & and69) | (or_sel & or69);
  assign y70 = (add_sel & s70) | (sub_sel & sub70) | (and_sel & and70) | (or_sel & or70);
  assign y71 = (add_sel & s71) | (sub_sel & sub71) | (and_sel & and71) | (or_sel & or71);
  assign y72 = (add_sel & s72) | (sub_sel & sub72) | (and_sel & and72) | (or_sel & or72);
  assign y73 = (add_sel & s73) | (sub_sel & sub73) | (and_sel & and73) | (or_sel & or73);
  assign y74 = (add_sel & s74) | (sub_sel & sub74) | (and_sel & and74) | (or_sel & or74);
  assign y75 = (add_sel & s75) | (sub_sel & sub75) | (and_sel & and75) | (or_sel & or75);
  assign y76 = (add_sel & s76) | (sub_sel & sub76) | (and_sel & and76) | (or_sel & or76);
  assign y77 = (add_sel & s77) | (sub_sel & sub77) | (and_sel & and77) | (or_sel & or77);
  assign y78 = (add_sel & s78) | (sub_sel & sub78) | (and_sel & and78) | (or_sel & or78);
  assign y79 = (add_sel & s79) | (sub_sel & sub79) | (and_sel & and79) | (or_sel & or79);
  assign y80 = (add_sel & s80) | (sub_sel & sub80) | (and_sel & and80) | (or_sel & or80);
  assign y81 = (add_sel & s81) | (sub_sel & sub81) | (and_sel & and81) | (or_sel & or81);
  assign y82 = (add_sel & s82) | (sub_sel & sub82) | (and_sel & and82) | (or_sel & or82);
  assign y83 = (add_sel & s83) | (sub_sel & sub83) | (and_sel & and83) | (or_sel & or83);
  assign y84 = (add_sel & s84) | (sub_sel & sub84) | (and_sel & and84) | (or_sel & or84);
  assign y85 = (add_sel & s85) | (sub_sel & sub85) | (and_sel & and85) | (or_sel & or85);
  assign y86 = (add_sel & s86) | (sub_sel & sub86) | (and_sel & and86) | (or_sel & or86);
  assign y87 = (add_sel & s87) | (sub_sel & sub87) | (and_sel & and87) | (or_sel & or87);
  assign y88 = (add_sel & s88) | (sub_sel & sub88) | (and_sel & and88) | (or_sel & or88);
  assign y89 = (add_sel & s89) | (sub_sel & sub89) | (and_sel & and89) | (or_sel & or89);
  assign y90 = (add_sel & s90) | (sub_sel & sub90) | (and_sel & and90) | (or_sel & or90);
  assign y91 = (add_sel & s91) | (sub_sel & sub91) | (and_sel & and91) | (or_sel & or91);
  assign y92 = (add_sel & s92) | (sub_sel & sub92) | (and_sel & and92) | (or_sel & or92);
  assign y93 = (add_sel & s93) | (sub_sel & sub93) | (and_sel & and93) | (or_sel & or93);
  assign y94 = (add_sel & s94) | (sub_sel & sub94) | (and_sel & and94) | (or_sel & or94);
  assign y95 = (add_sel & s95) | (sub_sel & sub95) | (and_sel & and95) | (or_sel & or95);
  assign y96 = (add_sel & s96) | (sub_sel & sub96) | (and_sel & and96) | (or_sel & or96);
  assign y97 = (add_sel & s97) | (sub_sel & sub97) | (and_sel & and97) | (or_sel & or97);
  assign y98 = (add_sel & s98) | (sub_sel & sub98) | (and_sel & and98) | (or_sel & or98);
  assign y99 = (add_sel & s99) | (sub_sel & sub99) | (and_sel & and99) | (or_sel & or99);
  assign y100 = (add_sel & s100) | (sub_sel & sub100) | (and_sel & and100) | (or_sel & or100);
  assign y101 = (add_sel & s101) | (sub_sel & sub101) | (and_sel & and101) | (or_sel & or101);
  assign y102 = (add_sel & s102) | (sub_sel & sub102) | (and_sel & and102) | (or_sel & or102);
  assign y103 = (add_sel & s103) | (sub_sel & sub103) | (and_sel & and103) | (or_sel & or103);
  assign y104 = (add_sel & s104) | (sub_sel & sub104) | (and_sel & and104) | (or_sel & or104);
  assign y105 = (add_sel & s105) | (sub_sel & sub105) | (and_sel & and105) | (or_sel & or105);
  assign y106 = (add_sel & s106) | (sub_sel & sub106) | (and_sel & and106) | (or_sel & or106);
  assign y107 = (add_sel & s107) | (sub_sel & sub107) | (and_sel & and107) | (or_sel & or107);
  assign y108 = (add_sel & s108) | (sub_sel & sub108) | (and_sel & and108) | (or_sel & or108);
  assign y109 = (add_sel & s109) | (sub_sel & sub109) | (and_sel & and109) | (or_sel & or109);
  assign y110 = (add_sel & s110) | (sub_sel & sub110) | (and_sel & and110) | (or_sel & or110);
  assign y111 = (add_sel & s111) | (sub_sel & sub111) | (and_sel & and111) | (or_sel & or111);
  assign y112 = (add_sel & s112) | (sub_sel & sub112) | (and_sel & and112) | (or_sel & or112);
  assign y113 = (add_sel & s113) | (sub_sel & sub113) | (and_sel & and113) | (or_sel & or113);
  assign y114 = (add_sel & s114) | (sub_sel & sub114) | (and_sel & and114) | (or_sel & or114);
  assign y115 = (add_sel & s115) | (sub_sel & sub115) | (and_sel & and115) | (or_sel & or115);
  assign y116 = (add_sel & s116) | (sub_sel & sub116) | (and_sel & and116) | (or_sel & or116);
  assign y117 = (add_sel & s117) | (sub_sel & sub117) | (and_sel & and117) | (or_sel & or117);
  assign y118 = (add_sel & s118) | (sub_sel & sub118) | (and_sel & and118) | (or_sel & or118);
  assign y119 = (add_sel & s119) | (sub_sel & sub119) | (and_sel & and119) | (or_sel & or119);
  assign y120 = (add_sel & s120) | (sub_sel & sub120) | (and_sel & and120) | (or_sel & or120);
  assign y121 = (add_sel & s121) | (sub_sel & sub121) | (and_sel & and121) | (or_sel & or121);
  assign y122 = (add_sel & s122) | (sub_sel & sub122) | (and_sel & and122) | (or_sel & or122);
  assign y123 = (add_sel & s123) | (sub_sel & sub123) | (and_sel & and123) | (or_sel & or123);
  assign y124 = (add_sel & s124) | (sub_sel & sub124) | (and_sel & and124) | (or_sel & or124);
  assign y125 = (add_sel & s125) | (sub_sel & sub125) | (and_sel & and125) | (or_sel & or125);
  assign y126 = (add_sel & s126) | (sub_sel & sub126) | (and_sel & and126) | (or_sel & or126);
  assign y127 = (add_sel & s127) | (sub_sel & sub127) | (and_sel & and127) | (or_sel & or127);
  assign y128 = (add_sel & s128) | (sub_sel & sub128) | (and_sel & and128) | (or_sel & or128);
  assign y129 = (add_sel & s129) | (sub_sel & sub129) | (and_sel & and129) | (or_sel & or129);
  assign y130 = (add_sel & s130) | (sub_sel & sub130) | (and_sel & and130) | (or_sel & or130);
  assign y131 = (add_sel & s131) | (sub_sel & sub131) | (and_sel & and131) | (or_sel & or131);
  assign y132 = (add_sel & s132) | (sub_sel & sub132) | (and_sel & and132) | (or_sel & or132);
  assign y133 = (add_sel & s133) | (sub_sel & sub133) | (and_sel & and133) | (or_sel & or133);
  assign y134 = (add_sel & s134) | (sub_sel & sub134) | (and_sel & and134) | (or_sel & or134);
  assign y135 = (add_sel & s135) | (sub_sel & sub135) | (and_sel & and135) | (or_sel & or135);
  assign y136 = (add_sel & s136) | (sub_sel & sub136) | (and_sel & and136) | (or_sel & or136);
  assign y137 = (add_sel & s137) | (sub_sel & sub137) | (and_sel & and137) | (or_sel & or137);
  assign y138 = (add_sel & s138) | (sub_sel & sub138) | (and_sel & and138) | (or_sel & or138);
  assign y139 = (add_sel & s139) | (sub_sel & sub139) | (and_sel & and139) | (or_sel & or139);
  assign y140 = (add_sel & s140) | (sub_sel & sub140) | (and_sel & and140) | (or_sel & or140);
  assign y141 = (add_sel & s141) | (sub_sel & sub141) | (and_sel & and141) | (or_sel & or141);
  assign y142 = (add_sel & s142) | (sub_sel & sub142) | (and_sel & and142) | (or_sel & or142);
  assign y143 = (add_sel & s143) | (sub_sel & sub143) | (and_sel & and143) | (or_sel & or143);
  assign y144 = (add_sel & s144) | (sub_sel & sub144) | (and_sel & and144) | (or_sel & or144);
  assign y145 = (add_sel & s145) | (sub_sel & sub145) | (and_sel & and145) | (or_sel & or145);
  assign y146 = (add_sel & s146) | (sub_sel & sub146) | (and_sel & and146) | (or_sel & or146);
  assign y147 = (add_sel & s147) | (sub_sel & sub147) | (and_sel & and147) | (or_sel & or147);
  assign y148 = (add_sel & s148) | (sub_sel & sub148) | (and_sel & and148) | (or_sel & or148);
  assign y149 = (add_sel & s149) | (sub_sel & sub149) | (and_sel & and149) | (or_sel & or149);
  assign y150 = (add_sel & s150) | (sub_sel & sub150) | (and_sel & and150) | (or_sel & or150);
  assign y151 = (add_sel & s151) | (sub_sel & sub151) | (and_sel & and151) | (or_sel & or151);
  assign y152 = (add_sel & s152) | (sub_sel & sub152) | (and_sel & and152) | (or_sel & or152);
  assign y153 = (add_sel & s153) | (sub_sel & sub153) | (and_sel & and153) | (or_sel & or153);
  assign y154 = (add_sel & s154) | (sub_sel & sub154) | (and_sel & and154) | (or_sel & or154);
  assign y155 = (add_sel & s155) | (sub_sel & sub155) | (and_sel & and155) | (or_sel & or155);
  assign y156 = (add_sel & s156) | (sub_sel & sub156) | (and_sel & and156) | (or_sel & or156);
  assign y157 = (add_sel & s157) | (sub_sel & sub157) | (and_sel & and157) | (or_sel & or157);
  assign y158 = (add_sel & s158) | (sub_sel & sub158) | (and_sel & and158) | (or_sel & or158);
  assign y159 = (add_sel & s159) | (sub_sel & sub159) | (and_sel & and159) | (or_sel & or159);
  assign y160 = (add_sel & s160) | (sub_sel & sub160) | (and_sel & and160) | (or_sel & or160);
  assign y161 = (add_sel & s161) | (sub_sel & sub161) | (and_sel & and161) | (or_sel & or161);
  assign y162 = (add_sel & s162) | (sub_sel & sub162) | (and_sel & and162) | (or_sel & or162);
  assign y163 = (add_sel & s163) | (sub_sel & sub163) | (and_sel & and163) | (or_sel & or163);
  assign y164 = (add_sel & s164) | (sub_sel & sub164) | (and_sel & and164) | (or_sel & or164);
  assign y165 = (add_sel & s165) | (sub_sel & sub165) | (and_sel & and165) | (or_sel & or165);
  assign y166 = (add_sel & s166) | (sub_sel & sub166) | (and_sel & and166) | (or_sel & or166);
  assign y167 = (add_sel & s167) | (sub_sel & sub167) | (and_sel & and167) | (or_sel & or167);
  assign y168 = (add_sel & s168) | (sub_sel & sub168) | (and_sel & and168) | (or_sel & or168);
  assign y169 = (add_sel & s169) | (sub_sel & sub169) | (and_sel & and169) | (or_sel & or169);
  assign y170 = (add_sel & s170) | (sub_sel & sub170) | (and_sel & and170) | (or_sel & or170);
  assign y171 = (add_sel & s171) | (sub_sel & sub171) | (and_sel & and171) | (or_sel & or171);
  assign y172 = (add_sel & s172) | (sub_sel & sub172) | (and_sel & and172) | (or_sel & or172);
  assign y173 = (add_sel & s173) | (sub_sel & sub173) | (and_sel & and173) | (or_sel & or173);
  assign y174 = (add_sel & s174) | (sub_sel & sub174) | (and_sel & and174) | (or_sel & or174);
  assign y175 = (add_sel & s175) | (sub_sel & sub175) | (and_sel & and175) | (or_sel & or175);
  assign y176 = (add_sel & s176) | (sub_sel & sub176) | (and_sel & and176) | (or_sel & or176);
  assign y177 = (add_sel & s177) | (sub_sel & sub177) | (and_sel & and177) | (or_sel & or177);
  assign y178 = (add_sel & s178) | (sub_sel & sub178) | (and_sel & and178) | (or_sel & or178);
  assign y179 = (add_sel & s179) | (sub_sel & sub179) | (and_sel & and179) | (or_sel & or179);
  assign y180 = (add_sel & s180) | (sub_sel & sub180) | (and_sel & and180) | (or_sel & or180);
  assign y181 = (add_sel & s181) | (sub_sel & sub181) | (and_sel & and181) | (or_sel & or181);
  assign y182 = (add_sel & s182) | (sub_sel & sub182) | (and_sel & and182) | (or_sel & or182);
  assign y183 = (add_sel & s183) | (sub_sel & sub183) | (and_sel & and183) | (or_sel & or183);
  assign y184 = (add_sel & s184) | (sub_sel & sub184) | (and_sel & and184) | (or_sel & or184);
  assign y185 = (add_sel & s185) | (sub_sel & sub185) | (and_sel & and185) | (or_sel & or185);
  assign y186 = (add_sel & s186) | (sub_sel & sub186) | (and_sel & and186) | (or_sel & or186);
  assign y187 = (add_sel & s187) | (sub_sel & sub187) | (and_sel & and187) | (or_sel & or187);
  assign y188 = (add_sel & s188) | (sub_sel & sub188) | (and_sel & and188) | (or_sel & or188);
  assign y189 = (add_sel & s189) | (sub_sel & sub189) | (and_sel & and189) | (or_sel & or189);
  assign y190 = (add_sel & s190) | (sub_sel & sub190) | (and_sel & and190) | (or_sel & or190);
  assign y191 = (add_sel & s191) | (sub_sel & sub191) | (and_sel & and191) | (or_sel & or191);
  assign y192 = (add_sel & s192) | (sub_sel & sub192) | (and_sel & and192) | (or_sel & or192);
  assign y193 = (add_sel & s193) | (sub_sel & sub193) | (and_sel & and193) | (or_sel & or193);
  assign y194 = (add_sel & s194) | (sub_sel & sub194) | (and_sel & and194) | (or_sel & or194);
  assign y195 = (add_sel & s195) | (sub_sel & sub195) | (and_sel & and195) | (or_sel & or195);
  assign y196 = (add_sel & s196) | (sub_sel & sub196) | (and_sel & and196) | (or_sel & or196);
  assign y197 = (add_sel & s197) | (sub_sel & sub197) | (and_sel & and197) | (or_sel & or197);
  assign y198 = (add_sel & s198) | (sub_sel & sub198) | (and_sel & and198) | (or_sel & or198);
  assign y199 = (add_sel & s199) | (sub_sel & sub199) | (and_sel & and199) | (or_sel & or199);
  assign y200 = (add_sel & s200) | (sub_sel & sub200) | (and_sel & and200) | (or_sel & or200);
  assign y201 = (add_sel & s201) | (sub_sel & sub201) | (and_sel & and201) | (or_sel & or201);
  assign y202 = (add_sel & s202) | (sub_sel & sub202) | (and_sel & and202) | (or_sel & or202);
  assign y203 = (add_sel & s203) | (sub_sel & sub203) | (and_sel & and203) | (or_sel & or203);
  assign y204 = (add_sel & s204) | (sub_sel & sub204) | (and_sel & and204) | (or_sel & or204);
  assign y205 = (add_sel & s205) | (sub_sel & sub205) | (and_sel & and205) | (or_sel & or205);
  assign y206 = (add_sel & s206) | (sub_sel & sub206) | (and_sel & and206) | (or_sel & or206);
  assign y207 = (add_sel & s207) | (sub_sel & sub207) | (and_sel & and207) | (or_sel & or207);
  assign y208 = (add_sel & s208) | (sub_sel & sub208) | (and_sel & and208) | (or_sel & or208);
  assign y209 = (add_sel & s209) | (sub_sel & sub209) | (and_sel & and209) | (or_sel & or209);
  assign y210 = (add_sel & s210) | (sub_sel & sub210) | (and_sel & and210) | (or_sel & or210);
  assign y211 = (add_sel & s211) | (sub_sel & sub211) | (and_sel & and211) | (or_sel & or211);
  assign y212 = (add_sel & s212) | (sub_sel & sub212) | (and_sel & and212) | (or_sel & or212);
  assign y213 = (add_sel & s213) | (sub_sel & sub213) | (and_sel & and213) | (or_sel & or213);
  assign y214 = (add_sel & s214) | (sub_sel & sub214) | (and_sel & and214) | (or_sel & or214);
  assign y215 = (add_sel & s215) | (sub_sel & sub215) | (and_sel & and215) | (or_sel & or215);
  assign y216 = (add_sel & s216) | (sub_sel & sub216) | (and_sel & and216) | (or_sel & or216);
  assign y217 = (add_sel & s217) | (sub_sel & sub217) | (and_sel & and217) | (or_sel & or217);
  assign y218 = (add_sel & s218) | (sub_sel & sub218) | (and_sel & and218) | (or_sel & or218);
  assign y219 = (add_sel & s219) | (sub_sel & sub219) | (and_sel & and219) | (or_sel & or219);
  assign y220 = (add_sel & s220) | (sub_sel & sub220) | (and_sel & and220) | (or_sel & or220);
  assign y221 = (add_sel & s221) | (sub_sel & sub221) | (and_sel & and221) | (or_sel & or221);
  assign y222 = (add_sel & s222) | (sub_sel & sub222) | (and_sel & and222) | (or_sel & or222);
  assign y223 = (add_sel & s223) | (sub_sel & sub223) | (and_sel & and223) | (or_sel & or223);
  assign y224 = (add_sel & s224) | (sub_sel & sub224) | (and_sel & and224) | (or_sel & or224);
  assign y225 = (add_sel & s225) | (sub_sel & sub225) | (and_sel & and225) | (or_sel & or225);
  assign y226 = (add_sel & s226) | (sub_sel & sub226) | (and_sel & and226) | (or_sel & or226);
  assign y227 = (add_sel & s227) | (sub_sel & sub227) | (and_sel & and227) | (or_sel & or227);
  assign y228 = (add_sel & s228) | (sub_sel & sub228) | (and_sel & and228) | (or_sel & or228);
  assign y229 = (add_sel & s229) | (sub_sel & sub229) | (and_sel & and229) | (or_sel & or229);
  assign y230 = (add_sel & s230) | (sub_sel & sub230) | (and_sel & and230) | (or_sel & or230);
  assign y231 = (add_sel & s231) | (sub_sel & sub231) | (and_sel & and231) | (or_sel & or231);
  assign y232 = (add_sel & s232) | (sub_sel & sub232) | (and_sel & and232) | (or_sel & or232);
  assign y233 = (add_sel & s233) | (sub_sel & sub233) | (and_sel & and233) | (or_sel & or233);
  assign y234 = (add_sel & s234) | (sub_sel & sub234) | (and_sel & and234) | (or_sel & or234);
  assign y235 = (add_sel & s235) | (sub_sel & sub235) | (and_sel & and235) | (or_sel & or235);
  assign y236 = (add_sel & s236) | (sub_sel & sub236) | (and_sel & and236) | (or_sel & or236);
  assign y237 = (add_sel & s237) | (sub_sel & sub237) | (and_sel & and237) | (or_sel & or237);
  assign y238 = (add_sel & s238) | (sub_sel & sub238) | (and_sel & and238) | (or_sel & or238);
  assign y239 = (add_sel & s239) | (sub_sel & sub239) | (and_sel & and239) | (or_sel & or239);
  assign y240 = (add_sel & s240) | (sub_sel & sub240) | (and_sel & and240) | (or_sel & or240);
  assign y241 = (add_sel & s241) | (sub_sel & sub241) | (and_sel & and241) | (or_sel & or241);
  assign y242 = (add_sel & s242) | (sub_sel & sub242) | (and_sel & and242) | (or_sel & or242);
  assign y243 = (add_sel & s243) | (sub_sel & sub243) | (and_sel & and243) | (or_sel & or243);
  assign y244 = (add_sel & s244) | (sub_sel & sub244) | (and_sel & and244) | (or_sel & or244);
  assign y245 = (add_sel & s245) | (sub_sel & sub245) | (and_sel & and245) | (or_sel & or245);
  assign y246 = (add_sel & s246) | (sub_sel & sub246) | (and_sel & and246) | (or_sel & or246);
  assign y247 = (add_sel & s247) | (sub_sel & sub247) | (and_sel & and247) | (or_sel & or247);
  assign y248 = (add_sel & s248) | (sub_sel & sub248) | (and_sel & and248) | (or_sel & or248);
  assign y249 = (add_sel & s249) | (sub_sel & sub249) | (and_sel & and249) | (or_sel & or249);
  assign y250 = (add_sel & s250) | (sub_sel & sub250) | (and_sel & and250) | (or_sel & or250);
  assign y251 = (add_sel & s251) | (sub_sel & sub251) | (and_sel & and251) | (or_sel & or251);
  assign y252 = (add_sel & s252) | (sub_sel & sub252) | (and_sel & and252) | (or_sel & or252);
  assign y253 = (add_sel & s253) | (sub_sel & sub253) | (and_sel & and253) | (or_sel & or253);
  assign y254 = (add_sel & s254) | (sub_sel & sub254) | (and_sel & and254) | (or_sel & or254);
  assign y255 = (add_sel & s255) | (sub_sel & sub255) | (and_sel & and255) | (or_sel & or255);
endmodule