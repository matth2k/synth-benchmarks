module chkn (
    x0,
    x1,
    x2,
    x3,
    x4,
    x5,
    x6,
    x7,
    x8,
    x9,
    x10,
    x11,
    x12,
    x13,
    x14,
    x15,
    x16,
    x17,
    x18,
    x19,
    x20,
    x21,
    x22,
    x23,
    x24,
    x25,
    x26,
    x27,
    x28,
    y0,
    y1,
    y2,
    y3,
    y4,
    y5,
    y6
);
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 ;
  output y0, y1, y2, y3, y4, y5, y6;
  wire n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 ;
  assign n30  = x23 & ~x26;
  assign n31  = (x23 & ~x24) | (x23 & n30) | (~x24 & n30);
  assign n32  = ~x21 & n31;
  assign n33  = (x20 & ~x22) | (x20 & n32) | (~x22 & n32);
  assign n34  = ~x20 & n33;
  assign n35  = ~x18 & n34;
  assign n36  = ~x19 & n35;
  assign n37  = x14 & n36;
  assign n38  = (x16 & x17) | (x16 & n37) | (x17 & n37);
  assign n39  = ~x17 & n38;
  assign n40  = x2 & x13;
  assign n41  = (x11 & ~n39) | (x11 & n40) | (~n39 & n40);
  assign n42  = n39 & n41;
  assign n43  = (x13 & ~x16) | (x13 & n42) | (~x16 & n42);
  assign n44  = x11 & ~n42;
  assign n45  = (x13 & ~n43) | (x13 & n44) | (~n43 & n44);
  assign n46  = ~x4 & x15;
  assign n47  = (x12 & n45) | (x12 & n46) | (n45 & n46);
  assign n48  = ~n45 & n47;
  assign n49  = ~x22 & x26;
  assign n50  = (x21 & x23) | (x21 & n49) | (x23 & n49);
  assign n51  = ~x21 & n50;
  assign n52  = ~x19 & n51;
  assign n53  = (x18 & ~x20) | (x18 & n52) | (~x20 & n52);
  assign n54  = ~x18 & n53;
  assign n55  = x13 & x14;
  assign n56  = (x15 & x17) | (x15 & n55) | (x17 & n55);
  assign n57  = ~x17 & n56;
  assign n58  = x12 & n57;
  assign n59  = (x2 & x11) | (x2 & n58) | (x11 & n58);
  assign n60  = ~x2 & n59;
  assign n64  = (x16 & ~n54) | (x16 & n60) | (~n54 & n60);
  assign n61  = x12 | x14;
  assign n62  = x11 | x15;
  assign n63  = (~x12 & n61) | (~x12 & n62) | (n61 & n62);
  assign n65  = x16 & ~n63;
  assign n66  = (n54 & n64) | (n54 & n65) | (n64 & n65);
  assign n67  = ~x4 & n66;
  assign n79  = (x2 & x25) | (x2 & x26) | (x25 & x26);
  assign n80  = x24 | n79;
  assign n81  = x21 & ~n80;
  assign n82  = (x22 & x23) | (x22 & n81) | (x23 & n81);
  assign n83  = ~x23 & n82;
  assign n84  = ~x19 & n83;
  assign n85  = (x18 & ~x20) | (x18 & n84) | (~x20 & n84);
  assign n86  = ~x18 & n85;
  assign n87  = ~x17 & n86;
  assign n88  = (~x12 & x15) | (~x12 & n87) | (x15 & n87);
  assign n89  = x12 & ~n88;
  assign n90  = ~x12 & x15;
  assign n91  = (~x2 & n89) | (~x2 & n90) | (n89 & n90);
  assign n92  = n89 | n91;
  assign n93  = x16 & ~n92;
  assign n94  = x13 & ~n93;
  assign n95  = x13 | n90;
  assign n96  = ~n94 & n95;
  assign n97  = x11 & ~n96;
  assign n76  = x15 & x16;
  assign n77  = x12 | x13;
  assign n78  = (x15 & ~n76) | (x15 & n77) | (~n76 & n77);
  assign n98  = x2 & ~n78;
  assign n99  = x11 | n98;
  assign n100 = ~n97 & n99;
  assign n101 = x14 & ~n100;
  assign n68  = (~x12 & x13) | (~x12 & x15) | (x13 & x15);
  assign n69  = ~x15 & n68;
  assign n70  = (x12 & x16) | (x12 & n69) | (x16 & n69);
  assign n71  = (n68 & n69) | (n68 & n70) | (n69 & n70);
  assign n72  = ~x12 & x16;
  assign n73  = ~x15 & n72;
  assign n74  = x2 | n73;
  assign n75  = (n71 & n73) | (n71 & n74) | (n73 & n74);
  assign n102 = ~x11 & n75;
  assign n103 = x14 | n102;
  assign n104 = ~n101 & n103;
  assign n105 = x3 & n104;
  assign n106 = ~x4 & n105;
  assign n181 = x13 & x16;
  assign n182 = x15 & n181;
  assign n147 = ~x23 & x26;
  assign n148 = x22 | n147;
  assign n149 = ~x23 & x24;
  assign n150 = (x22 & n147) | (x22 & n149) | (n147 & n149);
  assign n151 = n148 & ~n150;
  assign n152 = ~x9 & x23;
  assign n153 = ~x22 & n152;
  assign n154 = x25 & ~n153;
  assign n155 = (n151 & n153) | (n151 & ~n154) | (n153 & ~n154);
  assign n172 = (x2 & x21) | (x2 & n155) | (x21 & n155);
  assign n163 = x9 & ~x22;
  assign n164 = x9 | x24;
  assign n165 = (x26 & n163) | (x26 & n164) | (n163 & n164);
  assign n166 = x2 & ~n165;
  assign n167 = x22 | n166;
  assign n168 = (~x24 & n166) | (~x24 & n167) | (n166 & n167);
  assign n169 = x23 & n168;
  assign n156 = x22 & x26;
  assign n157 = (x22 & ~x25) | (x22 & n156) | (~x25 & n156);
  assign n160 = (x9 & x24) | (x9 & n157) | (x24 & n157);
  assign n158 = (~x2 & x22) | (~x2 & x26) | (x22 & x26);
  assign n159 = n79 & ~n158;
  assign n161 = x24 & n159;
  assign n162 = (~x9 & n160) | (~x9 & n161) | (n160 & n161);
  assign n170 = x23 | n162;
  assign n171 = (~x23 & n169) | (~x23 & n170) | (n169 & n170);
  assign n173 = ~x21 & n171;
  assign n174 = (n155 & ~n172) | (n155 & n173) | (~n172 & n173);
  assign n134 = ~x9 & x26;
  assign n135 = ~x25 & n134;
  assign n136 = x2 & n135;
  assign n131 = x23 & x25;
  assign n132 = x26 & n131;
  assign n133 = (x26 & n30) | (x26 & ~n132) | (n30 & ~n132);
  assign n137 = ~x2 & n133;
  assign n138 = (x21 & n136) | (x21 & ~n137) | (n136 & ~n137);
  assign n144 = (x22 & x24) | (x22 & n138) | (x24 & n138);
  assign n139 = x2 | x26;
  assign n140 = x21 | n139;
  assign n141 = ~x23 & x25;
  assign n142 = (x24 & ~n140) | (x24 & n141) | (~n140 & n141);
  assign n143 = n140 & n142;
  assign n145 = ~x22 & n143;
  assign n146 = (n138 & ~n144) | (n138 & n145) | (~n144 & n145);
  assign n175 = n146 & ~n174;
  assign n176 = x19 | x20;
  assign n177 = (n174 & n175) | (n174 & ~n176) | (n175 & ~n176);
  assign n178 = x14 & ~x18;
  assign n179 = (x17 & n177) | (x17 & n178) | (n177 & n178);
  assign n180 = ~x17 & n179;
  assign n183 = x11 & n180;
  assign n184 = x9 & ~x11;
  assign n185 = (n182 & ~n183) | (n182 & n184) | (~n183 & n184);
  assign n110 = ~x11 & x16;
  assign n276 = (x13 & x14) | (x13 & x16) | (x14 & x16);
  assign n211 = ~x21 & x25;
  assign n234 = x2 & x21;
  assign n235 = (x24 & n211) | (x24 & ~n234) | (n211 & ~n234);
  assign n245 = x26 & ~n235;
  assign n236 = x21 & x25;
  assign n237 = x24 & n236;
  assign n238 = ~x24 & x25;
  assign n239 = ~x21 & x26;
  assign n240 = x25 | n239;
  assign n241 = ~n238 & n240;
  assign n242 = (~x2 & x16) | (~x2 & n241) | (x16 & n241);
  assign n210 = x24 & x26;
  assign n212 = (~x24 & n210) | (~x24 & n211) | (n210 & n211);
  assign n243 = (x2 & x16) | (x2 & n212) | (x16 & n212);
  assign n244 = n242 & n243;
  assign n246 = n237 | n244;
  assign n247 = (n235 & n245) | (n235 & ~n246) | (n245 & ~n246);
  assign n248 = x2 & ~x24;
  assign n249 = x21 & n248;
  assign n250 = (x23 & n247) | (x23 & ~n249) | (n247 & ~n249);
  assign n189 = x25 & x26;
  assign n231 = (~x21 & x24) | (~x21 & n140) | (x24 & n140);
  assign n232 = n189 & n231;
  assign n233 = (n140 & ~n189) | (n140 & n232) | (~n189 & n232);
  assign n251 = (x23 & ~n233) | (x23 & n249) | (~n233 & n249);
  assign n252 = n250 & ~n251;
  assign n270 = (x20 & x22) | (x20 & ~n252) | (x22 & ~n252);
  assign n253 = x2 & ~x26;
  assign n254 = x24 & ~n253;
  assign n255 = (x25 & ~n253) | (x25 & n254) | (~n253 & n254);
  assign n256 = x23 & ~n255;
  assign n267 = (x21 & ~x22) | (x21 & n256) | (~x22 & n256);
  assign n257 = (x23 & ~x24) | (x23 & x25) | (~x24 & x25);
  assign n258 = x25 & ~n257;
  assign n259 = (x24 & n147) | (x24 & n257) | (n147 & n257);
  assign n260 = (x23 & n258) | (x23 & ~n259) | (n258 & ~n259);
  assign n264 = (x2 & ~x22) | (x2 & n260) | (~x22 & n260);
  assign n261 = x24 | x26;
  assign n262 = (~x23 & x25) | (~x23 & n261) | (x25 & n261);
  assign n263 = x23 | n262;
  assign n265 = x2 | n263;
  assign n266 = (~n260 & n264) | (~n260 & n265) | (n264 & n265);
  assign n268 = x21 | n266;
  assign n269 = (~n256 & n267) | (~n256 & n268) | (n267 & n268);
  assign n271 = x20 | n269;
  assign n272 = (n252 & n270) | (n252 & n271) | (n270 & n271);
  assign n273 = x18 | n272;
  assign n274 = (~x17 & x19) | (~x17 & n273) | (x19 & n273);
  assign n275 = x17 | n274;
  assign n277 = (~x13 & x16) | (~x13 & n275) | (x16 & n275);
  assign n278 = n276 & n277;
  assign n279 = (~x14 & n276) | (~x14 & n278) | (n276 & n278);
  assign n280 = x11 & ~n279;
  assign n281 = (x15 & n110) | (x15 & ~n280) | (n110 & ~n280);
  assign n282 = x7 & ~n281;
  assign n199 = x25 & ~x26;
  assign n200 = (x24 & x26) | (x24 & ~n199) | (x26 & ~n199);
  assign n201 = x21 & n200;
  assign n197 = ~x25 & x26;
  assign n198 = (x24 & x26) | (x24 & n197) | (x26 & n197);
  assign n202 = x2 & n198;
  assign n203 = x21 | n202;
  assign n204 = ~n201 & n203;
  assign n216 = x23 & n204;
  assign n205 = x21 & ~x26;
  assign n206 = (x2 & x24) | (x2 & n205) | (x24 & n205);
  assign n207 = ~x24 & n206;
  assign n208 = x21 & x24;
  assign n209 = (x21 & ~n189) | (x21 & n208) | (~n189 & n208);
  assign n213 = (~x2 & x23) | (~x2 & n209) | (x23 & n209);
  assign n214 = ~x2 & n212;
  assign n215 = (~n209 & n213) | (~n209 & n214) | (n213 & n214);
  assign n217 = n207 | n215;
  assign n218 = (n204 & ~n216) | (n204 & n217) | (~n216 & n217);
  assign n219 = ~x22 & n218;
  assign n186 = (~x2 & x24) | (~x2 & x26) | (x24 & x26);
  assign n187 = x2 & n186;
  assign n188 = (x25 & n186) | (x25 & n187) | (n186 & n187);
  assign n190 = x25 | n139;
  assign n191 = (x23 & n189) | (x23 & n190) | (n189 & n190);
  assign n192 = x24 & n191;
  assign n193 = (~x24 & n190) | (~x24 & n192) | (n190 & n192);
  assign n194 = x22 & ~n193;
  assign n195 = x23 | n194;
  assign n196 = (~n188 & n194) | (~n188 & n195) | (n194 & n195);
  assign n220 = n196 | n219;
  assign n221 = (~x21 & n219) | (~x21 & n220) | (n219 & n220);
  assign n222 = x18 | x20;
  assign n223 = (x19 & n221) | (x19 & n222) | (n221 & n222);
  assign n224 = n221 & ~n223;
  assign n225 = x15 & n224;
  assign n226 = (x16 & x17) | (x16 & n225) | (x17 & n225);
  assign n227 = ~x17 & n226;
  assign n228 = x11 & x14;
  assign n229 = (x13 & ~n227) | (x13 & n228) | (~n227 & n228);
  assign n230 = n227 & n229;
  assign n283 = n230 | n282;
  assign n284 = (x6 & n282) | (x6 & n283) | (n282 & n283);
  assign n285 = x5 | n284;
  assign n286 = (~n185 & n284) | (~n185 & n285) | (n284 & n285);
  assign n289 = (x14 & ~x15) | (x14 & x16) | (~x15 & x16);
  assign n290 = (~x13 & x14) | (~x13 & x15) | (x14 & x15);
  assign n291 = ~n289 & n290;
  assign n292 = x5 & ~x11;
  assign n293 = (x9 & n291) | (x9 & n292) | (n291 & n292);
  assign n294 = ~x9 & n293;
  assign n287 = x14 & ~x15;
  assign n288 = ~x16 & n287;
  assign n295 = (x7 & n288) | (x7 & n294) | (n288 & n294);
  assign n296 = x13 & ~n295;
  assign n297 = (x13 & n294) | (x13 & ~n296) | (n294 & ~n296);
  assign n298 = (x12 & n286) | (x12 & n297) | (n286 & n297);
  assign n111 = (x11 & ~x15) | (x11 & x16) | (~x15 & x16);
  assign n112 = (x14 & n110) | (x14 & ~n111) | (n110 & ~n111);
  assign n113 = x5 & n112;
  assign n107 = (x6 & x14) | (x6 & x16) | (x14 & x16);
  assign n108 = x7 & x14;
  assign n109 = (~x16 & n107) | (~x16 & n108) | (n107 & n108);
  assign n114 = n109 | n113;
  assign n115 = (~x11 & n113) | (~x11 & n114) | (n113 & n114);
  assign n116 = (~x9 & x11) | (~x9 & x16) | (x11 & x16);
  assign n117 = (x9 & x11) | (x9 & ~x13) | (x11 & ~x13);
  assign n118 = n116 & ~n117;
  assign n126 = (~x5 & x14) | (~x5 & n118) | (x14 & n118);
  assign n119 = (~x13 & x15) | (~x13 & x16) | (x15 & x16);
  assign n120 = ~n111 & n119;
  assign n121 = x11 & ~x15;
  assign n122 = (x8 & x13) | (x8 & n121) | (x13 & n121);
  assign n123 = ~x13 & n122;
  assign n124 = x7 | n123;
  assign n125 = (n120 & n123) | (n120 & n124) | (n123 & n124);
  assign n127 = ~x14 & n125;
  assign n128 = (n118 & ~n126) | (n118 & n127) | (~n126 & n127);
  assign n129 = x13 | n128;
  assign n130 = (n115 & n128) | (n115 & n129) | (n128 & n129);
  assign n299 = (~x12 & n130) | (~x12 & n297) | (n130 & n297);
  assign n300 = n298 | n299;
  assign n303 = (x4 & ~x10) | (x4 & n300) | (~x10 & n300);
  assign n301 = x7 & x28;
  assign n302 = (x7 & x27) | (x7 & n301) | (x27 & n301);
  assign n304 = x10 & n302;
  assign n305 = (n300 & ~n303) | (n300 & n304) | (~n303 & n304);
  assign n306 = x14 & x15;
  assign n323 = ~x24 & n190;
  assign n324 = (n189 & n190) | (n189 & n323) | (n190 & n323);
  assign n325 = x22 & ~n324;
  assign n326 = ~x23 & n325;
  assign n327 = ~x20 & n326;
  assign n328 = (x19 & ~x21) | (x19 & n327) | (~x21 & n327);
  assign n329 = ~x19 & n328;
  assign n330 = x16 & ~x18;
  assign n331 = (x17 & n329) | (x17 & n330) | (n329 & n330);
  assign n332 = ~x17 & n331;
  assign n314 = x11 & x13;
  assign n333 = (x12 & n314) | (x12 & ~n332) | (n314 & ~n332);
  assign n334 = n332 & n333;
  assign n308 = x22 & n149;
  assign n309 = ~x20 & n308;
  assign n310 = (x19 & ~x21) | (x19 & n309) | (~x21 & n309);
  assign n311 = ~x19 & n310;
  assign n312 = x16 & ~x17;
  assign n313 = ~x18 & n312;
  assign n315 = (x12 & ~n313) | (x12 & n314) | (~n313 & n314);
  assign n316 = n313 & n315;
  assign n320 = (x9 & n311) | (x9 & ~n316) | (n311 & ~n316);
  assign n317 = x12 | x16;
  assign n318 = (~x11 & x13) | (~x11 & n317) | (x13 & n317);
  assign n319 = x11 | n318;
  assign n321 = x9 | n319;
  assign n322 = (~n311 & n320) | (~n311 & n321) | (n320 & n321);
  assign n335 = n322 | n334;
  assign n336 = (n306 & n334) | (n306 & ~n335) | (n334 & ~n335);
  assign n307 = (~x13 & n181) | (~x13 & n306) | (n181 & n306);
  assign n337 = (x12 & n307) | (x12 & ~n336) | (n307 & ~n336);
  assign n338 = x11 & n337;
  assign n339 = (x11 & n336) | (x11 & ~n338) | (n336 & ~n338);
  assign n340 = x0 & n339;
  assign n341 = ~x4 & n340;
  assign n342 = (~x12 & x14) | (~x12 & x15) | (x14 & x15);
  assign n343 = x16 & ~n342;
  assign n344 = (x12 & ~x16) | (x12 & n343) | (~x16 & n343);
  assign n345 = ~x13 & x16;
  assign n346 = x14 | x15;
  assign n347 = (x13 & n345) | (x13 & ~n346) | (n345 & ~n346);
  assign n348 = (x3 & x11) | (x3 & n90) | (x11 & n90);
  assign n349 = ~x3 & n348;
  assign n350 = (x15 & x16) | (x15 & ~n349) | (x16 & ~n349);
  assign n351 = x11 & ~n349;
  assign n352 = (~x16 & n350) | (~x16 & n351) | (n350 & n351);
  assign n383 = (~x13 & x14) | (~x13 & n352) | (x14 & n352);
  assign n353 = x22 & ~x23;
  assign n354 = ~x26 & n353;
  assign n355 = ~x3 & x21;
  assign n356 = (x2 & n354) | (x2 & n355) | (n354 & n355);
  assign n357 = ~x2 & n356;
  assign n358 = (x21 & x22) | (x21 & ~n357) | (x22 & ~n357);
  assign n359 = x23 & n358;
  assign n360 = (x23 & n357) | (x23 & ~n359) | (n357 & ~n359);
  assign n371 = (x20 & x24) | (x20 & n360) | (x24 & n360);
  assign n361 = x23 | x25;
  assign n362 = x24 | n361;
  assign n363 = x22 & ~n362;
  assign n364 = (x3 & x21) | (x3 & n363) | (x21 & n363);
  assign n365 = ~x3 & n364;
  assign n366 = (~x22 & x23) | (~x22 & n365) | (x23 & n365);
  assign n367 = x24 & ~n366;
  assign n368 = (x24 & n365) | (x24 & ~n367) | (n365 & ~n367);
  assign n369 = ~x26 & n368;
  assign n370 = (~x2 & n368) | (~x2 & n369) | (n368 & n369);
  assign n372 = ~x20 & n370;
  assign n373 = (n360 & ~n371) | (n360 & n372) | (~n371 & n372);
  assign n374 = ~x18 & n373;
  assign n375 = (x17 & ~x19) | (x17 & n374) | (~x19 & n374);
  assign n376 = ~x17 & n375;
  assign n377 = x12 & ~n376;
  assign n378 = x3 | x12;
  assign n379 = (~x15 & n377) | (~x15 & n378) | (n377 & n378);
  assign n380 = x11 & x16;
  assign n381 = (x13 & n379) | (x13 & n380) | (n379 & n380);
  assign n382 = ~n379 & n381;
  assign n384 = x14 & n382;
  assign n385 = (~n352 & n383) | (~n352 & n384) | (n383 & n384);
  assign n386 = (~n344 & n347) | (~n344 & n385) | (n347 & n385);
  assign n387 = x11 & ~n385;
  assign n388 = (n344 & n386) | (n344 & ~n387) | (n386 & ~n387);
  assign n389 = x1 & n388;
  assign n390 = ~x4 & n389;
  assign n393 = (x11 & ~x12) | (x11 & x14) | (~x12 & x14);
  assign n394 = ~x16 & n393;
  assign n395 = (~x12 & x16) | (~x12 & n394) | (x16 & n394);
  assign n391 = x12 & ~n182;
  assign n392 = (x11 & ~n182) | (x11 & n391) | (~n182 & n391);
  assign n443 = (~x4 & x11) | (~x4 & x14) | (x11 & x14);
  assign n444 = x12 & n443;
  assign n445 = (x4 & x12) | (x4 & ~n444) | (x12 & ~n444);
  assign n446 = (~x13 & x15) | (~x13 & n445) | (x15 & n445);
  assign n400 = x26 | n30;
  assign n401 = x25 | n400;
  assign n402 = (~x23 & n30) | (~x23 & n401) | (n30 & n401);
  assign n403 = (x24 & n30) | (x24 & n402) | (n30 & n402);
  assign n419 = ~x2 & n403;
  assign n404 = (x22 & x23) | (x22 & x24) | (x23 & x24);
  assign n405 = x22 & ~n190;
  assign n406 = (~x23 & n404) | (~x23 & n405) | (n404 & n405);
  assign n407 = ~x2 & x23;
  assign n408 = x24 & ~n407;
  assign n409 = (x22 & ~n407) | (x22 & n408) | (~n407 & n408);
  assign n416 = x25 & ~n409;
  assign n410 = (~x2 & x22) | (~x2 & x23) | (x22 & x23);
  assign n411 = x23 & ~x24;
  assign n412 = (~x22 & n410) | (~x22 & n411) | (n410 & n411);
  assign n413 = x24 | n189;
  assign n414 = x2 | x22;
  assign n415 = (~n189 & n413) | (~n189 & n414) | (n413 & n414);
  assign n417 = ~n412 & n415;
  assign n418 = (n409 & n416) | (n409 & n417) | (n416 & n417);
  assign n420 = ~n406 & n418;
  assign n421 = (~n403 & n419) | (~n403 & n420) | (n419 & n420);
  assign n422 = (x24 & ~n189) | (x24 & n237) | (~n189 & n237);
  assign n423 = x23 | n237;
  assign n424 = (n189 & n422) | (n189 & n423) | (n422 & n423);
  assign n432 = (x2 & x22) | (x2 & n424) | (x22 & n424);
  assign n425 = x2 & x25;
  assign n426 = x26 & ~n425;
  assign n427 = (x24 & ~n425) | (x24 & n426) | (~n425 & n426);
  assign n429 = (x21 & ~x23) | (x21 & n427) | (~x23 & n427);
  assign n428 = (x2 & ~x24) | (x2 & n253) | (~x24 & n253);
  assign n430 = x21 & n428;
  assign n431 = (~n427 & n429) | (~n427 & n430) | (n429 & n430);
  assign n433 = ~x22 & n431;
  assign n434 = (n424 & ~n432) | (n424 & n433) | (~n432 & n433);
  assign n435 = (x21 & n421) | (x21 & ~n434) | (n421 & ~n434);
  assign n396 = ~x22 & n139;
  assign n397 = (x25 & n139) | (x25 & n396) | (n139 & n396);
  assign n398 = x24 | n397;
  assign n399 = x23 | n398;
  assign n436 = (x21 & ~n399) | (x21 & n434) | (~n399 & n434);
  assign n437 = n435 & ~n436;
  assign n438 = (x19 & n222) | (x19 & ~n437) | (n222 & ~n437);
  assign n439 = n437 | n438;
  assign n440 = x11 & ~n439;
  assign n441 = (x14 & x17) | (x14 & n440) | (x17 & n440);
  assign n442 = ~x17 & n441;
  assign n447 = (x13 & ~x15) | (x13 & n442) | (~x15 & n442);
  assign n448 = n446 | n447;
  assign n449 = n392 | n448;
  assign n450 = n395 | n449;
  assign y0   = n48;
  assign y1   = n67;
  assign y2   = n106;
  assign y3   = n305;
  assign y4   = n341;
  assign y5   = n390;
  assign y6   = n450;
endmodule
