// IWLS benchmark module "C432.iscas" printed on Wed May 29 16:28:22 2002
module C432 (\1GAT(0) , \4GAT(1) , \8GAT(2) , \11GAT(3) , \14GAT(4) , \17GAT(5) , \21GAT(6) , \24GAT(7) , \27GAT(8) , \30GAT(9) , \34GAT(10) , \37GAT(11) , \40GAT(12) , \43GAT(13) , \47GAT(14) , \50GAT(15) , \53GAT(16) , \56GAT(17) , \60GAT(18) , \63GAT(19) , \66GAT(20) , \69GAT(21) , \73GAT(22) , \76GAT(23) , \79GAT(24) , \82GAT(25) , \86GAT(26) , \89GAT(27) , \92GAT(28) , \95GAT(29) , \99GAT(30) , \102GAT(31) , \105GAT(32) , \108GAT(33) , \112GAT(34) , \115GAT(35) , \223GAT(84) , \329GAT(133) , \370GAT(163) , \421GAT(188) , \430GAT(193) , \431GAT(194) , \432GAT(195) );
input
  \40GAT(12) ,
  \43GAT(13) ,
  \76GAT(23) ,
  \50GAT(15) ,
  \56GAT(17) ,
  \115GAT(35) ,
  \47GAT(14) ,
  \66GAT(20) ,
  \11GAT(3) ,
  \17GAT(5) ,
  \69GAT(21) ,
  \53GAT(16) ,
  \21GAT(6) ,
  \95GAT(29) ,
  \4GAT(1) ,
  \27GAT(8) ,
  \63GAT(19) ,
  \60GAT(18) ,
  \92GAT(28) ,
  \30GAT(9) ,
  \82GAT(25) ,
  \86GAT(26) ,
  \89GAT(27) ,
  \102GAT(31) ,
  \14GAT(4) ,
  \108GAT(33) ,
  \73GAT(22) ,
  \99GAT(30) ,
  \105GAT(32) ,
  \8GAT(2) ,
  \37GAT(11) ,
  \34GAT(10) ,
  \24GAT(7) ,
  \1GAT(0) ,
  \112GAT(34) ,
  \79GAT(24) ;
output
  \430GAT(193) ,
  \329GAT(133) ,
  \223GAT(84) ,
  \431GAT(194) ,
  \370GAT(163) ,
  \432GAT(195) ,
  \421GAT(188) ;
wire
  \151GAT(36) ,
  \150GAT(37) ,
  \224GAT(101) ,
  \127GAT(48) ,
  \126GAT(49) ,
  \419GAT(184) ,
  \273GAT(112) ,
  \159GAT(77) ,
  \189GAT(67) ,
  \348GAT(160) ,
  \336GAT(148) ,
  \375GAT(168) ,
  \246GAT(100) ,
  \263GAT(119) ,
  \158GAT(78) ,
  \282GAT(106) ,
  \414GAT(173) ,
  \188GAT(69) ,
  \407GAT(175) ,
  \233GAT(95) ,
  \357GAT(161) ,
  \411GAT(174) ,
  \334GAT(150) ,
  \[0] ,
  \295GAT(103) ,
  \[1] ,
  \289GAT(115) ,
  \343GAT(135) ,
  \333GAT(145) ,
  \[2] ,
  \379GAT(164) ,
  \[3] ,
  \399GAT(177) ,
  \264GAT(118) ,
  \[4] ,
  \342GAT(142) ,
  \404GAT(176) ,
  \242GAT(102) ,
  \[5] ,
  \381GAT(180) ,
  \356GAT(152) ,
  \162GAT(74) ,
  \373GAT(170) ,
  \[6] ,
  \353GAT(155) ,
  \418GAT(185) ,
  \307GAT(123) ,
  \171GAT(65) ,
  \332GAT(147) ,
  \303GAT(127) ,
  \374GAT(169) ,
  \345GAT(138) ,
  \319GAT(132) ,
  \428GAT(191) ,
  \270GAT(114) ,
  \230GAT(97) ,
  \213GAT(83) ,
  \239GAT(91) ,
  \296GAT(122) ,
  \236GAT(93) ,
  \294GAT(105) ,
  \300GAT(130) ,
  \350GAT(158) ,
  \199GAT(81) ,
  \154GAT(80) ,
  \165GAT(71) ,
  \378GAT(165) ,
  \344GAT(140) ,
  \174GAT(62) ,
  \180GAT(56) ,
  \285GAT(104) ,
  \279GAT(108) ,
  \380GAT(181) ,
  \417GAT(186) ,
  \331GAT(149) ,
  \309GAT(131) ,
  \119GAT(52) ,
  \118GAT(53) ,
  \425GAT(190) ,
  \306GAT(124) ,
  \341GAT(137) ,
  \335GAT(143) ,
  \302GAT(128) ,
  \251GAT(85) ,
  \196GAT(57) ,
  \195GAT(58) ,
  \276GAT(110) ,
  \259GAT(86) ,
  \293GAT(107) ,
  \377GAT(166) ,
  \258GAT(88) ,
  \360GAT(162) ,
  \339GAT(139) ,
  \429GAT(189) ,
  \393GAT(178) ,
  \143GAT(40) ,
  \142GAT(41) ,
  \346GAT(136) ,
  \198GAT(54) ,
  \168GAT(68) ,
  \247GAT(87) ,
  \351GAT(157) ,
  \338GAT(146) ,
  \197GAT(55) ,
  \340GAT(144) ,
  \123GAT(50) ,
  \122GAT(51) ,
  \203GAT(82) ,
  \254GAT(96) ,
  \354GAT(154) ,
  \260GAT(120) ,
  \422GAT(192) ,
  \191GAT(64) ,
  \192GAT(63) ,
  \193GAT(61) ,
  \305GAT(125) ,
  \243GAT(89) ,
  \292GAT(109) ,
  \301GAT(129) ,
  \147GAT(38) ,
  \146GAT(39) ,
  \288GAT(117) ,
  \376GAT(167) ,
  \371GAT(172) ,
  \290GAT(113) ,
  \386GAT(179) ,
  \257GAT(90) ,
  \194GAT(60) ,
  \304GAT(126) ,
  \352GAT(156) ,
  \416GAT(182) ,
  \190GAT(66) ,
  \227GAT(99) ,
  \187GAT(70) ,
  \139GAT(42) ,
  \138GAT(43) ,
  \420GAT(183) ,
  \256GAT(92) ,
  \250GAT(98) ,
  \415GAT(187) ,
  \349GAT(159) ,
  \267GAT(116) ,
  \337GAT(141) ,
  \330GAT(151) ,
  \255GAT(94) ,
  \185GAT(73) ,
  \291GAT(111) ,
  \131GAT(46) ,
  \130GAT(47) ,
  \186GAT(72) ,
  \355GAT(153) ,
  \183GAT(76) ,
  \184GAT(75) ,
  \135GAT(44) ,
  \134GAT(45) ,
  \372GAT(171) ,
  \347GAT(134) ,
  \157GAT(79) ,
  \177GAT(59) ,
  \308GAT(121) ;
assign
  \151GAT(36)  = ~\108GAT(33) ,
  \150GAT(37)  = ~\102GAT(31) ,
  \430GAT(193)  = \[4] ,
  \224GAT(101)  = (~\154GAT(80)  & \203GAT(82) ) | (\154GAT(80)  & ~\203GAT(82) ),
  \127GAT(48)  = ~\30GAT(9) ,
  \126GAT(49)  = ~\24GAT(7) ,
  \419GAT(184)  = ~\407GAT(175) ,
  \329GAT(133)  = \[1] ,
  \273GAT(112)  = ~\189GAT(67)  | ~\236GAT(93) ,
  \159GAT(77)  = ~\17GAT(5)  | ~\122GAT(51) ,
  \189GAT(67)  = ~\135GAT(44)  & ~\60GAT(18) ,
  \348GAT(160)  = ~\300GAT(130)  | ~\330GAT(151) ,
  \336GAT(148)  = ~\21GAT(6)  | ~\319GAT(132) ,
  \375GAT(168)  = ~\66GAT(20)  | ~\360GAT(162) ,
  \246GAT(100)  = ~\11GAT(3)  | ~\213GAT(83) ,
  \263GAT(119)  = ~\158GAT(78)  | ~\224GAT(101) ,
  \223GAT(84)  = \[0] ,
  \158GAT(78)  = ~\119GAT(52)  & ~\14GAT(4) ,
  \282GAT(106)  = ~\195GAT(58)  | ~\247GAT(87) ,
  \414GAT(173)  = ~\108GAT(33)  | (~\379GAT(164)  | (~\347GAT(134)  | ~\259GAT(86) )),
  \188GAT(69)  = ~\131GAT(46)  & ~\53GAT(16) ,
  \407GAT(175)  = ~\82GAT(25)  | (~\377GAT(166)  | (~\345GAT(138)  | ~\257GAT(90) )),
  \233GAT(95)  = (~\165GAT(71)  & \203GAT(82) ) | (\165GAT(71)  & ~\203GAT(82) ),
  \357GAT(161)  = \356GAT(152)  & (\355GAT(153)  & (\354GAT(154)  & (\353GAT(155)  & (\352GAT(156)  & (\351GAT(157)  & (\350GAT(158)  & (\349GAT(159)  & \348GAT(160) ))))))),
  \411GAT(174)  = ~\95GAT(29)  | (~\378GAT(165)  | (~\346GAT(136)  | ~\258GAT(88) )),
  \334GAT(150)  = ~\319GAT(132)  | ~\8GAT(2) ,
  \[0]  = ~\199GAT(81) ,
  \295GAT(103)  = ~\198GAT(54)  | ~\251GAT(85) ,
  \[1]  = ~\296GAT(122) ,
  \289GAT(115)  = ~\186GAT(72)  | ~\230GAT(97) ,
  \343GAT(135)  = (~\285GAT(104)  & \309GAT(131) ) | (\285GAT(104)  & ~\309GAT(131) ),
  \333GAT(145)  = (~\270GAT(114)  & \309GAT(131) ) | (\270GAT(114)  & ~\309GAT(131) ),
  \[2]  = ~\357GAT(161) ,
  \379GAT(164)  = ~\115GAT(35)  | ~\360GAT(162) ,
  \[3]  = ~\416GAT(182)  & ~\415GAT(187) ,
  \399GAT(177)  = ~\56GAT(17)  | (~\375GAT(168)  | (~\342GAT(142)  | ~\255GAT(94) )),
  \264GAT(118)  = ~\183GAT(76)  | ~\227GAT(99) ,
  \[4]  = ~\399GAT(177)  | (~\422GAT(192)  | (~\386GAT(179)  | ~\381GAT(180) )),
  \342GAT(142)  = ~\60GAT(18)  | ~\319GAT(132) ,
  \404GAT(176)  = ~\69GAT(21)  | (~\376GAT(167)  | (~\344GAT(140)  | ~\256GAT(92) )),
  \242GAT(102)  = ~\213GAT(83)  | ~\1GAT(0) ,
  \[5]  = ~\428GAT(191)  | (~\425GAT(190)  | (~\386GAT(179)  | ~\381GAT(180) )),
  \381GAT(180)  = ~\17GAT(5)  | (~\372GAT(171)  | (~\336GAT(148)  | ~\246GAT(100) )),
  \431GAT(194)  = \[5] ,
  \356GAT(152)  = ~\308GAT(121)  | ~\343GAT(135) ,
  \162GAT(74)  = ~\30GAT(9)  | ~\126GAT(49) ,
  \373GAT(170)  = ~\40GAT(12)  | ~\360GAT(162) ,
  \[6]  = ~\429GAT(189)  | (~\425GAT(190)  | (~\422GAT(192)  | ~\381GAT(180) )),
  \353GAT(155)  = ~\305GAT(125)  | ~\337GAT(141) ,
  \418GAT(185)  = ~\404GAT(176) ,
  \307GAT(123)  = ~\294GAT(105) ,
  \171GAT(65)  = ~\69GAT(21)  | ~\138GAT(43) ,
  \332GAT(147)  = (~\267GAT(116)  & \309GAT(131) ) | (\267GAT(116)  & ~\309GAT(131) ),
  \303GAT(127)  = ~\290GAT(113) ,
  \374GAT(169)  = ~\53GAT(16)  | ~\360GAT(162) ,
  \345GAT(138)  = ~\86GAT(26)  | ~\319GAT(132) ,
  \319GAT(132)  = ~\296GAT(122) ,
  \428GAT(191)  = ~\419GAT(184)  | (~\393GAT(178)  | ~\399GAT(177) ),
  \370GAT(163)  = \[2] ,
  \270GAT(114)  = ~\187GAT(70)  | ~\233GAT(95) ,
  \230GAT(97)  = (~\162GAT(74)  & \203GAT(82) ) | (\162GAT(74)  & ~\203GAT(82) ),
  \213GAT(83)  = ~\199GAT(81) ,
  \239GAT(91)  = (~\171GAT(65)  & \203GAT(82) ) | (\171GAT(65)  & ~\203GAT(82) ),
  \296GAT(122)  = \285GAT(104)  & (\282GAT(106)  & (\279GAT(108)  & (\276GAT(110)  & (\273GAT(112)  & (\270GAT(114)  & (\267GAT(116)  & (\264GAT(118)  & \260GAT(120) ))))))),
  \236GAT(93)  = (~\168GAT(68)  & \203GAT(82) ) | (\168GAT(68)  & ~\203GAT(82) ),
  \294GAT(105)  = ~\196GAT(57)  | ~\247GAT(87) ,
  \300GAT(130)  = ~\263GAT(119) ,
  \350GAT(158)  = ~\302GAT(128)  | ~\332GAT(147) ,
  \199GAT(81)  = \180GAT(56)  & (\177GAT(59)  & (\174GAT(62)  & (\171GAT(65)  & (\168GAT(68)  & (\165GAT(71)  & (\162GAT(74)  & (\159GAT(77)  & \154GAT(80) ))))))),
  \154GAT(80)  = ~\4GAT(1)  | ~\118GAT(53) ,
  \165GAT(71)  = ~\43GAT(13)  | ~\130GAT(47) ,
  \378GAT(165)  = ~\105GAT(32)  | ~\360GAT(162) ,
  \344GAT(140)  = ~\73GAT(22)  | ~\319GAT(132) ,
  \174GAT(62)  = ~\82GAT(25)  | ~\142GAT(41) ,
  \180GAT(56)  = ~\108GAT(33)  | ~\150GAT(37) ,
  \285GAT(104)  = ~\197GAT(55)  | ~\251GAT(85) ,
  \279GAT(108)  = ~\193GAT(61)  | ~\243GAT(89) ,
  \380GAT(181)  = ~\371GAT(172)  | (~\334GAT(150)  | (~\242GAT(102)  | ~\4GAT(1) )),
  \432GAT(195)  = \[6] ,
  \417GAT(186)  = ~\393GAT(178) ,
  \331GAT(149)  = (~\264GAT(118)  & \309GAT(131) ) | (\264GAT(118)  & ~\309GAT(131) ),
  \309GAT(131)  = ~\296GAT(122) ,
  \421GAT(188)  = \[3] ,
  \119GAT(52)  = ~\4GAT(1) ,
  \118GAT(53)  = ~\1GAT(0) ,
  \425GAT(190)  = ~\399GAT(177)  | (~\418GAT(185)  | (~\393GAT(178)  | ~\386GAT(179) )),
  \306GAT(124)  = ~\293GAT(107) ,
  \341GAT(137)  = (~\282GAT(106)  & \309GAT(131) ) | (\282GAT(106)  & ~\309GAT(131) ),
  \335GAT(143)  = (~\273GAT(112)  & \309GAT(131) ) | (\273GAT(112)  & ~\309GAT(131) ),
  \302GAT(128)  = ~\289GAT(115) ,
  \251GAT(85)  = (~\180GAT(56)  & \203GAT(82) ) | (\180GAT(56)  & ~\203GAT(82) ),
  \196GAT(57)  = ~\147GAT(38)  & ~\105GAT(32) ,
  \195GAT(58)  = ~\147GAT(38)  & ~\99GAT(30) ,
  \276GAT(110)  = ~\191GAT(64)  | ~\239GAT(91) ,
  \259GAT(86)  = ~\102GAT(31)  | ~\213GAT(83) ,
  \293GAT(107)  = ~\194GAT(60)  | ~\243GAT(89) ,
  \377GAT(166)  = ~\92GAT(28)  | ~\360GAT(162) ,
  \258GAT(88)  = ~\89GAT(27)  | ~\213GAT(83) ,
  \360GAT(162)  = ~\357GAT(161) ,
  \339GAT(139)  = (~\279GAT(108)  & \309GAT(131) ) | (\279GAT(108)  & ~\309GAT(131) ),
  \429GAT(189)  = ~\420GAT(183)  | (~\407GAT(175)  | (~\393GAT(178)  | ~\386GAT(179) )),
  \393GAT(178)  = ~\43GAT(13)  | (~\374GAT(169)  | (~\340GAT(144)  | ~\254GAT(96) )),
  \143GAT(40)  = ~\82GAT(25) ,
  \142GAT(41)  = ~\76GAT(23) ,
  \346GAT(136)  = ~\99GAT(30)  | ~\319GAT(132) ,
  \198GAT(54)  = ~\151GAT(36)  & ~\115GAT(35) ,
  \168GAT(68)  = ~\56GAT(17)  | ~\134GAT(45) ,
  \247GAT(87)  = (~\177GAT(59)  & \203GAT(82) ) | (\177GAT(59)  & ~\203GAT(82) ),
  \351GAT(157)  = ~\303GAT(127)  | ~\333GAT(145) ,
  \338GAT(146)  = ~\34GAT(10)  | ~\319GAT(132) ,
  \197GAT(55)  = ~\151GAT(36)  & ~\112GAT(34) ,
  \340GAT(144)  = ~\47GAT(14)  | ~\319GAT(132) ,
  \123GAT(50)  = ~\17GAT(5) ,
  \122GAT(51)  = ~\11GAT(3) ,
  \203GAT(82)  = ~\199GAT(81) ,
  \254GAT(96)  = ~\37GAT(11)  | ~\213GAT(83) ,
  \354GAT(154)  = ~\306GAT(124)  | ~\339GAT(139) ,
  \260GAT(120)  = ~\157GAT(79)  | ~\224GAT(101) ,
  \422GAT(192)  = ~\417GAT(186)  | ~\386GAT(179) ,
  \191GAT(64)  = ~\139GAT(42)  & ~\73GAT(22) ,
  \192GAT(63)  = ~\139GAT(42)  & ~\79GAT(24) ,
  \193GAT(61)  = ~\143GAT(40)  & ~\86GAT(26) ,
  \305GAT(125)  = ~\292GAT(109) ,
  \243GAT(89)  = (~\174GAT(62)  & \203GAT(82) ) | (\174GAT(62)  & ~\203GAT(82) ),
  \292GAT(109)  = ~\192GAT(63)  | ~\239GAT(91) ,
  \301GAT(129)  = ~\288GAT(117) ,
  \147GAT(38)  = ~\95GAT(29) ,
  \146GAT(39)  = ~\89GAT(27) ,
  \288GAT(117)  = ~\184GAT(75)  | ~\227GAT(99) ,
  \376GAT(167)  = ~\79GAT(24)  | ~\360GAT(162) ,
  \371GAT(172)  = ~\360GAT(162)  | ~\14GAT(4) ,
  \290GAT(113)  = ~\188GAT(69)  | ~\233GAT(95) ,
  \386GAT(179)  = ~\30GAT(9)  | (~\373GAT(170)  | (~\338GAT(146)  | ~\250GAT(98) )),
  \257GAT(90)  = ~\76GAT(23)  | ~\213GAT(83) ,
  \194GAT(60)  = ~\143GAT(40)  & ~\92GAT(28) ,
  \304GAT(126)  = ~\291GAT(111) ,
  \352GAT(156)  = ~\304GAT(126)  | ~\335GAT(143) ,
  \416GAT(182)  = \414GAT(173)  & (\411GAT(174)  & (\407GAT(175)  & (\404GAT(176)  & (\399GAT(177)  & (\393GAT(178)  & (\386GAT(179)  & \381GAT(180) )))))),
  \190GAT(66)  = ~\135GAT(44)  & ~\66GAT(20) ,
  \227GAT(99)  = (~\159GAT(77)  & \203GAT(82) ) | (\159GAT(77)  & ~\203GAT(82) ),
  \187GAT(70)  = ~\131GAT(46)  & ~\47GAT(14) ,
  \139GAT(42)  = ~\69GAT(21) ,
  \138GAT(43)  = ~\63GAT(19) ,
  \420GAT(183)  = ~\411GAT(174) ,
  \256GAT(92)  = ~\63GAT(19)  | ~\213GAT(83) ,
  \250GAT(98)  = ~\24GAT(7)  | ~\213GAT(83) ,
  \415GAT(187)  = ~\380GAT(181) ,
  \349GAT(159)  = ~\301GAT(129)  | ~\331GAT(149) ,
  \267GAT(116)  = ~\185GAT(73)  | ~\230GAT(97) ,
  \337GAT(141)  = (~\276GAT(110)  & \309GAT(131) ) | (\276GAT(110)  & ~\309GAT(131) ),
  \330GAT(151)  = (~\260GAT(120)  & \309GAT(131) ) | (\260GAT(120)  & ~\309GAT(131) ),
  \255GAT(94)  = ~\50GAT(15)  | ~\213GAT(83) ,
  \185GAT(73)  = ~\127GAT(48)  & ~\34GAT(10) ,
  \291GAT(111)  = ~\190GAT(66)  | ~\236GAT(93) ,
  \131GAT(46)  = ~\43GAT(13) ,
  \130GAT(47)  = ~\37GAT(11) ,
  \186GAT(72)  = ~\127GAT(48)  & ~\40GAT(12) ,
  \355GAT(153)  = ~\307GAT(123)  | ~\341GAT(137) ,
  \183GAT(76)  = ~\123GAT(50)  & ~\21GAT(6) ,
  \184GAT(75)  = ~\123GAT(50)  & ~\27GAT(8) ,
  \135GAT(44)  = ~\56GAT(17) ,
  \134GAT(45)  = ~\50GAT(15) ,
  \372GAT(171)  = ~\27GAT(8)  | ~\360GAT(162) ,
  \347GAT(134)  = ~\112GAT(34)  | ~\319GAT(132) ,
  \157GAT(79)  = ~\119GAT(52)  & ~\8GAT(2) ,
  \177GAT(59)  = ~\95GAT(29)  | ~\146GAT(39) ,
  \308GAT(121)  = ~\295GAT(103) ;
endmodule

