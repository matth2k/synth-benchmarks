// IWLS benchmark module "C7552.iscas" printed on Wed May 29 16:30:29 2002
module C7552 (\1(0) , \5(1) , \9(2) , \12(3) , \15(4) , \18(5) , \23(6) , \26(7) , \29(8) , \32(9) , \35(10) , \38(11) , \41(12) , \44(13) , \47(14) , \50(15) , \53(16) , \54(17) , \55(18) , \56(19) , \57(20) , \58(21) , \59(22) , \60(23) , \61(24) , \62(25) , \63(26) , \64(27) , \65(28) , \66(29) , \69(30) , \70(31) , \73(32) , \74(33) , \75(34) , \76(35) , \77(36) , \78(37) , \79(38) , \80(39) , \81(40) , \82(41) , \83(42) , \84(43) , \85(44) , \86(45) , \87(46) , \88(47) , \89(48) , \94(49) , \97(50) , \100(51) , \103(52) , \106(53) , \109(54) , \110(55) , \111(56) , \112(57) , \113(58) , \114(59) , \115(60) , \118(61) , \121(62) , \124(63) , \127(64) , \130(65) , \133(66) , \134(67) , \135(68) , \138(69) , \141(70) , \144(71) , \147(72) , \150(73) , \151(74) , \152(75) , \153(76) , \154(77) , \155(78) , \156(79) , \157(80) , \158(81) , \159(82) , \160(83) , \161(84) , \162(85) , \163(86) , \164(87) , \165(88) , \166(89) , \167(90) , \168(91) , \169(92) , \170(93) , \171(94) , \172(95) , \173(96) , \174(97) , \175(98) , \176(99) , \177(100) , \178(101) , \179(102) , \180(103) , \181(104) , \182(105) , \183(106) , \184(107) , \185(108) , \186(109) , \187(110) , \188(111) , \189(112) , \190(113) , \191(114) , \192(115) , \193(116) , \194(117) , \195(118) , \196(119) , \197(120) , \198(121) , \199(122) , \200(123) , \201(124) , \202(125) , \203(126) , \204(127) , \205(128) , \206(129) , \207(130) , \208(131) , \209(132) , \210(133) , \211(134) , \212(135) , \213(136) , \214(137) , \215(138) , \216(139) , \217(140) , \218(141) , \219(142) , \220(143) , \221(144) , \222(145) , \223(146) , \224(147) , \225(148) , \226(149) , \227(150) , \228(151) , \229(152) , \230(153) , \231(154) , \232(155) , \233(156) , \234(157) , \235(158) , \236(159) , \237(160) , \238(161) , \239(162) , \240(163) , \IN-339(164) , \1197(165) , \1455(166) , \1459(167) , \1462(168) , \1469(169) , \1480(170) , \1486(171) , \1492(172) , \1496(173) , \2204(174) , \2208(175) , \2211(176) , \2218(177) , \2224(178) , \2230(179) , \2236(180) , \2239(181) , \2247(182) , \2253(183) , \2256(184) , \3698(185) , \3701(186) , \3705(187) , \3711(188) , \3717(189) , \3723(190) , \3729(191) , \3737(192) , \3743(193) , \3749(194) , \4393(195) , \4394(196) , \4400(197) , \4405(198) , \4410(199) , \4415(200) , \4420(201) , \4427(202) , \4432(203) , \4437(204) , \4526(205) , \4528(206) , \339(164) , \2(313) , \3(312) , \450(288) , \448(284) , \444(282) , \442(280) , \440(277) , \438(274) , \496(271) , \494(267) , \492(265) , \490(263) , \488(260) , \486(258) , \484(256) , \482(253) , \480(250) , \560(248) , \542(246) , \558(244) , \556(242) , \554(240) , \552(238) , \550(236) , \548(234) , \546(232) , \544(230) , \540(227) , \538(224) , \536(222) , \534(220) , \532(218) , \530(216) , \528(214) , \526(212) , \524(210) , \279(304) , \436(286) , \478(269) , \522(226) , \402(395) , \404(390) , \406(388) , \408(385) , \410(387) , \432(428) , \446(393) , \284(384) , \286(419) , \289(383) , \292(392) , \341(420) , \281(547) , \453(596) , \278(536) , \373(2994) , \246(3110) , \258(3122) , \264(3121) , \270(3109) , \388(3093) , \391(3094) , \394(3095) , \397(3097) , \376(3206) , \379(3207) , \382(3148) , \385(3151) , \412(3369) , \414(3338) , \416(3368) , \249(3418) , \295(3352) , \324(3363) , \252(3450) , \276(3401) , \310(3393) , \313(3396) , \316(3397) , \319(3398) , \327(3408) , \330(3411) , \333(3416) , \336(3412) , \418(3449) , \273(3402) , \298(3387) , \301(3388) , \304(3390) , \307(3389) , \344(3382) , \422(3451) , \469(3452) , \419(3444) , \471(3445) , \359(3426) , \362(3429) , \365(3430) , \368(3431) , \347(3420) , \350(3421) , \353(3425) , \356(3424) , \321(3715) , \338(3716) , \370(3718) , \399(3717) );
input
  \4437(204) ,
  \200(123) ,
  \3743(193) ,
  \147(72) ,
  \158(81) ,
  \225(148) ,
  \169(92) ,
  \228(151) ,
  \106(53) ,
  \211(134) ,
  \183(106) ,
  \70(31) ,
  \12(3) ,
  \239(162) ,
  \81(40) ,
  \4420(201) ,
  \222(145) ,
  \197(120) ,
  \180(103) ,
  \109(54) ,
  \62(25) ,
  \73(32) ,
  \3729(191) ,
  \2218(177) ,
  \84(43) ,
  \2204(174) ,
  \236(159) ,
  \194(117) ,
  \54(17) ,
  \3701(186) ,
  \65(28) ,
  \1462(168) ,
  \76(35) ,
  \233(156) ,
  \150(73) ,
  \87(46) ,
  \191(114) ,
  \5(1) ,
  \208(131) ,
  \161(84) ,
  \35(10) ,
  \172(95) ,
  \3737(192) ,
  \57(20) ,
  \3723(190) ,
  \219(142) ,
  \230(153) ,
  \79(38) ,
  \3698(185) ,
  \177(100) ,
  \153(76) ,
  \164(87) ,
  \4528(206) ,
  \205(128) ,
  \38(11) ,
  \175(98) ,
  \112(57) ,
  \134(67) ,
  \216(139) ,
  \202(125) ,
  \156(79) ,
  \167(90) ,
  \1459(167) ,
  \185(108) ,
  \115(60) ,
  \213(136) ,
  \1492(172) ,
  \188(111) ,
  \159(82) ,
  \224(147) ,
  \199(122) ,
  \2256(184) ,
  \227(150) ,
  \182(105) ,
  \210(133) ,
  \60(23) ,
  \118(61) ,
  \238(161) ,
  \82(41) ,
  \221(144) ,
  \2253(183) ,
  \41(12) ,
  \29(8) ,
  \196(119) ,
  \3717(189) ,
  \63(26) ,
  \74(33) ,
  \85(44) ,
  \235(158) ,
  \193(116) ,
  \15(4) ,
  \4400(197) ,
  \44(13) ,
  \170(93) ,
  \55(18) ,
  \66(29) ,
  \232(155) ,
  \77(36) ,
  \151(74) ,
  \179(102) ,
  \88(47) ,
  \190(113) ,
  \2239(181) ,
  \207(130) ,
  \162(85) ,
  \3711(188) ,
  \1486(171) ,
  \23(6) ,
  \47(14) ,
  \173(96) ,
  \110(55) ,
  \58(21) ,
  \2211(176) ,
  \218(141) ,
  \121(62) ,
  \69(30) ,
  \1197(165) ,
  \2236(180) ,
  \154(77) ,
  \1(0) ,
  \240(163) ,
  \204(127) ,
  \165(88) ,
  \4427(202) ,
  \176(99) ,
  \4394(196) ,
  \113(58) ,
  \2247(182) ,
  \124(63) ,
  \215(138) ,
  \135(68) ,
  \201(124) ,
  \1480(170) ,
  \157(80) ,
  \168(91) ,
  \226(149) ,
  \IN-339(164) ,
  \229(152) ,
  \212(135) ,
  \184(107) ,
  \187(110) ,
  \127(64) ,
  \138(69) ,
  \80(39) ,
  \2230(179) ,
  \1469(169) ,
  \1455(166) ,
  \2208(175) ,
  \223(146) ,
  \198(121) ,
  \181(104) ,
  \50(15) ,
  \4405(198) ,
  \61(24) ,
  \4432(203) ,
  \3705(187) ,
  \32(9) ,
  \237(160) ,
  \220(143) ,
  \83(42) ,
  \94(49) ,
  \9(2) ,
  \195(118) ,
  \53(16) ,
  \64(27) ,
  \75(34) ,
  \234(157) ,
  \86(45) ,
  \192(115) ,
  \209(132) ,
  \97(50) ,
  \160(83) ,
  \171(94) ,
  \56(19) ,
  \130(65) ,
  \231(154) ,
  \78(37) ,
  \141(70) ,
  \152(75) ,
  \4410(199) ,
  \178(101) ,
  \89(48) ,
  \3749(194) ,
  \163(86) ,
  \206(129) ,
  \100(51) ,
  \174(97) ,
  \2224(178) ,
  \4415(200) ,
  \59(22) ,
  \111(56) ,
  \217(140) ,
  \18(5) ,
  \133(66) ,
  \1496(173) ,
  \144(71) ,
  \155(78) ,
  \203(126) ,
  \166(89) ,
  \4393(195) ,
  \4526(205) ,
  \103(52) ,
  \114(59) ,
  \186(109) ,
  \214(137) ,
  \189(112) ,
  \26(7) ;
output
  \336(3412) ,
  \492(265) ,
  \356(3424) ,
  \471(3445) ,
  \442(280) ,
  \276(3401) ,
  \298(3387) ,
  \284(384) ,
  \313(3396) ,
  \339(164) ,
  \550(236) ,
  \478(269) ,
  \270(3109) ,
  \450(288) ,
  \528(214) ,
  \419(3444) ,
  \385(3151) ,
  \373(2994) ,
  \249(3418) ,
  \359(3426) ,
  \292(392) ,
  \258(3122) ,
  \406(388) ,
  \3(312) ,
  \536(222) ,
  \522(226) ,
  \316(3397) ,
  \486(258) ,
  \436(286) ,
  \416(3368) ,
  \388(3093) ,
  \558(244) ,
  \289(383) ,
  \301(3388) ,
  \469(3452) ,
  \544(230) ,
  \494(267) ,
  \376(3206) ,
  \480(250) ,
  \530(216) ,
  \444(282) ,
  \281(547) ,
  \414(3338) ,
  \370(3718) ,
  \552(238) ,
  \347(3420) ,
  \319(3398) ,
  \327(3408) ,
  \246(3110) ,
  \304(3390) ,
  \362(3429) ,
  \344(3382) ,
  \560(248) ,
  \324(3363) ,
  \286(419) ,
  \379(3207) ,
  \408(385) ,
  \488(260) ,
  \278(536) ,
  \538(224) ,
  \338(3716) ,
  \391(3094) ,
  \252(3450) ,
  \524(210) ,
  \438(274) ,
  \422(3451) ,
  \2(313) ,
  \453(596) ,
  \365(3430) ,
  \496(271) ,
  \546(232) ,
  \482(253) ,
  \532(218) ,
  \307(3389) ,
  \264(3121) ,
  \330(3411) ,
  \341(420) ,
  \350(3421) ,
  \402(395) ,
  \554(240) ,
  \412(3369) ,
  \394(3095) ,
  \490(263) ,
  \410(387) ,
  \540(227) ,
  \440(277) ,
  \368(3431) ,
  \418(3449) ,
  \321(3715) ,
  \279(304) ,
  \333(3416) ,
  \446(393) ,
  \526(212) ,
  \353(3425) ,
  \295(3352) ,
  \382(3148) ,
  \273(3402) ,
  \310(3393) ,
  \397(3097) ,
  \548(234) ,
  \399(3717) ,
  \432(428) ,
  \534(220) ,
  \448(284) ,
  \484(256) ,
  \404(390) ,
  \556(242) ,
  \542(246) ;
wire
  \260(2889) ,
  \4872(2649) ,
  \5531(2823) ,
  \1514(406) ,
  \7117(3661) ,
  \7127(3660) ,
  \7050(2914) ,
  \5796(960) ,
  \1037(1561) ,
  \573(311) ,
  \7368(1627) ,
  \6732(1295) ,
  \5145(3488) ,
  \7548(1683) ,
  \4881(375) ,
  \5911(460) ,
  \7442(2814) ,
  \1143(3177) ,
  \6538(1055) ,
  \3228(2097) ,
  \2049(803) ,
  \4977(1835) ,
  \6269(2878) ,
  \980(3210) ,
  \3216(1462) ,
  \5753(354) ,
  \7070(3252) ,
  \4024(2268) ,
  \3119(2180) ,
  \2163(976) ,
  \4979(2200) ,
  \2501(2335) ,
  \5107(2690) ,
  \2149(808) ,
  \7538(1686) ,
  \4852(2352) ,
  \315(3281) ,
  \3471(2997) ,
  \1721(2410) ,
  \5682(2674) ,
  \4993(1203) ,
  \5937(2610) ,
  \3143(2738) ,
  \1239(1734) ,
  \4175(1007) ,
  \3079(1370) ,
  \1781(3684) ,
  \6535(984) ,
  \6458(1036) ,
  \6669(2767) ,
  \4250(2709) ,
  \6370(1065) ,
  \3249(2223) ,
  \5261(1447) ,
  \845(980) ,
  \4160(993) ,
  \5006(3226) ,
  \275(3286) ,
  \6498(1032) ,
  \2930(613) ,
  \2055(785) ,
  \4945(2743) ,
  \2343(1982) ,
  \2481(1721) ,
  \6103(3519) ,
  \5881(341) ,
  \4221(2171) ,
  \4983(1191) ,
  \1321(2460) ,
  \2872(430) ,
  \6972(2555) ,
  \621(532) ,
  \2925(514) ,
  \4291(2173) ,
  \2291(618) ,
  \577(631) ,
  \7567(1310) ,
  \2938(860) ,
  \6093(3463) ,
  \2511(2348) ,
  \7504(1150) ,
  \702(638) ,
  \2519(2361) ,
  \1372(522) ,
  \6213(3510) ,
  \6012(1287) ,
  \348(3371) ,
  \6968(2226) ,
  \4965(3227) ,
  \1597(1527) ,
  \6982(2565) ,
  \5780(1081) ,
  \5591(2952) ,
  \7272(1399) ,
  \7482(898) ,
  \6036(1383) ,
  \4341(1392) ,
  \6131(3149) ,
  \6952(2576) ,
  \4490(1000) ,
  \2226(264) ,
  \6173(1723) ,
  \1129(2434) ,
  \6896(1302) ,
  \4290(1911) ,
  \1092(1572) ,
  \7227(1358) ,
  \4239(2141) ,
  \6471(1307) ,
  \5138(3413) ,
  \4635(2727) ,
  \7228(1606) ,
  \395(3023) ,
  \3081(1641) ,
  \6884(1694) ,
  \6527(932) ,
  \2171(992) ,
  \3661(496) ,
  \6962(2572) ,
  \2546(3010) ,
  \6924(1613) ,
  \7471(902) ,
  \4716(2094) ,
  \2851(3008) ,
  \6163(3534) ,
  \1333(3069) ,
  \6347(3057) ,
  \5417(360) ,
  \3135(2868) ,
  \5718(3483) ,
  \4434(211) ,
  \5529(1519) ,
  \2852(2785) ,
  \1745(2084) ,
  \6978(2235) ,
  \4988(2834) ,
  \1198(299) ,
  \3151(2974) ,
  \1326(3135) ,
  \1902(1537) ,
  \4522(3128) ,
  \1735(2080) ,
  \7069(3323) ,
  \1725(2081) ,
  \1184(294) ,
  \6958(2248) ,
  \3351(1476) ,
  \7044(2590) ,
  \2789(2365) ,
  \5783(479) ,
  \3270(2892) ,
  \4179(1608) ,
  \4897(548) ,
  \4636(2976) ,
  \2849(3692) ,
  \5029(3114) ,
  \2839(3690) ,
  \6744(1601) ,
  \7291(1868) ,
  \1322(2847) ,
  \6357(3063) ,
  \4187(1884) ,
  \7009(3312) ,
  \7281(1860) ,
  \5007(1201) ,
  \2544(2919) ,
  \1226(1959) ,
  \4675(482) ,
  \6909(324) ,
  \3281(1464) ,
  \4911(507) ,
  \2914(591) ,
  \1320(2696) ,
  \328(3361) ,
  \7293(953) ,
  \6374(1420) ,
  \2564(2929) ,
  \4785(3237) ,
  \6153(3479) ,
  \1556(1807) ,
  \6614(1602) ,
  \1112(1553) ,
  \1546(1803) ,
  \4443(3309) ,
  \2117(577) ,
  \1572(1517) ,
  \4505(1014) ,
  \3745(231) ,
  \1369(646) ,
  \1300(2146) ,
  \4090(2757) ,
  \1206(306) ,
  \3019(1581) ,
  \4871(2985) ,
  \3444(2246) ,
  \5122(2443) ,
  \3376(1119) ,
  \5825(2383) ,
  \7185(3553) ,
  \3609(2984) ,
  \6631(334) ,
  \7138(2913) ,
  \3352(1773) ,
  \6240(2643) ,
  \5255(1092) ,
  \3282(1763) ,
  \3434(2230) ,
  \7562(1314) ,
  \4372(2520) ,
  \6509(1649) ,
  \2494(2333) ,
  \6009(345) ,
  \3488(2771) ,
  \5484(3103) ,
  \2532(2788) ,
  \3526(1610) ,
  \1125(2104) ,
  \6047(455) ,
  \7337(1902) ,
  \6220(2646) ,
  \2542(2786) ,
  \300(3267) ,
  \4760(2455) ,
  \1997(2944) ,
  \4904(1448) ,
  \3731(235) ,
  \2816(3019) ,
  \6589(435) ,
  \975(3157) ,
  \693(524) ,
  \6182(3065) ,
  \7286(1264) ,
  \6260(2636) ,
  \3567(1878) ,
  \7496(1516) ,
  \5183(498) ,
  \3608(2741) ,
  \2099(970) ,
  \6250(2638) ,
  \3622(407) ,
  \2854(2916) ,
  \2508(2630) ,
  \5776(1433) ,
  \6230(2633) ,
  \6294(2746) ,
  \1987(2942) ,
  \2768(2619) ,
  \587(402) ,
  \1776(3649) ,
  \6875(436) ,
  \1750(2078) ,
  \2753(2603) ,
  \5492(2402) ,
  \393(2937) ,
  \2571(3018) ,
  \5178(399) ,
  \1740(2071) ,
  \4585(1908) ,
  \4575(1909) ,
  \2520(2522) ,
  \2800(2530) ,
  \7490(887) ,
  \1766(3073) ,
  \7021(3475) ,
  \7081(3477) ,
  \2552(2794) ,
  \4680(683) ,
  \7256(1022) ,
  \2085(986) ,
  \3489(2906) ,
  \6598(1704) ,
  \4368(2855) ,
  \6702(1216) ,
  \363(3380) ,
  \1336(405) ,
  \5967(2796) ,
  \1014(560) ,
  \6856(1327) ,
  \5539(3104) ,
  \4745(3222) ,
  \5503(3465) ,
  \3469(2900) ,
  \4590(2499) ,
  \3061(1672) ,
  \3035(2374) ,
  \3479(2902) ,
  \3807(834) ,
  \5599(3107) ,
  \7396(1045) ,
  \1921(1832) ,
  \6992(3002) ,
  \7296(811) ,
  \5924(1382) ,
  \3051(1669) ,
  \6825(2469) ,
  \6658(2233) ,
  \7248(1668) ,
  \4485(711) ,
  \4149(742) ,
  \2616(1491) ,
  \3490(3195) ,
  \2124(731) ,
  \5836(2008) ,
  \4017(2569) ,
  \5761(357) ,
  \5447(487) ,
  \4496(999) ,
  \7469(1186) ,
  \5432(1242) ,
  \3033(2092) ,
  \3527(2160) ,
  \955(3172) ,
  \7100(3551) ,
  \1955(2073) ,
  \5521(3560) ,
  \2790(2526) ,
  \1965(2074) ,
  \1436(3029) ,
  \601(422) ,
  \6511(429) ,
  \4605(2405) ,
  \6057(1136) ,
  \6941(3141) ,
  \7060(3079) ,
  \989(3676) ,
  \4625(2678) ,
  \5210(1094) ,
  \3600(2838) ,
  \3279(3072) ,
  \6933(2908) ,
  \375(3090) ,
  \4567(2501) ,
  \4258(2716) ,
  \2272(594) ,
  \5175(372) ,
  \6788(1719) ,
  \5641(3583) ,
  \2749(2307) ,
  \2144(663) ,
  \2971(1744) ,
  \2058(654) ,
  \3130(2513) ,
  \5563(3481) ,
  \1170(3367) ,
  \4832(2597) ,
  \4919(605) ,
  \3658(681) ,
  \5482(2661) ,
  \1982(2816) ,
  \3695(1050) ,
  \7433(2949) ,
  \6241(3646) ,
  \1544(1148) ,
  \6567(319) ,
  \2143(806) ,
  \323(3238) ,
  \6973(3531) ,
  \3142(2478) ,
  \1960(2059) ,
  \3620(3117) ,
  \1503(303) ,
  \5840(2386) ,
  \7159(3377) ,
  \7172(2291) ,
  \2063(789) ,
  \5119(3175) ,
  \5952(2607) ,
  \1945(2019) ,
  \2296(715) ,
  \917(1190) ,
  \1281(1859) ,
  \2371(1788) ,
  \7145(3080) ,
  \7003(3247) ,
  \624(635) ,
  \3168(828) ,
  \3207(936) ,
  \710(642) ,
  \6070(2612) ,
  \7221(1020) ,
  \926(2163) ,
  \6251(3634) ,
  \997(2432) ,
  \4278(2739) ,
  \6853(318) ,
  \1024(1209) ,
  \2946(858) ,
  \5021(2960) ,
  \5112(2687) ,
  \2384(1132) ,
  \2005(2824) ,
  \5566(2000) ,
  \3559(2205) ,
  \3245(3230) ,
  \5570(2376) ,
  \707(544) ,
  \3548(1924) ,
  \3473(2759) ,
  \4520(3243) ,
  \3614(3044) ,
  \2819(3610) ,
  \711(852) ,
  \1992(2820) ,
  \2676(1994) ,
  \4276(2967) ,
  \5017(1219) ,
  \4058(3569) ,
  \4935(722) ,
  \7047(1485) ,
  \5420(1082) ,
  \1530(411) ,
  \4908(1096) ,
  \2286(554) ,
  \6083(3332) ,
  \1418(819) ,
  \4007(2231) ,
  \2158(677) ,
  \1157(1699) ,
  \5491(3269) ,
  \6514(397) ,
  \5892(1250) ,
  \984(3668) ,
  \6851(3120) ,
  \3926(1120) ,
  \2452(1506) ,
  \3854(1466) ,
  \337(3712) ,
  \7423(1687) ,
  \3909(1478) ,
  \6534(1408) ,
  \5576(2013) ,
  \6362(2849) ,
  \3558(1938) ,
  \7058(2912) ,
  \5425(363) ,
  \4255(2488) ,
  \3503(1221) ,
  \3465(3201) ,
  \1380(539) ,
  \7376(1599) ,
  \6953(3374) ,
  \6360(2697) ,
  \1234(1760) ,
  \1971(3165) ,
  \5061(3527) ,
  \6558(556) ,
  \3796(725) ,
  \3804(833) ,
  \3210(1026) ,
  \7000(2763) ,
  \6479(1339) ,
  \2220(266) ,
  \6223(3557) ,
  \5560(2396) ,
  \7383(1685) ,
  \5556(2024) ,
  \6439(1333) ,
  \5743(3647) ,
  \633(843) ,
  \4839(316) ,
  \6378(1066) ,
  \2863(3127) ,
  \4189(2176) ,
  \4764(2102) ,
  \6113(3574) ,
  \3786(568) ,
  \3799(799) ,
  \4146(743) ,
  \7618(2498) ,
  \5580(2390) ,
  \958(3228) ,
  \4493(998) ,
  \5855(1161) ,
  \5549(3268) ,
  \6768(1023) ,
  \5300(1052) ,
  \4141(690) ,
  \3855(1765) ,
  \7158(3251) ,
  \3449(2267) ,
  \4812(2269) ,
  \5546(2038) ,
  \4823(3327) ,
  \7506(1507) ,
  \1495(276) ,
  \6477(1639) ,
  \4488(752) ,
  \1224(1756) ,
  \3439(2252) ,
  \7245(1331) ,
  \1377(649) ,
  \346(3311) ,
  \1154(1928) ,
  \6655(2568) ,
  \2844(3625) ,
  \5197(501) ,
  \4086(3630) ,
  \5791(480) ,
  \5027(3053) ,
  \5672(2418) ,
  \2775(2803) ,
  \902(1199) ,
  \1867(1170) ,
  \6845(3058) ,
  \946(2122) ,
  \7385(1324) ,
  \6597(438) ,
  \296(3340) ,
  \7494(1164) ,
  \1999(2400) ,
  \4683(468) ,
  \7195(3606) ,
  \4720(2430) ,
  \5692(2413) ,
  \5465(885) ,
  \5748(1085) ,
  \2599(1786) ,
  \696(628) ,
  \1857(1169) ,
  \7573(1643) ,
  \5804(958) ,
  \941(2161) ,
  \3353(1972) ,
  \2878(386) ,
  \3283(1964) ,
  \4063(3570) ,
  \7182(2262) ,
  \1705(2010) ,
  \7299(1232) ,
  \956(2124) ,
  \1363(647) ,
  \5609(3277) ,
  \1156(1368) ,
  \6836(1833) ,
  \5071(3585) ,
  \4270(2459) ,
  \263(2858) ,
  \1175(3403) ,
  \2824(3611) ,
  \6017(346) ,
  \380(3086) ,
  \4474(759) ,
  \3214(1571) ,
  \3274(2999) ,
  \6883(439) ,
  \7192(2278) ,
  \3150(3241) ,
  \1940(2032) ,
  \7451(3123) ,
  \1607(1171) ,
  \5186(398) ,
  \7461(3125) ,
  \991(3405) ,
  \3666(698) ,
  \6610(1266) ,
  \907(1028) ,
  \5455(475) ,
  \3092(1888) ,
  \2701(1995) ,
  \1935(2004) ,
  \1136(3174) ,
  \6437(1187) ,
  \4743(3282) ,
  \5102(2481) ,
  \616(729) ,
  \1993(2659) ,
  \3971(1124) ,
  \3194(1617) ,
  \5679(2951) ,
  \2972(1515) ,
  \6917(335) ,
  \2436(1993) ,
  \1950(2047) ,
  \3549(1696) ,
  \2554(3085) ,
  \3755(412) ,
  \5148(3487) ,
  \1192(251) ,
  \6961(3457) ,
  \3235(2435) ,
  \6318(2632) ,
  \7479(890) ,
  \5940(2310) ,
  \4344(2188) ,
  \7617(2506) ,
  \268(3028) ,
  \2299(782) ,
  \318(3283) ,
  \6128(2611) ,
  \2764(2319) ,
  \3474(2998) ,
  \2504(2334) ,
  \5511(3503) ,
  \6935(3077) ,
  \4666(687) ,
  \5213(672) ,
  \5424(1437) ,
  \5009(3225) ,
  \2804(2327) ,
  \4076(3670) ,
  \6328(2642) ,
  \311(3349) ,
  \2754(2314) ,
  \6740(1265) ,
  \3026(2020) ,
  \763(723) ,
  \5314(1415) ,
  \6762(1689) ,
  \4966(1198) ,
  \2883(314) ,
  \7345(2154) ,
  \4889(378) ,
  \5173(3469) ,
  \6397(1167) ,
  \5631(3525) ,
  \3468(2898) ,
  \2002(2947) ,
  \4203(1923) ,
  \5368(2541) ,
  \6308(2647) ,
  \1230(2221) ,
  \2905(426) ,
  \1324(2461) ,
  \6106(3518) ,
  \1771(3137) ,
  \5597(3043) ,
  \4976(829) ,
  \3379(1480) ,
  \6594(1375) ,
  \4360(2699) ,
  \4143(744) ,
  \825(1279) ,
  \1138(2134) ,
  \5214(1449) ,
  \5904(1623) ,
  \6575(320) ,
  \1128(2132) ,
  \6340(2539) ,
  \7237(1701) ,
  \4132(707) ,
  \2152(660) ,
  \4381(2964) ,
  \1929(910) ,
  \6074(2793) ,
  \7432(1724) ,
  \5919(461) ,
  \2051(804) ,
  \5117(3113) ,
  \6670(2563) ,
  \5474(2948) ,
  \4570(1896) ,
  \2837(3682) ,
  \5980(2330) ,
  \6096(3460) ,
  \6407(903) ,
  \4042(2289) ,
  \4638(2723) ,
  \5540(2660) ,
  \3703(245) ,
  \1590(882) ,
  \3517(2120) ,
  \4647(580) ,
  \7033(3548) ,
  \3082(2179) ,
  \3267(3035) ,
  \7120(3608) ,
  \7110(3609) ,
  \2151(809) ,
  \6864(1352) ,
  \6134(3146) ,
  \3107(1305) ,
  \6861(321) ,
  \361(3324) ,
  \4710(762) ,
  \1074(1846) ,
  \4631(2866) ,
  \4442(290) ,
  \2629(1133) ,
  \6582(1688) ,
  \3571(2096) ,
  \971(3356) ,
  \1331(3188) ,
  \2052(658) ,
  \2341(1488) ,
  \2560(2800) ,
  \4544(2062) ,
  \5571(3523) ,
  \5315(965) ,
  \4968(3224) ,
  \6143(3383) ,
  \4094(584) ,
  \4417(217) ,
  \303(3271) ,
  \1991(3031) ,
  \1117(1193) ,
  \7157(3322) ,
  \1387(812) ,
  \2579(3011) ,
  \4783(3299) ,
  \6729(1301) ,
  \6543(937) ,
  \3801(824) ,
  \1025(1560) ,
  \5792(1243) ,
  \2812(2995) ,
  \6350(2514) ,
  \5889(343) ,
  \5639(3564) ,
  \4639(2973) ,
  \1329(3132) ,
  \5059(3507) ,
  \5579(3559) ,
  \4477(693) ,
  \3910(1775) ,
  \1710(2028) ,
  \7200(3699) ,
  \1133(2115) ,
  \4860(2358) ,
  \3131(2733) ,
  \1155(2201) ,
  \2537(2915) ,
  \4912(1451) ,
  \1249(1952) ,
  \5304(1407) ,
  \5250(1101) ,
  \2919(518) ,
  \3015(912) ,
  \701(541) ,
  \1291(2543) ,
  \3156(2706) ,
  \4081(3679) ,
  \6920(1276) ,
  \3652(668) ,
  \1323(2695) ,
  \4012(2255) ,
  \5433(364) ,
  \6033(350) ,
  \6815(2504) ,
  \2654(1795) ,
  \7487(881) ,
  \3660(608) ,
  \2924(610) ,
  \2833(317) ,
  \2285(616) ,
  \4949(2954) ,
  \4037(2298) ,
  \3164(2980) ,
  \2399(1792) ,
  \3891(1114) ,
  \6546(1057) ,
  \4027(2299) ,
  \1325(2848) ,
  \4154(996) ,
  \1257(1737) ,
  \6784(1396) ,
  \5729(3582) ,
  \615(529) ,
  \1247(1732) ,
  \6211(3491) ,
  \1545(1509) ,
  \6525(1207) ,
  \3522(1839) ,
  \5644(2064) ,
  \3540(2491) ,
  \6329(3641) ,
  \575(309) ,
  \7521(1652) ,
  \1412(818) ,
  \2861(3189) ,
  \6690(780) ,
  \581(421) ,
  \7079(3459) ,
  \2557(2928) ,
  \4618(2496) ,
  \2130(593) ,
  \1791(3701) ,
  \5258(1097) ,
  \641(841) ,
  \6677(1474) ,
  \4978(1926) ,
  \4508(1013) ,
  \6301(3490) ,
  \5218(1095) ,
  \5149(3528) ,
  \7271(1620) ,
  \2577(2920) ,
  \7188(3550) ,
  \5041(3360) ,
  \293(3285) ,
  \400(297) ,
  \6311(3537) ,
  \3856(1966) ,
  \7019(3456) ,
  \1366(528) ,
  \5848(2385) ,
  \2419(1796) ,
  \343(3258) ,
  \5318(816) ,
  \6835(3049) ,
  \6999(3140) ,
  \7515(1317) ,
  \4315(1877) ,
  \4880(566) ,
  \1555(1514) ,
  \7255(1364) ,
  \3232(2169) ,
  \2294(571) ,
  \1161(3229) ,
  \3595(2688) ,
  \3122(2158) ,
  \1609(1820) ,
  \2491(2608) ,
  \4235(1855) ,
  \2842(3681) ,
  \4375(2521) ,
  \4962(919) ,
  \1738(2067) ,
  \2545(2787) ,
  \3785(623) ,
  \6161(3520) ,
  \5664(2052) ,
  \6280(3096) ,
  \5654(2054) ,
  \1068(981) ,
  \6239(3633) ,
  \6565(1223) ,
  \6466(1019) ,
  \3793(796) ,
  \2335(1044) ,
  \7249(1024) ,
  \4669(490) ,
  \2777(2357) ,
  \4793(3203) ,
  \4140(745) ,
  \243(3032) ,
  \1779(3648) ,
  \3700(247) ,
  \5279(1458) ,
  \7581(1677) ,
  \4613(2728) ,
  \7575(1338) ,
  \6345(3054) ,
  \5269(1459) ,
  \5326(956) ,
  \4444(582) ,
  \4482(755) ,
  \1743(2070) ,
  \2979(886) ,
  \7235(1381) ,
  \4267(2143) ,
  \7348(2148) ,
  \3017(1524) ,
  \6025(349) ,
  \366(3381) ,
  \3102(2177) ,
  \3258(2546) ,
  \6279(3155) ,
  \3163(2861) ,
  \4552(1664) ,
  \7591(1671) ,
  \3673(821) ,
  \7585(1334) ,
  \6891(442) ,
  \6110(2318) ,
  \7169(3476) ,
  \2312(836) ,
  \6892(1603) ,
  \4539(1533) ,
  \3613(3108) ,
  \7436(2394) ,
  \3502(1573) ,
  \7602(2021) ,
  \1757(3594) ,
  \3028(2372) ,
  \5991(449) ,
  \7570(1308) ,
  \5812(966) ,
  \6876(1706) ,
  \5624(2076) ,
  \4577(2183) ,
  \2487(2312) ,
  \1920(1544) ,
  \6221(3536) ,
  \3140(2494) ,
  \6718(921) ,
  \6125(3087) ,
  \396(2941) ,
  \3031(2061) ,
  \3052(2192) ,
  \4052(2292) ,
  \6490(1299) ,
  \7132(2589) ,
  \7152(2584) ,
  \3739(233) ,
  \2157(792) ,
  \6151(3462) ,
  \7400(1398) ,
  \3062(2194) ,
  \827(1874) ,
  \3586(2704) ,
  \6189(3187) ,
  \7360(2216) ,
  \1869(1819) ,
  \1859(1818) ,
  \4529(1545) ,
  \6944(3139) ,
  \4668(701) ,
  \3169(597) ,
  \7068(2775) ,
  \7048(2777) ,
  \7364(1292) ,
  \2512(2354) ,
  \1166(3292) ,
  \3725(237) ,
  \5081(3640) ,
  \6382(1421) ,
  \7312(952) ,
  \6727(1611) ,
  \1173(3357) ,
  \5960(2614) ,
  \3380(1777) ,
  \2828(208) ,
  \5109(2959) ,
  \4841(2804) ,
  \6366(2963) ,
  \5039(3296) ,
  \3220(1761) ,
  \4314(1248) ,
  \378(3091) ,
  \1733(2057) ,
  \1723(2058) ,
  \6981(3568) ,
  \6352(2734) ,
  \5475(3038) ,
  \2954(1740) ,
  \4916(400) ,
  \5463(489) ,
  \5611(3348) ,
  \5614(2091) ,
  \4151(997) ,
  \2589(1981) ,
  \5369(2989) ,
  \5091(3639) ,
  \4352(2149) ,
  \7146(2911) ,
  \7061(3199) ,
  \7340(1931) ,
  \7229(1037) ,
  \5784(1436) ,
  \6787(1621) ,
  \7001(3193) ,
  \4540(1822) ,
  \4515(3099) ,
  \1985(2817) ,
  \3007(1575) ,
  \2304(728) ,
  \4059(3604) ,
  \7148(3078) ,
  \7304(948) ,
  \6418(947) ,
  \4674(684) ,
  \3525(1873) ,
  \1995(2819) ,
  \5551(3344) ,
  \5769(358) ,
  \351(3372) ,
  \606(403) ,
  \5927(464) ,
  \5254(1456) ,
  \251(3365) ,
  \6423(888) ,
  \6710(1213) ,
  \1953(2050) ,
  \2065(985) ,
  \6583(322) ,
  \7404(1042) ,
  \5687(3106) ,
  \5191(376) ,
  \2792(2355) ,
  \7211(1609) ,
  \6080(2343) ,
  \241(2837) ,
  \5494(3273) ,
  \5945(2609) ,
  \4518(3183) ,
  \5472(2822) ,
  \2179(977) ,
  \2962(867) ,
  \6077(3261) ,
  \3535(1885) ,
  \2918(736) ,
  \5621(3468) ,
  \3545(2155) ,
  \271(3354) ,
  \4572(2187) ,
  \4193(2493) ,
  \5561(3466) ,
  \3212(1367) ,
  \3222(1366) ,
  \1270(1583) ,
  \1948(2027) ,
  \4451(732) ,
  \826(1614) ,
  \2060(655) ,
  \1784(3617) ,
  \3242(3098) ,
  \3243(3171) ,
  \1178(261) ,
  \6415(907) ,
  \6086(3334) ,
  \5323(959) ,
  \2492(2313) ,
  \3979(1126) ,
  \1475(295) ,
  \3949(1122) ,
  \1762(3595) ,
  \3897(1475) ,
  \4439(209) ,
  \7239(1005) ,
  \7315(1427) ,
  \2279(739) ,
  \2417(1138) ,
  \987(3667) ,
  \4948(2680) ,
  \6666(2232) ,
  \6728(1278) ,
  \7012(3315) ,
  \6827(2700) ,
  \4768(2442) ,
  \4523(3246) ,
  \2734(1987) ,
  \4350(1861) ,
  \790(1208) ,
  \1395(814) ,
  \6121(1790) ,
  \6438(1233) ,
  \1957(2411) ,
  \2320(1025) ,
  \4728(2412) ,
  \7279(1595) ,
  \6090(2328) ,
  \2724(1722) ,
  \331(3364) ,
  \6141(3331) ,
  \5330(1235) ,
  \5897(344) ,
  \4224(1574) ,
  \6181(2987) ,
  \5069(3566) ,
  \3128(2509) ,
  \1445(2895) ,
  \3898(1772) ,
  \5844(2007) ,
  \5629(3505) ,
  \1964(3162) ,
  \5440(1240) ,
  \1500(296) ,
  \6991(2907) ,
  \6971(3513) ,
  \7224(1270) ,
  \3045(2651) ,
  \2801(2645) ,
  \5948(2311) ,
  \2791(2637) ,
  \6231(3593) ,
  \2982(1816) ,
  \6942(2764) ,
  \3655(550) ,
  \3911(1974) ,
  \2932(614) ,
  \4207(2198) ,
  \6888(1267) ,
  \6454(1354) ,
  \6287(3264) ,
  \719(850) ,
  \4138(689) ,
  \4234(1577) ,
  \623(533) ,
  \2771(2634) ,
  \4210(1712) ,
  \6100(2309) ,
  \2293(619) ,
  \2927(515) ,
  \4800(2598) ,
  \7204(3706) ,
  \6557(741) ,
  \2057(786) ,
  \618(632) ,
  \7059(3143) ,
  \5999(452) ,
  \7443(3061) ,
  \4791(3301) ,
  \6751(1705) ,
  \1450(2996) ,
  \4271(2857) ,
  \3116(1271) ,
  \6321(3592) ,
  \1004(3708) ,
  \5205(502) ,
  \2856(3709) ,
  \704(639) ,
  \961(3291) ,
  \2160(679) ,
  \349(3314) ,
  \4279(2982) ,
  \4064(3605) ,
  \1464(285) ,
  \5441(367) ,
  \5366(2217) ,
  \7477(1174) ,
  \7453(3062) ,
  \6622(1636) ,
  \6720(1189) ,
  \6605(440) ,
  \1990(2943) ,
  \4471(699) ,
  \4753(3158) ,
  \5569(3504) ,
  \4724(2048) ,
  \6916(1703) ,
  \2847(3624) ,
  \4980(2511) ,
  \3611(2718) ,
  \7566(1648) ,
  \3612(2970) ,
  \3101(1907) ,
  \939(2125) ,
  \1371(652) ,
  \7603(2196) ,
  \2992(1821) ,
  \4376(2714) ,
  \299(3341) ,
  \5399(466) ,
  \4623(2420) ,
  \1718(2046) ,
  \2866(3115) ,
  \1288(2219) ,
  \6259(3663) ,
  \4514(292) ,
  \3482(3075) ,
  \949(2129) ,
  \256(2991) ,
  \7301(949) ,
  \383(3089) ,
  \4101(734) ,
  \4955(3046) ,
  \6817(2744) ,
  \2998(896) ,
  \3472(2901) ,
  \994(3407) ,
  \727(848) ,
  \6829(2957) ,
  \3838(1004) ,
  \4868(2371) ,
  \4820(2281) ,
  \1943(2034) ,
  \1374(537) ,
  \4610(2502) ,
  \5871(450) ,
  \4317(2170) ,
  \2014(3274) ,
  \5542(3102) ,
  \2868(3308) ,
  \6426(1070) ,
  \4091(2899) ,
  \3663(493) ,
  \3029(2043) ,
  \6925(1115) ,
  \6132(2792) ,
  \4355(2207) ,
  \4927(508) ,
  \2547(3084) ,
  \5833(2393) ,
  \6434(954) ,
  \3457(2282) ,
  \5334(962) ,
  \5523(1158) ,
  \3872(1468) ,
  \906(1554) ,
  \1787(3678) ,
  \5337(1435) ,
  \1309(2545) ,
  \1996(2658) ,
  \5478(2388) ,
  \4422(215) ,
  \4998(3111) ,
  \957(1836) ,
  \3248(3293) ,
  \3987(1472) ,
  \4010(2552) ,
  \5799(485) ,
  \1986(2653) ,
  \1334(3190) ,
  \6542(1410) ,
  \5588(2672) ,
  \4677(477) ,
  \1777(3675) ,
  \2767(2341) ,
  \5608(2670) ,
  \1938(2006) ,
  \5977(1493) ,
  \2019(576) ,
  \4327(2186) ,
  \6447(1335) ,
  \3616(3184) ,
  \3202(1566) ,
  \1715(2391) ,
  \6249(3673) ,
  \6386(1069) ,
  \3988(1770) ,
  \2266(587) ,
  \5550(2401) ,
  \3873(1767) ,
  \7149(3198) ,
  \1007(773) ,
  \7384(1594) ,
  \5634(2045) ,
  \6678(2571) ,
  \4772(2105) ,
  \5514(3502) ,
  \4848(2631) ,
  \7393(1319) ,
  \2145(810) ,
  \5278(1103) ,
  \6695(983) ,
  \7309(1072) ,
  \944(2114) ,
  \2409(1989) ,
  \5719(3526) ,
  \6964(3454) ,
  \2507(2337) ,
  \1713(2030) ,
  \6844(2979) ,
  \3566(1940) ,
  \4707(763) ,
  \3601(2856) ,
  \5287(1413) ,
  \5159(3584) ,
  \4676(702) ,
  \1262(1234) ,
  \1685(1163) ,
  \3193(1731) ,
  \6840(2867) ,
  \4363(2465) ,
  \1299(2536) ,
  \7289(1628) ,
  \4831(3329) ,
  \6663(2567) ,
  \7335(1742) ,
  \3213(1735) ,
  \784(559) ,
  \6171(3573) ,
  \5661(3637) ,
  \4135(688) ,
  \2990(1579) ,
  \266(2956) ,
  \5064(2099) ,
  \4283(2694) ,
  \5651(3638) ,
  \4043(2301) ,
  \4593(1889) ,
  \4079(3669) ,
  \1307(2463) ,
  \6951(3313) ,
  \791(1559) ,
  \695(525) ,
  \1308(2752) ,
  \326(3294) ,
  \4281(2740) ,
  \3381(1976) ,
  \2617(1787) ,
  \3046(2813) ,
  \7391(1662) ,
  \7343(2191) ,
  \7325(1746) ,
  \6938(2562) ,
  \6219(3529) ,
  \4084(3627) ,
  \364(3326) ,
  \5756(1086) ,
  \5697(3276) ,
  \7424(1587) ,
  \6737(1360) ,
  \3550(2199) ,
  \2864(3245) ,
  \5084(2108) ,
  \1310(2887) ,
  \7074(2306) ,
  \7529(1661) ,
  \5051(3471) ,
  \4634(2863) ,
  \6277(3130) ,
  \5115(3052) ,
  \5900(1288) ,
  \4045(2288) ,
  \5094(2106) ,
  \3452(2295) ,
  \3679(776) ,
  \6687(943) ,
  \7307(1228) ,
  \261(2992) ,
  \4324(1284) ,
  \5238(1195) ,
  \950(2448) ,
  \4385(3060) ,
  \1186(254) ,
  \6487(1313) ,
  \5375(3070) ,
  \1253(2214) ,
  \1461(287) ,
  \2502(2317) ,
  \1790(2815) ,
  \4682(670) ,
  \6591(325) ,
  \4025(2277) ,
  \3215(1852) ,
  \3828(1035) ,
  \4035(2276) ,
  \2026(730) ,
  \4808(2583) ,
  \4913(497) ,
  \915(1029) ,
  \306(3270) ,
  \3563(2517) ,
  \2454(1996) ,
  \4997(1555) ,
  \320(3711) ,
  \6209(3464) ,
  \7540(1914) ,
  \2073(971) ,
  \4487(710) ,
  \1981(2655) ,
  \3192(931) ,
  \6405(1172) ,
  \4092(3705) ,
  \3583(2472) ,
  \4751(3284) ,
  \6993(3076) ,
  \1584(877) ,
  \5392(2885) ,
  \5129(3359) ,
  \5777(361) ,
  \7550(1910) ,
  \6309(3522) ,
  \3618(3244) ,
  \3173(717) ,
  \678(414) ,
  \6872(1377) ,
  \7408(1391) ,
  \1072(1214) ,
  \3483(2577) ,
  \3453(2578) ,
  \3195(1876) ,
  \7213(1306) ,
  \5037(3236) ,
  \4833(207) ,
  \6342(2750) ,
  \6168(2320) ,
  \6602(1359) ,
  \7219(1638) ,
  \7077(3428) ,
  \6148(2329) ,
  \5823(2657) ,
  \5263(1104) ,
  \2045(801) ,
  \933(2683) ,
  \1205(305) ,
  \417(3415) ,
  \7554(1011) ,
  \7456(2737) ,
  \4801(3250) ,
  \6502(1371) ,
  \5685(3042) ,
  \2146(661) ,
  \6164(3517) ,
  \4015(2257) ,
  \6869(323) ,
  \5968(2613) ,
  \626(636) ,
  \650(423) ,
  \7051(3007) ,
  \2955(1508) ,
  \2762(2326) ,
  \5038(2686) ,
  \5699(3347) ,
  \4137(746) ,
  \3442(2251) ,
  \4298(1867) ,
  \6064(2924) ,
  \885(832) ,
  \3649(511) ,
  \2597(1129) ,
  \6989(1769) ,
  \3398(1779) ,
  \3397(1482) ,
  \4040(2285) ,
  \5552(3272) ,
  \3899(1971) ,
  \5030(3051) ,
  \4704(764) ,
  \2817(3590) ,
  \6138(2342) ,
  \3635(408) ,
  \2354(1983) ,
  \7578(1312) ,
  \7518(1322) ,
  \4986(2742) ,
  \5992(1625) ,
  \3209(942) ,
  \1702(1999) ,
  \4849(2807) ,
  \5182(563) ,
  \4836(2745) ,
  \2970(872) ,
  \6613(441) ,
  \2298(716) ,
  \6299(3472) ,
  \2258(249) ,
  \3170(866) ,
  \5127(3295) ,
  \2921(512) ,
  \7020(2573) ,
  \1276(2145) ,
  \3265(3034) ,
  \709(545) ,
  \7446(2726) ,
  \7441(3039) ,
  \6075(3205) ,
  \7010(2575) ,
  \6055(1403) ,
  \5088(2447) ,
  \6772(1363) ,
  \6860(1665) ,
  \2198(974) ,
  \6291(3385) ,
  \6201(3386) ,
  \5098(2446) ,
  \6698(938) ,
  \5089(3621) ,
  \4713(3136) ,
  \7031(3530) ,
  \2288(555) ,
  \6753(1932) ,
  \4351(1917) ,
  \4942(1551) ,
  \792(1841) ,
  \2563(2756) ,
  \3598(2692) ,
  \5501(3441) ,
  \1868(1529) ,
  \1858(1528) ,
  \7263(1393) ,
  \7588(1336) ,
  \7091(3532) ,
  \386(3020) ,
  \5079(3622) ,
  \5068(2440) ,
  \3798(713) ,
  \3676(777) ,
  \1755(3580) ,
  \1217(1960) ,
  \5044(2136) ,
  \6482(1304) ,
  \1820(1157) ,
  \4020(2264) ,
  \2046(673) ,
  \7203(3657) ,
  \5800(1239) ,
  \2642(1794) ,
  \4178(1872) ,
  \2853(2784) ,
  \7470(915) ,
  \2899(590) ,
  \3240(3026) ,
  \1834(878) ,
  \1608(1530) ,
  \4188(1887) ,
  \1073(1565) ,
  \2137(738) ,
  \3271(3101) ,
  \4732(2051) ,
  \5600(3041) ,
  \1406(817) ,
  \1382(540) ,
  \6367(869) ,
  \5054(2121) ,
  \7610(2508) ,
  \3146(2871) ,
  \6049(1049) ,
  \6763(1918) ,
  \7040(2566) ,
  \7030(2554) ,
  \3342(1473) ,
  \3989(1969) ,
  \6041(342) ,
  \4660(581) ,
  \7558(1341) ,
  \3120(1871) ,
  \3788(552) ,
  \5953(2618) ,
  \4202(1362) ,
  \1171(3307) ,
  \6912(1374) ,
  \6154(3461) ,
  \1379(645) ,
  \4373(2519) ,
  \1736(2053) ,
  \6199(3337) ,
  \7282(1865) ,
  \5936(1949) ,
  \6832(1546) ,
  \6645(2762) ,
  \3123(2497) ,
  \4987(1549) ,
  \4671(488) ,
  \6533(1212) ,
  \2796(2529) ,
  \5988(1290) ,
  \3069(1934) ,
  \3343(1771) ,
  \6158(2308) ,
  \7458(2870) ,
  \6693(1222) ,
  \1365(644) ,
  \5712(2077) ,
  \6327(3612) ,
  \2526(2549) ,
  \3100(1886) ,
  \6899(443) ,
  \3874(1968) ,
  \4970(718) ,
  \3833(1016) ,
  \2822(3591) ,
  \5234(918) ,
  \5266(1091) ,
  \1477(394) ,
  \1141(2133) ,
  \5338(1241) ,
  \3327(1111) ,
  \5607(3221) ,
  \877(939) ,
  \3578(2437) ,
  \7448(2862) ,
  \4123(708) ,
  \7523(1323) ,
  \4905(380) ,
  \5709(3467) ,
  \5872(1626) ,
  \7167(3458) ,
  \6289(3335) ,
  \698(629) ,
  \7513(1325) ,
  \6807(1866) ,
  \1988(2818) ,
  \2301(783) ,
  \4621(2724) ,
  \3099(1268) ,
  \4134(747) ,
  \3435(2238) ,
  \5727(3563) ,
  \5448(1236) ,
  \5468(2665) ,
  \5581(911) ,
  \2587(1487) ,
  \5880(1596) ,
  \2559(2624) ,
  \4685(465) ,
  \2323(1038) ,
  \7351(2471) ,
  \4476(758) ,
  \4701(765) ,
  \7292(1881) ,
  \1519(374) ,
  \5078(2484) ,
  \3497(3319) ,
  \354(3375) ,
  \4595(2178) ,
  \6797(1862) ,
  \6735(1634) ,
  \3520(1564) ,
  \2840(3671) ,
  \2652(1139) ,
  \5049(3448) ,
  \5744(3698) ,
  \3110(2175) ,
  \2612(1131) ,
  \5074(2167) ,
  \1760(3581) ,
  \6210(2881) ,
  \4379(2854) ,
  \5067(3546) ,
  \2471(2209) ,
  \3312(1467) ,
  \4220(1619) ,
  \1447(3100) ,
  \1687(1813) ,
  \3241(2859) ,
  \2192(991) ,
  \2004(2666) ,
  \1332(3134) ,
  \5732(2063) ,
  \274(3353) ,
  \6430(1425) ,
  \2795(2368) ,
  \1741(2083) ,
  \4028(2579) ,
  \3719(239) ,
  \6485(1678) ,
  \4547(1532) ,
  \3665(600) ,
  \269(2896) ,
  \5649(3620) ,
  \1708(2378) ,
  \6024(1718) ,
  \6445(1670) ,
  \314(3350) ,
  \5905(347) ,
  \6826(2467) ,
  \5376(1961) ,
  \1788(2375) ,
  \5245(830) ,
  \2081(988) ,
  \5105(1569) ,
  \2418(1502) ,
  \3313(1766) ,
  \802(924) ,
  \7428(1404) ,
  \6319(3577) ,
  \995(3691) ,
  \572(427) ,
  \1174(3290) ,
  \6144(3333) ,
  \5638(2409) ,
  \7087(3497) ,
  \1018(606) ,
  \334(3362) ,
  \5659(3619) ,
  \4884(1105) ,
  \5048(2454) ,
  \6974(3512) ,
  \3114(1298) ,
  \4511(1012) ,
  \6805(1624) ,
  \5647(3597) ,
  \7022(3455) ,
  \4626(2404) ,
  \1017(831) ,
  \6390(1424) ,
  \5199(377) ,
  \1956(2087) ,
  \7257(1043) ,
  \6115(1494) ,
  \1966(2089) ,
  \5675(1541) ,
  \5536(2387) ,
  \3594(2719) ,
  \5785(362) ,
  \6900(1635) ,
  \5396(1084) ,
  \1507(418) ,
  \2859(3133) ,
  \6252(3614) ,
  \1151(2681) ,
  \5058(2451) ,
  \3020(1543) ,
  \6877(326) ,
  \3362(1117) ,
  \4761(3233) ,
  \2531(2547) ,
  \4624(2829) ,
  \5377(2988) ,
  \3440(2234) ,
  \2154(664) ,
  \6373(1147) ,
  \7399(1656) ,
  \4932(1547) ,
  \7135(1780) ,
  \5648(2422) ,
  \2053(805) ,
  \3568(2172) ,
  \294(3223) ,
  \4023(2582) ,
  \2871(315) ,
  \3090(1356) ,
  \3543(1869) ,
  \5702(2090) ,
  \6242(3635) ,
  \6779(1713) ,
  \6192(3154) ,
  \5628(2426) ,
  \6848(2851) ,
  \6007(453) ,
  \6559(944) ,
  \6462(1380) ,
  \4274(2852) ,
  \5618(2429) ,
  \3512(1616) ,
  \3484(2772) ,
  \3006(901) ,
  \3000(1534) ,
  \5668(2416) ,
  \5658(2417) ,
  \6510(1607) ,
  \5147(3508) ,
  \4230(2140) ,
  \7606(2197) ,
  \908(1192) ,
  \1272(1858) ,
  \2342(1784) ,
  \6431(914) ,
  \3399(1978) ,
  \3203(1847) ,
  \5221(505) ,
  \895(1850) ,
  \3018(1814) ,
  \5190(562) ,
  \1789(2652) ,
  \6819(2152) ,
  \5222(1450) ,
  \1606(892) ,
  \7333(1419) ,
  \937(2162) ,
  \6229(3579) ,
  \3485(2909) ,
  \3654(682) ,
  \4243(1747) ,
  \5449(359) ,
  \5407(470) ,
  \3475(3074) ,
  \2287(620) ,
  \5752(1440) ,
  \2465(1144) ,
  \7323(1423) ,
  \6674(2245) ,
  \4721(3217) ,
  \4131(748) ,
  \4780(2168) ,
  \3238(2684) ,
  \5262(1452) ,
  \4008(2242) ,
  \5868(1291) ,
  \280(391) ,
  \6621(444) ,
  \765(774) ,
  \1126(2165) ,
  \5943(2791) ,
  \620(633) ,
  \4958(3048) ,
  \4266(2458) ,
  \4479(694) ,
  \1782(3616) ,
  \1946(2033) ,
  \4353(1720) ,
  \4242(1580) ,
  \985(3653) ,
  \7101(3589) ,
  \5856(2398) ,
  \5807(486) ,
  \5152(2098) ,
  \7242(1018) ,
  \6056(1948) ,
  \4776(2445) ,
  \4297(1293) ,
  \7412(1039) ,
  \7147(3142) ,
  \2942(859) ,
  \6297(3436) ,
  \6406(1230) ,
  \617(530) ,
  \4048(2594) ,
  \5717(3506) ,
  \6945(3248) ,
  \5020(2844) ,
  \4736(2415) ,
  \2926(611) ,
  \5237(720) ,
  \3175(1558) ,
  \703(542) ,
  \4847(2932) ,
  \398(3713) ,
  \5281(1058) ,
  \1989(2654) ,
  \5956(2316) ,
  \1961(2072) ,
  \3491(3249) ,
  \2054(676) ,
  \1822(1811) ,
  \5331(1080) ,
  \3662(601) ,
  \6336(3704) ,
  \6268(2808) ,
  \3233(2119) ,
  \3792(714) ,
  \4698(766) ,
  \7156(2774) ,
  \7136(2776) ,
  \7212(1277) ,
  \1368(520) ,
  \893(1220) ,
  \3292(1107) ,
  \5921(351) ,
  \4356(2466) ,
  \7372(1263) ,
  \803(1211) ,
  \7232(1033) ,
  \3657(504) ,
  \4601(2406) ,
  \3619(3181) ,
  \4799(3259) ,
  \247(3310) ,
  \3670(778) ,
  \2032(592) ,
  \6288(2805) ,
  \6506(1272) ,
  \3604(2853) ,
  \1225(1755) ,
  \381(3092) ,
  \6135(3260) ,
  \5879(451) ,
  \4828(2293) ,
  \927(2112) ,
  \6630(1631) ,
  \6954(3316) ,
  \5018(2713) ,
  \2732(1496) ,
  \947(2113) ,
  \1458(289) ,
  \7179(3533) ,
  \7500(873) ,
  \2407(1499) ,
  \1050(930) ,
  \894(1570) ,
  \5617(3395) ,
  \7611(2193) ,
  \371(2754) ,
  \3221(557) ,
  \3787(624) ,
  \4809(3253) ,
  \1215(1758) ,
  \3185(1563) ,
  \4046(2303) ,
  \953(1197) ,
  \1524(301) ,
  \4602(2041) ,
  \1856(2037) ,
  \3782(553) ,
  \4286(2693) ,
  \804(1562) ,
  \5242(917) ,
  \2167(990) ,
  \4335(1653) ,
  \7485(1166) ,
  \6087(3435) ,
  \5696(2669) ,
  \4386(2698) ,
  \3244(1962) ,
  \3795(797) ,
  \3152(3305) ,
  \6809(2190) ,
  \5311(1060) ,
  \7574(1640) ,
  \3344(1970) ,
  \4640(409) ,
  \3596(2450) ,
  \6375(874) ,
  \7108(2592) ,
  \6394(1073) ,
  \4484(754) ,
  \6261(1944) ,
  \7121(3643) ,
  \3016(1745) ,
  \367(3328) ,
  \4637(2864) ,
  \5428(963) ,
  \1313(2886) ,
  \5526(2662) ,
  \5000(3169) ,
  \2001(2825) ,
  \2845(3626) ,
  \4361(2470) ,
  \1373(648) ,
  \7111(3644) ,
  \5619(3443) ,
  \1848(1160) ,
  \4470(761) ,
  \329(3298) ,
  \2867(3239) ,
  \5139(3470) ,
  \7098(2581) ,
  \4299(1912) ,
  \6721(1274) ,
  \4888(1460) ,
  \1706(2015) ,
  \5912(1717) ,
  \1296(2212) ,
  \3544(1922) ,
  \4402(223) ,
  \4364(2720) ,
  \5118(3050) ,
  \4499(1001) ,
  \4038(2271) ,
  \1567(876) ,
  \4521(3186) ,
  \992(3404) ,
  \4219(1942) ,
  \6646(2556) ,
  \5841(2392) ,
  \4129(691) ,
  \4924(1099) ,
  \692(626) ,
  \2965(1805) ,
  \2556(2801) ,
  \5532(2946) ,
  \5157(3565) ,
  \3127(2725) ,
  \5975(1498) ,
  \7593(1905) ,
  \4524(3265) ,
  \6701(1281) ,
  \3027(2040) ,
  \5355(1438) ,
  \5637(3542) ,
  \5751(467) ,
  \4382(2972) ,
  \6781(1286) ,
  \254(2888) ,
  \2255(252) ,
  \5932(1726) ,
  \309(3275) ,
  \5347(1750) ,
  \342(3330) ,
  \6626(1297) ,
  \3686(838) ,
  \4013(2236) ,
  \5722(2044) ,
  \1628(1176) ,
  \967(3355) ,
  \6795(1591) ,
  \5559(3440) ,
  \2741(2210) ,
  \2159(793) ,
  \5393(352) ,
  \7507(1002) ,
  \5808(1237) ,
  \3956(1778) ,
  \7361(1343) ,
  \3995(1486) ,
  \5357(1753) ,
  \4928(1454) ,
  \6290(3262) ,
  \6745(1376) ,
  \7165(3427) ,
  \7216(1300) ,
  \6518(558) ,
  \6455(1337) ,
  \6122(2923) ,
  \5226(1100) ,
  \5913(348) ,
  \664(574) ,
  \6550(1412) ,
  \4251(2476) ,
  \5852(2026) ,
  \3955(1481) ,
  \6599(327) ,
  \1553(870) ,
  \6686(2570) ,
  \5676(2671) ,
  \6332(3697) ,
  \4856(2639) ,
  \6493(1647) ,
  \6478(1604) ,
  \302(3342) ,
  \1327(3071) ,
  \5688(3040) ,
  \4169(1009) ,
  \1287(2544) ,
  \7029(3514) ,
  \2505(2336) ,
  \4254(2708) ,
  \1280(1751) ,
  \942(2110) ,
  \574(308) ,
  \3314(1967) ,
  \2850(3083) ,
  \5572(3501) ,
  \2241(257) ,
  \757(856) ,
  \3996(1782) ,
  \4282(2983) ,
  \6355(3119) ,
  \5125(3234) ,
  \4695(767) ,
  \352(3318) ,
  \2653(1501) ,
  \3445(2254) ,
  \1883(1177) ,
  \6541(1282) ,
  \7089(3515) ,
  \5793(365) ,
  \1221(2222) ,
  \6885(329) ,
  \7002(3138) ,
  \3201(1733) ,
  \6066(3015) ,
  \3108(1883) ,
  \990(3685) ,
  \1535(302) ,
  \4041(2300) ,
  \2295(781) ,
  \5077(3601) ,
  \7401(1318) ,
  \805(1844) ,
  \7557(1651) ,
  \4334(1939) ,
  \6852(2965) ,
  \5764(1075) ,
  \6341(2538) ,
  \4561(1897) ,
  \4571(1898) ,
  \1775(3666) ,
  \6365(3129) ,
  \4457(583) ,
  \2765(2324) ,
  \2755(2325) ,
  \7353(1954) ,
  \1541(275) ,
  \3713(241) ,
  \2860(3068) ,
  \3466(2558) ,
  \5908(1394) ,
  \1711(2012) ,
  \7238(1708) ,
  \4077(3659) ,
  \4180(2159) ,
  \2352(1489) ,
  \1152(1369) ,
  \5246(1194) ,
  \5657(3651) ,
  \5667(3650) ,
  \1693(1184) ,
  \6996(2561) ,
  \5345(1429) ,
  \4609(2729) ,
  \5485(3213) ,
  \6015(458) ,
  \6765(1365) ,
  \5504(3438) ,
  \6495(1311) ,
  \4354(1943) ,
  \7099(3572) ,
  \1238(1727) ,
  \2838(3672) ,
  \2799(2531) ,
  \1312(2542) ,
  \1653(1179) ,
  \2062(657) ,
  \6868(1690) ,
  \5142(2123) ,
  \389(3021) ,
  \3478(3001) ,
  \7327(1064) ,
  \5415(472) ,
  \913(1027) ,
  \3460(2284) ,
  \5372(1759) ,
  \1803(1152) ,
  \5888(1593) ,
  \5985(336) ,
  \579(840) ,
  \2162(659) ,
  \4936(1834) ,
  \6706(933) ,
  \6413(1175) ,
  \5388(2751) ,
  \3930(1479) ,
  \3508(2138) ,
  \5530(2821) ,
  \4816(2586) ,
  \3211(827) ,
  \4082(3687) ,
  \4126(692) ,
  \2675(1798) ,
  \2950(865) ,
  \2500(2322) ,
  \6267(2208) ,
  \7537(1684) ,
  \332(3304) ,
  \821(929) ,
  \322(3302) ,
  \7317(1068) ,
  \6298(2880) ,
  \1780(3674) ,
  \4312(1256) ,
  \1739(2082) ,
  \7420(1249) ,
  \5132(2135) ,
  \7547(1680) ,
  \1108(1196) ,
  \3227(1925) ,
  \4938(2202) ,
  \7039(3567) ,
  \3450(2274) ,
  \3531(2480) ,
  \3459(3196) ,
  \4946(1837) ,
  \6114(2615) ,
  \7595(1801) ,
  \4316(1899) ,
  \5457(368) ,
  \7139(3006) ,
  \2929(516) ,
  \1086(935) ,
  \3415(1484) ,
  \777(370) ,
  \3816(1021) ,
  \1383(815) ,
  \5400(1439) ,
  \3931(1776) ,
  \3093(2156) ,
  \4300(2153) ,
  \706(640) ,
  \7128(2587) ,
  \7088(2595) ,
  \625(534) ,
  \5831(2656) ,
  \2059(787) ,
  \2290(569) ,
  \1343(575) ,
  \7118(2588) ,
  \5590(2833) ,
  \1792(3707) ,
  \3768(595) ,
  \2518(2353) ,
  \6717(916) ,
  \4952(1204) ,
  \5156(2439) ,
  \5174(3700) ,
  \1248(1730) ,
  \5533(3037) ,
  \5295(1409) ,
  \6398(1428) ,
  \2779(2527) ,
  \6703(927) ,
  \1914(905) ,
  \5270(1446) ,
  \2548(2922) ,
  \5383(3066) ,
  \1311(2753) ,
  \6060(2799) ,
  \6908(1630) ,
  \4629(2730) ,
  \2715(1145) ,
  \7078(2600) ,
  \1357(589) ,
  \5815(491) ,
  \2372(1986) ,
  \6222(3521) ,
  \4876(401) ,
  \6907(445) ,
  \2920(615) ,
  \6880(1361) ,
  \1304(2147) ,
  \6226(2347) ,
  \4473(697) ,
  \3416(1781) ,
  \4784(2485) ,
  \3591(2490) ,
  \3259(2874) ,
  \6743(1693) ,
  \2529(2548) ,
  \3350(2261) ,
  \3651(509) ,
  \2862(3185) ,
  \4535(2093) ,
  \6551(599) ,
  \7416(1386) ,
  \5003(920) ,
  \3513(1848) ,
  \4796(2304) ,
  \2806(2755) ,
  \384(3016) ,
  \6307(3509) ,
  \1686(1522) ,
  \4107(585) ,
  \7246(1355) ,
  \3117(1930) ,
  \1134(2131) ,
  \357(3376) ,
  \5887(454) ,
  \5976(2623) ,
  \6097(3498) ,
  \4226(1854) ,
  \3790(551) ,
  \7522(1660) ,
  \4692(768) ,
  \6264(2640) ,
  \2536(2789) ,
  \6383(880) ,
  \7526(1320) ,
  \7175(3496) ,
  \3438(2239) ,
  \3129(2516) ,
  \764(603) ,
  \6351(2505) ,
  \4087(3695) ,
  \2843(3689) ,
  \4769(3242) ,
  \4056(3005) ,
  \4464(733) ,
  \3068(1353) ,
  \244(3033) ,
  \2788(2356) ,
  \4879(495) ,
  \7497(868) ,
  \5359(1957) ,
  \2757(2602) ,
  \3008(1539) ,
  \2635(1135) ,
  \250(3417) ,
  \1805(1806) ,
  \4921(381) ,
  \2514(2523) ,
  \2881(3339) ,
  \3781(621) ,
  \7392(1618) ,
  \2524(2525) ,
  \387(2931) ,
  \5322(955) ,
  \3821(1034) ,
  \2989(889) ,
  \6284(2635) ,
  \5436(961) ,
  \7592(1674) ,
  \2808(2917) ,
  \7016(2249) ,
  \7049(2781) ,
  \4759(3211) ,
  \629(844) ,
  \4553(1663) ,
  \2778(2366) ,
  \4729(3218) ,
  \1376(546) ,
  \4558(2189) ,
  \1744(2085) ,
  \7189(3588) ,
  \5040(3232) ,
  \2798(2367) ,
  \1795(1804) ,
  \5108(2843) ,
  \5929(1048) ,
  \3149(3182) ,
  \4225(1225) ,
  \5339(1074) ,
  \7236(1372) ,
  \4947(2836) ,
  \6562(1059) ,
  \6638(1612) ,
  \4679(476) ,
  \3032(2079) ,
  \1055(1875) ,
  \4306(1864) ,
  \317(3351) ,
  \7036(2237) ,
  \2848(3693) ,
  \5961(2617) ,
  \3621(3240) ,
  \7080(3433) ,
  \5028(2842) ,
  \7026(2225) ,
  \2761(2783) ,
  \3141(2492) ,
  \4614(2495) ,
  \1235(1958) ,
  \5627(3485) ,
  \6522(1063) ,
  \697(526) ,
  \4678(703) ,
  \5349(1083) ,
  \2700(1799) ,
  \6337(2961) ,
  \611(573) ,
  \7551(1316) ,
  \1121(1552) ,
  \2794(2528) ,
  \7162(2305) ,
  \5207(549) ,
  \2813(2930) ,
  \1969(2088) ,
  \7247(1691) ,
  \3957(1977) ,
  \6653(2761) ,
  \6812(2204) ,
  \2807(2648) ,
  \4128(749) ,
  \5167(3446) ,
  \6084(2626) ,
  \4740(2066) ,
  \5289(1054) ,
  \4627(2827) ,
  \2513(2362) ,
  \2523(2363) ,
  \3425(1125) ,
  \6271(3064) ,
  \3335(1113) ,
  \3136(2475) ,
  \6212(3473) ,
  \2435(1797) ,
  \2007(3161) ,
  \7437(2373) ,
  \1655(1827) ,
  \2153(791) ,
  \7495(1523) ,
  \2453(1800) ,
  \5824(2380) ,
  \6094(2620) ,
  \1734(2068) ,
  \5137(3447) ,
  \1724(2069) ,
  \1695(1829) ,
  \4150(704) ,
  \2797(2644) ,
  \2670(1141) ,
  \6104(2605) ,
  \5155(3547) ,
  \3148(3059) ,
  \6928(2770) ,
  \3183(926) ,
  \4114(735) ,
  \5473(2826) ,
  \4670(686) ,
  \2448(1142) ,
  \4396(225) ,
  \5126(2685) ,
  \7109(3632) ,
  \7119(3631) ,
  \3477(2766) ,
  \6816(2515) ,
  \3200(982) ,
  \1939(2017) ,
  \3997(1980) ,
  \3775(740) ,
  \4531(1830) ,
  \4989(2679) ,
  \751(857) ,
  \5695(3219) ,
  \4387(2850) ,
  \6052(1725) ,
  \6032(1714) ,
  \4263(2142) ,
  \3467(2760) ,
  \7425(1047) ,
  \2300(726) ,
  \6000(1597) ,
  \2493(2321) ,
  \5097(3654) ,
  \6179(1946) ,
  \1314(2749) ,
  \5876(1259) ,
  \3667(779) ,
  \5087(3655) ,
  \4554(1900) ,
  \1271(1584) ,
  \4684(669) ,
  \7300(946) ,
  \5384(1953) ,
  \1261(1582) ,
  \6023(459) ,
  \5471(1162) ,
  \4369(2486) ,
  \4277(2876) ,
  \2550(3013) ,
  \1785(3618) ,
  \6983(1470) ,
  \2175(975) ,
  \3176(1840) ,
  \5726(2408) ,
  \1954(2060) ,
  \7614(2181) ,
  \5380(1736) ,
  \3070(1675) ,
  \7541(1342) ,
  \5106(2712) ,
  \6107(3555) ,
  \6186(2811) ,
  \2793(2364) ,
  \6554(396) ,
  \3186(1845) ,
  \3603(2969) ,
  \988(3652) ,
  \4857(2810) ,
  \6133(3204) ,
  \7054(2779) ,
  \1240(1950) ,
  \1793(1149) ,
  \4606(2503) ,
  \6442(1006) ,
  \4563(2184) ,
  \4887(500) ,
  \6828(2701) ,
  \2213(268) ,
  \2809(2893) ,
  \4630(2977) ,
  \4121(228) ,
  \1885(1825) ,
  \5404(1087) ,
  \7265(1285) ,
  \4525(862) ,
  \5993(339) ,
  \5737(3636) ,
  \6453(1673) ,
  \7531(1346) ,
  \4259(2487) ,
  \1821(1518) ,
  \3582(2705) ,
  \1949(2036) ,
  \5935(1402) ,
  \6755(1328) ,
  \6932(2905) ,
  \1153(1700) ,
  \6118(2798) ,
  \6799(1289) ,
  \5423(478) ,
  \6629(446) ,
  \4489(709) ,
  \4990(2953) ,
  \7205(1273) ,
  \6714(775) ,
  \1897(900) ,
  \2980(1748) ,
  \1488(279) ,
  \628(637) ,
  \2047(802) ,
  \5284(1051) ,
  \7478(1181) ,
  \7369(1344) ,
  \7367(1681) ,
  \7006(2259) ,
  \7409(1321) ,
  \3932(1975) ,
  \5047(3410) ,
  \5863(1520) ,
  \3536(2174) ,
  \1207(307) ,
  \2147(807) ,
  \6893(330) ,
  \4807(3321) ,
  \3410(1123) ,
  \1391(813) ,
  \6642(2227) ,
  \6752(1702) ,
  \5321(1244) ,
  \3602(2711) ,
  \1210(298) ,
  \5162(2166) ,
  \2048(653) ,
  \5146(2452) ,
  \5136(2453) ,
  \1630(1824) ,
  \5735(3596) ,
  \4057(3586) ,
  \6236(2360) ,
  \4719(3192) ,
  \5996(1260) ,
  \6202(3336) ,
  \5669(1182) ,
  \3629(578) ,
  \6789(1253) ,
  \5057(3489) ,
  \6965(3492) ,
  \4211(1716) ,
  \5229(510) ,
  \6317(3558) ,
  \1158(1927) ,
  \886(604) ,
  \715(851) ,
  \4959(3170) ,
  \6216(2369) ,
  \6639(2560) ,
  \5895(456) ,
  \2923(513) ,
  \1316(2882) ,
  \4481(696) ,
  \1023(1205) ,
  \1647(899) ,
  \868(934) ,
  \7407(1654) ,
  \6246(2351) ,
  \7601(1997) ,
  \5230(1455) ,
  \6570(1329) ,
  \5280(1457) ,
  \1381(651) ,
  \6915(437) ,
  \6256(2350) ,
  \257(2860) ,
  \2470(1945) ,
  \6145(3434) ,
  \5760(1441) ,
  \6682(2244) ,
  \1370(521) ,
  \3607(2875) ,
  \5610(3216) ,
  \7177(3516) ,
  \3458(2294) ,
  \700(630) ,
  \3800(700) ,
  \6124(3014) ,
  \2186(989) ,
  \2655(1991) ,
  \1440(3030) ,
  \4284(2456) ,
  \7380(1257) ,
  \4198(2157) ,
  \2039(737) ,
  \4157(1010) ,
  \5864(2397) ,
  \5070(3545) ,
  \1709(2016) ,
  \5444(957) ,
  \6904(1296) ,
  \5951(2790) ,
  \5820(2002) ,
  \3648(665) ,
  \2148(678) ,
  \5839(2664) ,
  \3147(3116) ,
  \4727(3278) ,
  \4929(564) ,
  \2238(259) ,
  \5589(2677) ,
  \4996(3045) ,
  \5385(2962) ,
  \5660(3598) ,
  \5650(3599) ,
  \3184(1729) ,
  \3417(1979) ,
  \6748(1373) ,
  \3843(1463) ,
  \2111(987) ,
  \6818(2732) ,
  \3025(2005) ,
  \1749(2022) ,
  \637(842) ,
  \4184(2479) ,
  \1499(273) ,
  \7431(1401) ,
  \5401(355) ,
  \5011(941) ,
  \7067(3256) ,
  \2600(1984) ,
  \5736(2421) ,
  \5408(1442) ,
  \6020(1395) ,
  \3464(3200) ,
  \6578(1350) ,
  \6470(1357) ,
  \723(849) ,
  \2522(2550) ,
  \2578(3082) ,
  \962(2839) ,
  \5706(2428) ,
  \3762(586) ,
  \3579(2473) ,
  \7260(1040) ,
  \5166(2483) ,
  \7090(3494) ,
  \5716(2427) ,
  \594(572) ,
  \372(2890) ,
  \3174(1738) ,
  \1880(895) ,
  \1850(1812) ,
  \4581(2500) ,
  \3557(1935) ,
  \2818(3575) ,
  \4308(2151) ,
  \4855(2935) ,
  \4788(2118) ,
  \3844(1762) ,
  \6607(328) ,
  \3021(1831) ,
  \4744(2423) ,
  \851(1217) ,
  \4516(3024) ,
  \1233(1754) ,
  \305(3343) ,
  \4216(2206) ,
  \5801(366) ,
  \5896(1588) ,
  \5964(2315) ,
  \4673(483) ,
  \4272(2710) ,
  \4062(3587) ,
  \6176(2809) ,
  \1714(2031) ,
  \7336(1739) ,
  \6193(3263) ,
  \6196(2806) ,
  \6414(1229) ,
  \6711(772) ,
  \2308(835) ,
  \2303(784) ,
  \2472(2532) ,
  \4262(2715) ,
  \4817(3254) ,
  \5215(379) ,
  \5598(2831) ,
  \7326(1743) ,
  \6634(1275) ,
  \6391(891) ,
  \355(3317) ,
  \2259(413) ,
  \6486(1637) ,
  \5759(469) ,
  \852(1568) ,
  \3001(1823) ,
  \6048(1589) ,
  \5128(3231) ,
  \3034(2403) ,
  \7438(2650) ,
  \7505(1511) ,
  \1596(1168) ,
  \7583(1891) ,
  \7582(1646) ,
  \2784(2802) ,
  \3463(2296) ,
  \6758(1351) ,
  \5707(3442) ,
  \7168(3432) ,
  \1284(2220) ,
  \7176(2596) ,
  \7166(2599) ,
  \2161(794) ,
  \4085(3629) ,
  \4478(757) ,
  \5483(3160) ,
  \5920(1715) ,
  \5678(2832) ,
  \7208(978) ,
  \6232(3578) ,
  \5181(494) ,
  \3118(1644) ,
  \5705(3394) ,
  \4748(2075) ,
  \4011(2243) ,
  \4051(2247) ,
  \4343(1658) ,
  \7356(1955) ,
  \6654(2557) ,
  \1315(2534) ,
  \2973(1808) ,
  \3155(3366) ,
  \5725(3543) ,
  \4026(2287) ,
  \945(2128) ,
  \1471(283) ,
  \1244(2211) ,
  \262(2993) ,
  \691(523) ,
  \4036(2286) ,
  \6822(2150) ,
  \7308(1227) ,
  \6719(1202) ,
  \7196(2591) ,
  \2249(255) ,
  \2210(270) ,
  \5816(1245) ,
  \1778(3665) ,
  \2763(2338) ,
  \6031(462) ,
  \2588(1783) ,
  \4594(1890) ,
  \4584(1893) ,
  \2933(861) ,
  \4197(1921) ,
  \7493(1155) ,
  \7503(1146) ,
  \3121(1894) ,
  \1038(1843) ,
  \4072(3202) ,
  \4865(2877) ,
  \6063(1495) ,
  \374(3152) ,
  \6709(1206) ,
  \4307(1915) ,
  \6943(3194) ,
  \912(1550) ,
  \4519(3124) ,
  \6573(432) ,
  \5969(1137) ,
  \1751(2828) ,
  \2892(416) ,
  \297(3266) ,
  \3575(2095) ,
  \5594(2675) ,
  \4767(3297) ,
  \2503(2323) ,
  \7598(1809) ,
  \916(1030) ,
  \6155(3499) ,
  \2981(1526) ,
  \1944(2009) ,
  \1145(3179) ,
  \3554(2510) ,
  \4864(2641) ,
  \3277(2891) ,
  \335(3300) ,
  \6335(3656) ,
  \267(3027) ,
  \5515(3539) ,
  \6773(1388) ,
  \2305(826) ,
  \6764(1901) ,
  \4689(769) ,
  \1571(1156) ,
  \2370(1492) ,
  \3091(1870) ,
  \1006(602) ,
  \1941(2379) ,
  \4483(712) ,
  \4305(1262) ,
  \3231(2109) ,
  \4895(503) ,
  \2156(662) ,
  \4285(2845) ,
  \6065(2927) ,
  \4967(3288) ,
  \1127(2116) ,
  \6637(447) ,
  \5288(1406) ,
  \2823(3576) ,
  \6095(3478) ,
  \2641(1500) ,
  \1137(2117) ,
  \5194(1106) ,
  \7447(2735) ,
  \7457(2736) ,
  \3885(1112) ,
  \2155(800) ,
  \3022(1998) ,
  \6685(1768) ,
  \6606(1692) ,
  \5860(2025) ,
  \4016(2258) ,
  \5772(1078) ,
  \1295(2537) ,
  \4348(1385) ,
  \1053(1280) ,
  \4549(1815) ,
  \6549(1215) ,
  \5431(481) ,
  \6955(3423) ,
  \6180(2936) ,
  \3443(2253) ,
  \242(2955) ,
  \1116(1031) ,
  \2991(1531) ,
  \6183(3131) ,
  \2909(417) ,
  \6190(2939) ,
  \853(1849) ,
  \3707(243) ,
  \5367(2540) ,
  \1303(2462) ,
  \5303(1417) ,
  \2003(2399) ,
  \6016(1622) ,
  \2865(3180) ,
  \737(854) ,
  \7359(2215) ,
  \5313(1416) ,
  \4407(221) ,
  \5488(2039) ,
  \[100] ,
  \4342(1936) ,
  \[101] ,
  \[102] ,
  \1256(1728) ,
  \6923(448) ,
  \[103] ,
  \[104] ,
  \4617(2722) ,
  \6346(2884) ,
  \[105] ,
  \[106] ,
  \6200(2933) ,
  \5562(3439) ,
  \5916(1390) ,
  \2931(517) ,
  \[107] ,
  \5231(561) ,
  \1019(923) ,
  \4576(1650) ,
  \1754(2950) ,
  \1482(281) ,
  \2495(2601) ,
  \2549(2795) ,
  \2061(788) ,
  \1267(2144) ,
  \5495(3392) ,
  \6421(1180) ,
  \5008(3289) ,
  \6463(1309) ,
  \622(634) ,
  \6761(1666) ,
  \1002(2682) ,
  \7565(1679) ,
  \925(2103) ,
  \6754(1933) ,
  \6105(3535) ,
  \7178(3495) ,
  \5239(719) ,
  \2329(1041) ,
  \2558(3017) ,
  \6028(1389) ,
  \1849(1521) ,
  \5865(337) ,
  \2928(612) ,
  \2527(2524) ,
  \5498(2023) ,
  \4333(1397) ,
  \3656(667) ,
  \6008(1592) ,
  \619(531) ,
  \6671(1116) ,
  \7280(1586) ,
  \3486(3004) ,
  \5640(3541) ,
  \7510(1003) ,
  \2420(1992) ,
  \4289(1880) ,
  \2289(617) ,
  \6694(945) ,
  \2056(674) ,
  \2232(262) ,
  \4032(2773) ,
  \4840(2879) ,
  \1279(1585) ,
  \705(543) ,
  \645(847) ,
  \7462(2981) ,
  \1160(3173) ,
  \1629(1535) ,
  \1140(3176) ,
  \6172(2616) ,
  \6356(2869) ,
  \312(3279) ,
  \3363(1477) ,
  \6618(1303) ,
  \1669(904) ,
  \3076(1379) ,
  \4147(705) ,
  \7559(1340) ,
  \7186(2580) ,
  \6044(1251) ,
  \6004(1254) ,
  \4172(1008) ,
  \7013(3422) ,
  \6314(2346) ,
  \4212(1937) ,
  \7097(3552) ,
  \6381(1151) ,
  \1258(1951) ,
  \7320(1071) ,
  \2857(293) ,
  \5391(3055) ,
  \4374(2518) ,
  \7032(3511) ,
  \2400(1988) ,
  \3293(1465) ,
  \2733(1791) ,
  \1367(650) ,
  \6142(2625) ,
  \4686(770) ,
  \7057(3081) ,
  \7452(2975) ,
  \3794(724) ,
  \2406(2344) ,
  \2297(790) ,
  \6808(1879) ,
  \5024(2689) ,
  \272(3287) ,
  \1756(3561) ,
  \4892(1090) ,
  \671(424) ,
  \3659(499) ,
  \3789(625) ,
  \5348(1749) ,
  \5090(3602) ,
  \2408(1793) ,
  \1737(2056) ,
  \6152(2621) ,
  \5329(1238) ,
  \3797(798) ,
  \3617(3126) ,
  \3294(1764) ,
  \3597(2841) ,
  \6771(1697) ,
  \4777(3235) ,
  \5080(3603) ,
  \3784(567) ,
  \1375(643) ,
  \3139(2474) ,
  \3845(1963) ,
  \7530(1657) ,
  \5817(2384) ,
  \5247(1098) ,
  \4937(1929) ,
  \2740(1947) ,
  \3364(1774) ,
  \3599(2436) ,
  \1901(1178) ,
  \5984(2622) ,
  \4486(753) ,
  \1884(1536) ,
  \4093(3710) ,
  \2742(2533) ,
  \1598(1817) ,
  \4080(3658) ,
  \4939(2512) ,
  \5223(382) ,
  \345(3370) ,
  \4125(750) ,
  \1512(300) ,
  \4472(760) ,
  \2091(969) ,
  \2693(1143) ,
  \4681(471) ,
  \5601(3166) ,
  \5034(2444) ,
  \5541(3159) ,
  \5768(1430) ,
  \3521(1557) ,
  \7514(1326) ,
  \2543(3009) ,
  \1146(2431) ,
  \2316(837) ,
  \4244(1856) ,
  \4548(1525) ,
  \7264(1387) ,
  \6474(1269) ,
  \6798(1863) ,
  \694(627) ,
  \5019(2691) ,
  \392(3022) ,
  \2876(389) ,
  \3481(3000) ,
  \6206(2747) ,
  \7187(3571) ,
  \5158(3544) ,
  \1866(893) ,
  \920(2100) ,
  \265(2835) ,
  \1694(1542) ,
  \1115(371) ,
  \1317(2748) ,
  \3605(2703) ,
  \5698(3215) ,
  \3511(1567) ,
  \7344(2203) ,
  \4896(1445) ,
  \5959(2797) ,
  \7388(1283) ,
  \7220(1633) ,
  \887(922) ,
  \2553(3012) ,
  \1794(1510) ,
  \5198(1461) ,
  \940(2107) ,
  \4530(1185) ,
  \5715(3484) ,
  \1330(3067) ,
  \7330(1067) ,
  \7544(1345) ,
  \5116(2840) ,
  \2841(3662) ,
  \1903(1826) ,
  \5165(3600) ,
  \4737(3220) ,
  \1654(1538) ,
  \6934(3003) ,
  \4844(2345) ,
  \5767(473) ,
  \7283(1294) ,
  \6530(1053) ,
  \3462(3197) ,
  \6001(340) ,
  \3223(1698) ,
  \5828(2003) ,
  \1804(1513) ,
  \2598(1490) ,
  \4633(2978) ,
  \3606(2966) ,
  \6402(951) ,
  \4586(2182) ,
  \5297(1062) ,
  \6581(433) ,
  \2069(968) ,
  \7534(1348) ,
  \6615(331) ,
  \5308(846) ,
  \7268(1046) ,
  \3050(1903) ,
  \3751(229) ,
  \3071(2195) ,
  \2618(1985) ,
  \325(3358) ,
  \3504(1851) ,
  \3308(1109) ,
  \5464(1246) ,
  \2541(2918) ,
  \6233(3613) ,
  \4196(1605) ,
  \4538(1540) ,
  \1968(3163) ,
  \6661(2768) ,
  \4973(1548) ,
  \3441(2240) ,
  \4632(2731) ,
  \3030(2055) ,
  \4502(1015) ,
  \4824(2593) ,
  \6300(3453) ,
  \4517(3156) ,
  \6986(2769) ,
  \1761(3562) ,
  \6901(332) ,
  \[37] ,
  \6073(3150) ,
  \5505(3480) ,
  \5274(864) ,
  \1742(2065) ,
  \1093(1853) ,
  \2551(2921) ,
  \7352(2464) ,
  \2963(1741) ,
  \4653(410) ,
  \4089(2553) ,
  \2561(2925) ,
  \3574(2438) ,
  \6310(3500) ,
  \2555(2627) ,
  \4144(706) ,
  \4775(3303) ,
  \5832(2381) ,
  \[41] ,
  \[42] ,
  \5543(3212) ,
  \[43] ,
  \360(3379) ,
  \5014(2482) ,
  \5481(3105) ,
  \6503(1315) ,
  \[44] ,
  \6859(431) ,
  \2499(2782) ,
  \[45] ,
  \1102(940) ,
  \4920(565) ,
  \2008(3214) ,
  \6253(3645) ,
  \1573(1810) ,
  \[48] ,
  \6736(1629) ,
  \5740(3694) ,
  \[49] ,
  \2999(1578) ,
  \965(2958) ,
  \1841(883) ,
  \1994(2945) ,
  \5903(457) ,
  \1122(2101) ,
  \2515(2628) ,
  \6450(1017) ,
  \3009(1828) ,
  \4429(213) ,
  \1319(2883) ,
  \5508(2001) ,
  \929(2433) ,
  \1263(1857) ,
  \7273(1258) ,
  \[50] ,
  \745(853) ,
  \5362(1956) ,
  \[51] ,
  \6975(3549) ,
  \[52] ,
  \657(404) ,
  \[53] ,
  \6162(2604) ,
  \[55] ,
  \7290(1600) ,
  \[56] ,
  \2366(1130) ,
  \[57] ,
  \390(2934) ,
  \6281(3209) ,
  \[58] ,
  \3431(2229) ,
  \3393(1121) ,
  \4903(671) ,
  \[59] ,
  \5099(1218) ,
  \1350(415) ,
  \4122(751) ,
  \3908(1118) ,
  \5944(2606) ,
  \7334(1422) ,
  \3534(1882) ,
  \6040(1710) ,
  \5253(1453) ,
  \6931(1471) ,
  \2000(2667) ,
  \2353(1785) ,
  \731(855) ,
  \7197(3642) ,
  \[60] ,
  \4053(2910) ,
  \4287(2457) ,
  \[61] ,
  \1947(2035) ,
  \[62] ,
  \5788(964) ,
  \3813(822) ,
  \6461(1676) ,
  \[63] ,
  \6270(2986) ,
  \4598(2042) ,
  \[64] ,
  \4999(3047) ,
  \[65] ,
  \4873(373) ,
  \6519(928) ,
  \[66] ,
  \5884(1255) ,
  \5518(2011) ,
  \7041(1127) ,
  \3476(2903) ,
  \[67] ,
  \7324(1426) ,
  \4388(2971) ,
  \2050(656) ,
  \[68] ,
  \5873(338) ,
  \5512(2377) ,
  \[69] ,
  \5170(3696) ,
  \4166(995) ,
  \3109(1892) ,
  \7417(1349) ,
  \1783(3615) ,
  \1973(3167) ,
  \4622(2673) ,
  \7094(2263) ,
  \5745(353) ,
  \2434(1503) ,
  \6191(3208) ,
  \5189(607) ,
  \5342(1079) ,
  \7377(1347) ,
  \2064(675) ,
  \1399(820) ,
  \6165(3554) ,
  \7023(3493) ,
  \1172(3419) ,
  \5630(3482) ,
  \[70] ,
  \627(535) ,
  \1677(909) ,
  \[71] ,
  \708(641) ,
  \245(2897) ,
  \[72] ,
  \7549(1913) ,
  \2150(680) ,
  \4475(695) ,
  \[73] ,
  \5305(845) ,
  \5452(1077) ,
  \[74] ,
  \5352(1088) ,
  \[75] ,
  \[76] ,
  \6650(2228) ,
  \5292(1056) ,
  \4067(3144) ,
  \[77] ,
  \2398(1497) ,
  \[78] ,
  \1328(3191) ,
  \369(3714) ,
  \[79] ,
  \3590(2717) ,
  \1962(2086) ,
  \986(3677) ,
  \5522(2389) ,
  \6274(2812) ,
  \6990(2904) ,
  \2207(272) ,
  \6843(3118) ,
  \3650(666) ,
  \4233(1576) ,
  \7539(1916) ,
  \5412(1076) ,
  \7375(1682) ,
  \5502(2395) ,
  \[80] ,
  \1726(2407) ,
  \6526(1418) ,
  \6566(1414) ,
  \[81] ,
  \1454(2894) ,
  \[82] ,
  \7137(2780) ,
  \[83] ,
  \4815(3325) ,
  \5584(2419) ,
  \3653(506) ,
  \3080(1920) ,
  \5135(3409) ,
  \[84] ,
  \6304(2370) ,
  \[85] ,
  \914(1200) ,
  \6501(1645) ,
  \[86] ,
  \1003(3702) ,
  \7252(825) ,
  \308(3346) ,
  \[87] ,
  \7466(771) ,
  \7071(3378) ,
  \4804(2266) ,
  \1364(519) ,
  \5460(967) ,
  \[88] ,
  \6361(2702) ,
  \7011(3373) ,
  \[89] ,
  \5983(1789) ,
  \6469(1642) ,
  \938(2111) ,
  \5493(3345) ,
  \5202(1089) ,
  \4201(1695) ,
  \4247(2477) ,
  \3060(1919) ,
  \2699(1505) ,
  \1216(1757) ,
  \5271(863) ,
  \5857(1159) ,
  \7486(1173) ,
  \[90] ,
  \5365(2218) ,
  \996(3683) ,
  \[91] ,
  \4047(2302) ,
  \1005(721) ,
  \2846(3623) ,
  \4326(1655) ,
  \5031(3178) ,
  \2855(3703) ,
  \6085(3384) ,
  \6278(2940) ,
  \1378(538) ,
  \1942(2018) ,
  \2431(1140) ,
  \[96] ,
  \[97] ,
  \[98] ,
  \5604(2414) ,
  \[99] ,
  \6837(3056) ,
  \5312(1061) ,
  \5587(1183) ,
  \2292(570) ,
  \3853(1108) ,
  \2391(1134) ,
  \3234(2137) ,
  \6590(1707) ,
  \3295(1965) ,
  \7415(1659) ,
  \3365(1973) ,
  \3480(2765) ,
  \5708(3399) ,
  \255(2990) ,
  \4628(2865) ,
  \2643(1990) ,
  \5409(356) ,
  \7107(3607) ,
  \1318(2535) ,
  \928(2126) ,
  \3783(622) ,
  \5809(369) ,
  \7114(2272) ,
  \4014(2241) ,
  \2780(2629) ,
  \3470(2758) ,
  \1132(2164) ,
  \2105(972) ,
  \358(3320) ,
  \4273(2968) ,
  \993(3406) ,
  \4039(2275) ,
  \4756(2139) ,
  \2756(2339) ,
  \5728(3540) ,
  \1054(1615) ,
  \1998(3036) ,
  \7584(1906) ,
  \948(2130) ,
  \7124(2270) ,
  \6647(2559) ,
  \4667(492) ,
  \7104(2279) ,
  \924(2441) ,
  \4792(2449) ,
  \3642(579) ,
  \2956(1802) ,
  \3615(3168) ,
  \3239(3025) ,
  \5847(2663) ,
  \7594(1904) ,
  \377(3153) ,
  \6324(2359) ,
  \3013(906) ,
  \5346(1434) ,
  \401(310) ,
  \3791(795) ,
  \4280(2872) ,
  \4957(3112) ,
  \4735(3280) ,
  \1518(278) ,
  \4336(2185) ,
  \2776(2349) ,
  \1816(875) ,
  \2964(1512) ,
  \7316(1231) ,
  \4863(2938) ,
  \6796(1590) ,
  \6203(3437) ,
  \4088(3688) ,
  \1707(2029) ,
  \6517(598) ,
  \6399(897) ,
  \699(527) ,
  \3810(823) ,
  \5775(474) ,
  \7084(2290) ,
  \4480(756) ,
  \3587(2489) ,
  \5358(1752) ,
  \1036(1210) ,
  \2766(2340) ,
  \7609(2507) ,
  \5677(2676) ,
  \4078(3680) ,
  \3456(2273) ,
  \4412(219) ,
  \4004(2224) ,
  \7142(2778) ,
  \4163(994) ,
  \2977(879) ,
  \4288(2846) ,
  \6802(1261) ,
  \1802(871) ,
  \2351(1128) ,
  \6806(1598) ,
  \1786(3686) ,
  \3446(2265) ,
  \6446(1332) ,
  \6429(1165) ,
  \6410(950) ,
  \4362(2468) ,
  \5416(1431) ,
  \3682(839) ,
  \1501(291) ,
  \5277(1102) ,
  \6623(333) ,
  \2922(609) ,
  \5553(3391) ,
  \6792(1252) ,
  \6039(463) ,
  \2506(2332) ,
  \5050(3414) ,
  \3868(1110) ,
  \5456(1432) ,
  \6776(1384) ,
  \5356(1443) ,
  \5060(3486) ,
  \6422(1226) ,
  \6780(1711) ,
  \6123(2926) ,
  \6724(979) ,
  \6389(1154) ,
  \1554(1153) ,
  \4275(2707) ,
  \5928(1709) ,
  \5296(1411) ,
  \4009(2256) ,
  \1176(1838) ,
  \4349(1400) ,
  \3487(2574) ,
  \6586(1378) ,
  \7129(1483) ,
  \6320(3556) ,
  \4752(2425) ,
  \7276(1247) ,
  \1746(2424) ,
  \7155(3255) ,
  \2674(1504) ,
  \6574(1667) ,
  \5206(1444) ,
  \3059(1330) ,
  \3436(2250) ,
  \4389(1405) ,
  \6243(3664) ,
  \1974(2382) ,
  \248(3306) ,
  \3461(2297) ,
  \6494(1632) ,
  \4825(3257) ,
  \5686(2830) ,
  \6067(3088) ,
  \5849(884) ,
  \4083(3628) ,
  \4044(2280) ,
  \2580(3145) ,
  \2886(425) ,
  \6662(2564) ,
  \6679(1469) ,
  \5972(2331) ,
  \3610(2873) ,
  \1722(2049) ,
  \943(2127) ,
  \3437(2551) ,
  \4325(1941) ,
  \4672(685) ,
  \1712(2014) ,
  \2302(727) ,
  \5513(3524) ,
  \7064(2585) ,
  \6867(434) ,
  \4380(2721) ,
  \4900(1093) ,
  \1292(2213) ,
  \6963(3474) ,
  \5689(3164) ,
  \685(588) ,
  \1730(2668) ,
  \4562(1895) ,
  \4956(1556) ,
  \7463(913) ,
  \1026(1842) ,
  \6076(3147) ,
  \6948(2260) ,
  \2077(973) ,
  \5620(3400) ,
  \7474(908) ,
  \5439(484) ,
  \3451(2283) ,
  \5573(3538) ,
  \1624(894) ,
  \1919(1188) ,
  \1035(925) ,
  \1091(1224) ;
assign
  \260(2889)  = \3249(2223)  & \3046(2813) ,
  \4872(2649)  = ~\4868(2371) ,
  \5531(2823)  = ~\5529(1519)  | ~\5526(2662) ,
  \1514(406)  = ~\1512(300) ,
  \7117(3661)  = ~\7111(3644) ,
  \7127(3660)  = ~\7121(3643) ,
  \7050(2914)  = ~\7048(2777)  | ~\7041(1127) ,
  \5796(960)  = \1412(818) ,
  \1037(1561)  = ~\5206(1444)  | ~\5199(377) ,
  \573(311)  = \1(0) ,
  \7368(1627)  = ~\7364(1292) ,
  \6732(1295)  = \2186(989) ,
  \5145(3488)  = ~\5139(3470) ,
  \7548(1683)  = ~\7544(1345) ,
  \4881(375)  = \1488(279) ,
  \5911(460)  = ~\5905(347) ,
  \7442(2814)  = ~\7438(2650) ,
  \336(3412)  = \[84] ,
  \1143(3177)  = \1074(1846)  & (\1093(1853)  & \3271(3101) ),
  \6538(1055)  = \637(842) ,
  \3228(2097)  = \3176(1840)  & (\3186(1845)  & (\3195(1876)  & (\3203(1847)  & \3215(1852) ))),
  \2049(803)  = \2026(730)  & \202(125) ,
  \4977(1835)  = ~\4973(1548) ,
  \6269(2878)  = ~\6267(2208)  | ~\6264(2640) ,
  \980(3210)  = ~\975(3157) ,
  \3216(1462)  = \3170(866)  & \3212(1367) ,
  \5753(354)  = \1186(254) ,
  \7070(3252)  = ~\7068(2775)  | ~\7061(3199) ,
  \4024(2268)  = \3926(1120)  & \3899(1971) ,
  \3119(2180)  = ~\3118(1644)  | ~\3117(1930) ,
  \2163(976)  = \2146(661)  | \2145(810) ,
  \4979(2200)  = ~\4977(1835)  | ~\4970(718) ,
  \2501(2335)  = \2354(1983)  & (\2391(1134)  & \2372(1986) ),
  \5107(2690)  = ~\5105(1569)  | ~\5102(2481) ,
  \2149(808)  = \2124(731)  & \195(118) ,
  \7538(1686)  = ~\7534(1348) ,
  \492(265)  = \2224(178) ,
  \4852(2352)  = \2420(1992) ,
  \315(3281)  = ~\4744(2423)  | ~\4737(3220) ,
  \3471(2997)  = ~\3470(2758)  | ~\3469(2900) ,
  \1721(2410)  = ~\1718(2046) ,
  \5682(2674)  = ~\1746(2424) ,
  \4993(1203)  = \887(922) ,
  \5937(2610)  = \2502(2317)  | (\2501(2335)  | (\2500(2322)  | \2366(1130) )),
  \3143(2738)  = \3142(2478)  | (\3141(2492)  | (\3140(2494)  | (\3139(2474)  | \3090(1356) ))),
  \1239(1734)  = ~\5288(1406)  | ~\5281(1058) ,
  \4175(1007)  = \4150(704)  | \4149(742) ,
  \3079(1370)  = \3804(833)  & \4166(995) ,
  \1781(3684)  = ~\1780(3674) ,
  \6535(984)  = \3673(821) ,
  \6458(1036)  = \3807(834) ,
  \6669(2767)  = ~\6663(2567) ,
  \4250(2709)  = ~\4247(2477) ,
  \6370(1065)  = \727(848) ,
  \3249(2223)  = \3228(2097)  & \3216(1462) ,
  \5261(1447)  = ~\5255(1092) ,
  \845(980)  = \2942(859)  & \1477(394) ,
  \4160(993)  = \4135(688)  | \4134(747) ,
  \5006(3226)  = ~\5000(3169) ,
  \275(3286)  = \908(1192)  & \958(3228) ,
  \6498(1032)  = \3804(833) ,
  \2930(613)  = \2929(516)  | \2914(591) ,
  \2055(785)  = \2039(737)  & \235(158) ,
  \4945(2743)  = ~\4939(2512) ,
  \2343(1982)  = ~\2342(1784)  | ~\2341(1488) ,
  \2481(1721)  = \4389(1405)  & \3682(839) ,
  \6103(3519)  = ~\6097(3498) ,
  \5881(341)  = \3739(233) ,
  \4221(2171)  = ~\4220(1619)  | ~\4219(1942) ,
  \4983(1191)  = ~\915(1029)  & ~\777(370) ,
  \1321(2460)  = \1300(2146)  & (\1263(1857)  & \1272(1858) ),
  \2872(430)  = ~\2871(315) ,
  \6972(2555)  = ~\6968(2226) ,
  \621(532)  = \587(402)  & \167(90) ,
  \356(3424)  = \[103] ,
  \2925(514)  = \2892(416)  & \214(137) ,
  \4291(2173)  = ~\4290(1911)  | ~\4289(1880) ,
  \2291(618)  = \2266(587)  & \206(129) ,
  \577(631)  = \615(529)  | \594(572) ,
  \7567(1310)  = \4163(994) ,
  \2938(860)  = \2886(425)  & \2922(609) ,
  \6093(3463)  = ~\6087(3435) ,
  \2511(2348)  = \2431(1140)  & \2409(1989) ,
  \7504(1150)  = ~\7500(873) ,
  \702(638)  = \701(541)  | \685(588) ,
  \2519(2361)  = \2420(1992)  & (\2465(1144)  & \2436(1993) ),
  \1372(522)  = \1336(405)  & \178(101) ,
  \6213(3510)  = ~\6212(3473)  | ~\6211(3491) ,
  \6012(1287)  = \2085(986) ,
  \348(3371)  = \3497(3319)  & \3482(3075) ,
  \6968(2226)  = \3845(1963) ,
  \4965(3227)  = ~\4959(3170) ,
  \1597(1527)  = ~\5424(1437)  | ~\5417(360) ,
  \6982(2565)  = ~\6978(2235) ,
  \5780(1081)  = \731(855) ,
  \5591(2952)  = ~\5590(2833)  | ~\5589(2677) ,
  \7272(1399)  = ~\7268(1046) ,
  \7482(898)  = \4695(767) ,
  \6036(1383)  = \2323(1038) ,
  \4341(1392)  = \2312(836)  & \4493(998) ,
  \6131(3149)  = ~\6125(3087) ,
  \6952(2576)  = ~\6948(2260) ,
  \4490(1000)  = \4475(695)  | \4474(759) ,
  \2226(264)  = ~\2224(178) ,
  \471(3445)  = \1175(3403) ,
  \6173(1723)  = ~\4389(1405)  & ~\3682(839) ,
  \1129(2434)  = \1128(2132)  | (\1127(2116)  | (\1126(2165)  | (\1125(2104)  | \1035(925) ))),
  \6896(1302)  = \2192(991) ,
  \4290(1911)  = ~\7368(1627)  | ~\7361(1343) ,
  \1092(1572)  = ~\5230(1455)  | ~\5223(382) ,
  \7227(1358)  = ~\7221(1020) ,
  \4239(2141)  = ~\4235(1855) ,
  \6471(1307)  = \4160(993) ,
  \5138(3413)  = ~\5136(2453)  | ~\5129(3359) ,
  \442(280)  = \1486(171) ,
  \4635(2727)  = \4614(2495)  & (\4577(2183)  & \4586(2182) ),
  \7228(1606)  = ~\7224(1270) ,
  \395(3023)  = ~\4871(2985)  | ~\4868(2371) ,
  \3081(1641)  = ~\6470(1357)  | ~\6463(1309) ,
  \6884(1694)  = ~\6880(1361) ,
  \6527(932)  = \3676(777) ,
  \2171(992)  = \2150(680)  | \2149(808) ,
  \3661(496)  = \3635(408)  & \1495(276) ,
  \6962(2572)  = ~\6958(2248) ,
  \2546(3010)  = ~\2545(2787)  | ~\2544(2919) ,
  \6924(1613)  = ~\6920(1276) ,
  \7471(902)  = \4692(768) ,
  \4716(2094)  = \1921(1832) ,
  \2851(3008)  = \2757(2602)  & \2809(2893) ,
  \6163(3534)  = ~\6161(3520)  | ~\6158(2308) ,
  \1333(3069)  = ~\5392(2885)  | ~\5385(2962) ,
  \6347(3057)  = ~\4273(2968)  | ~\4276(2967) ,
  \5417(360)  = \1178(261) ,
  \3135(2868)  = ~\3131(2733) ,
  \5718(3483)  = ~\5716(2427)  | ~\5709(3467) ,
  \4434(211)  = ~\4432(203) ,
  \5529(1519)  = ~\5523(1158) ,
  \2852(2785)  = \2771(2634)  & \2749(2307) ,
  \1745(2084)  = \1677(909)  & \1655(1827) ,
  \6978(2235)  = \3856(1966) ,
  \4988(2834)  = ~\4986(2742)  | ~\4983(1191) ,
  \1198(299)  = \38(11) ,
  \3151(2974)  = ~\3127(2725)  | ~\3135(2868) ,
  \1326(3135)  = ~\5375(3070)  | ~\5372(1759) ,
  \1902(1537)  = ~\5808(1237)  | ~\5801(366) ,
  \276(3401)  = \[76] ,
  \4522(3128)  = ~\7462(2981)  | ~\7453(3062) ,
  \1735(2080)  = \1609(1820)  & (\1677(909)  & (\1630(1824)  & \1655(1827) )),
  \7069(3323)  = ~\7067(3256)  | ~\7064(2585) ,
  \1725(2081)  = \1609(1820)  & (\1677(909)  & (\1598(1817)  & (\1630(1824)  & \1655(1827) ))),
  \298(3387)  = \[87] ,
  \1184(294)  = \133(66)  & \134(67) ,
  \6958(2248)  = \3874(1968) ,
  \3351(1476)  = ~\6605(440)  | ~\6602(1359) ,
  \7044(2590)  = \4044(2280)  | (\4043(2301)  | (\4042(2289)  | \3949(1122) )),
  \284(384)  = \[48] ,
  \2789(2365)  = \2655(1991)  & (\2715(1145)  & \2676(1994) ),
  \5783(479)  = ~\5777(361) ,
  \3270(2892)  = \1974(2382)  & (\3466(2558)  & (\2532(2788)  & \4526(205) )),
  \4179(1608)  = ~\7212(1277)  | ~\7205(1273) ,
  \4897(548)  = \1477(394) ,
  \4636(2976)  = ~\4635(2727)  & ~\4634(2863) ,
  \2849(3692)  = \2839(3690)  & \2828(208) ,
  \5029(3114)  = ~\5027(3053)  | ~\5024(2689) ,
  \2839(3690)  = ~\2838(3672)  | ~\2837(3682) ,
  \6744(1601)  = ~\6740(1265) ,
  \7291(1868)  = ~\7289(1628)  | ~\7286(1264) ,
  \1322(2847)  = ~\1321(2460)  & ~\1320(2696) ,
  \6357(3063)  = ~\4279(2982)  | ~\4282(2983) ,
  \4187(1884)  = ~\7219(1638)  | ~\7216(1300) ,
  \7009(3312)  = ~\7003(3247) ,
  \7281(1860)  = ~\7279(1595)  | ~\7276(1247) ,
  \5007(1201)  = ~\5003(920) ,
  \2544(2919)  = ~\5951(2790)  | ~\5948(2311) ,
  \1226(1959)  = ~\1225(1755)  | ~\1224(1756) ,
  \4675(482)  = \4640(409)  & \2232(262) ,
  \6909(324)  = \4422(215) ,
  \313(3396)  = \[78] ,
  \3281(1464)  = ~\6573(432)  | ~\6570(1329) ,
  \4911(507)  = ~\4905(380) ,
  \2914(591)  = ~\2909(417) ,
  \1320(2696)  = \1303(2462)  & (\1272(1858)  & \1267(2144) ),
  \328(3361)  = ~\4775(3303)  | ~\4772(2105) ,
  \7293(953)  = \1383(815) ,
  \6374(1420)  = ~\6370(1065) ,
  \2564(2929)  = \2563(2756)  | \2515(2628) ,
  \4785(3237)  = \1145(3179)  | \1102(940) ,
  \6153(3479)  = ~\6151(3462)  | ~\6148(2329) ,
  \1556(1807)  = ~\1555(1514)  | ~\1554(1153) ,
  \6614(1602)  = ~\6610(1266) ,
  \1112(1553)  = ~\1108(1196) ,
  \1546(1803)  = ~\1545(1509)  | ~\1544(1148) ,
  \339(164)  = \IN-339(164) ,
  \4443(3309)  = \3621(3240)  & (\3618(3244)  & (\1334(3190)  & \1328(3191) )),
  \2117(577)  = \1514(406) ,
  \1572(1517)  = ~\5416(1431)  | ~\5409(356) ,
  \4505(1014)  = \4485(711)  | \4484(754) ,
  \3745(231)  = ~\3743(193) ,
  \1369(646)  = \1343(575)  & \144(71) ,
  \1300(2146)  = \1281(1859) ,
  \4090(2757)  = \4028(2579)  & \4004(2224) ,
  \1206(306)  = ~\9(2)  | ~\12(3) ,
  \3019(1581)  = ~\6437(1187)  | ~\6434(954) ,
  \4871(2985)  = ~\4865(2877) ,
  \3444(2246)  = \3314(1967)  & \3344(1970) ,
  \5122(2443)  = ~\943(2127)  & (~\942(2110)  & (~\941(2161)  & ~\821(929) )),
  \3376(1119)  = \2198(974)  & \4412(219) ,
  \5825(2383)  = ~\1946(2033)  & (~\1945(2019)  & ~\1816(875) ),
  \7185(3553)  = ~\7179(3533) ,
  \3609(2984)  = ~\3608(2741)  & ~\3607(2875) ,
  \6631(334)  = \4396(225) ,
  \7138(2913)  = ~\7136(2776)  | ~\7129(1483) ,
  \3352(1773)  = ~\6606(1692)  | ~\6599(327) ,
  \6240(2643)  = ~\6236(2360) ,
  \5255(1092)  = \2942(859) ,
  \3282(1763)  = ~\6574(1667)  | ~\6567(319) ,
  \3434(2230)  = \3308(1109)  & \3283(1964) ,
  \7562(1314)  = \4154(996) ,
  \4372(2520)  = \4333(1397)  & \4317(2170) ,
  \6509(1649)  = ~\6503(1315) ,
  \2494(2333)  = \2354(1983)  & (\2391(1134)  & (\2343(1982)  & \2372(1986) )),
  \6009(345)  = \3725(237) ,
  \3488(2771)  = ~\6686(2570)  | ~\6679(1469) ,
  \5484(3103)  = ~\5482(2661)  | ~\5475(3038) ,
  \2532(2788)  = \2508(2630)  & \2487(2312) ,
  \3526(1610)  = ~\6728(1278)  | ~\6721(1274) ,
  \1125(2104)  = \1050(930)  & \1026(1842) ,
  \6047(455)  = ~\6041(342) ,
  \7337(1902)  = ~\7248(1668)  | ~\7247(1691) ,
  \6220(2646)  = ~\6216(2369) ,
  \2542(2786)  = ~\5944(2606)  | ~\5937(2610) ,
  \300(3267)  = \1994(2945)  & \2008(3214) ,
  \4760(2455)  = ~\4756(2139) ,
  \1997(2944)  = ~\1996(2658)  | ~\1995(2819) ,
  \4904(1448)  = ~\4900(1093) ,
  \3731(235)  = ~\3729(191) ,
  \2816(3019)  = ~\2813(2930) ,
  \6589(435)  = ~\6583(322) ,
  \975(3157)  = \1447(3100) ,
  \693(524)  = \657(404)  & \176(99) ,
  \6182(3065)  = ~\6180(2936)  | ~\6173(1723) ,
  \7286(1264)  = \2077(973) ,
  \6260(2636)  = ~\6256(2350) ,
  \3567(1878)  = ~\6788(1719)  | ~\6781(1286) ,
  \7496(1516)  = ~\7494(1164)  | ~\7487(881) ,
  \5183(498)  = \1519(374) ,
  \3608(2741)  = \3587(2489)  & (\3550(2199)  & \3559(2205) ),
  \2099(970)  = \2060(655)  | \2059(787) ,
  \6250(2638)  = ~\6246(2351) ,
  \3622(407)  = \1524(301) ,
  \2854(2916)  = \2853(2784)  | \2757(2602) ,
  \2508(2630)  = \2454(1996)  & (\2409(1989)  & (\2436(1993)  & (\2472(2532)  & \2420(1992) ))),
  \5776(1433)  = ~\5772(1078) ,
  \6230(2633)  = ~\6226(2347) ,
  \6294(2746)  = \2742(2533) ,
  \1987(2942)  = ~\1986(2653)  | ~\1985(2817) ,
  \2768(2619)  = \2767(2341)  | \2629(1133) ,
  \587(402)  = \1512(300) ,
  \1776(3649)  = ~\5658(2417)  | ~\5651(3638) ,
  \6875(436)  = ~\6869(323) ,
  \1750(2078)  = \1655(1827)  & \1695(1829) ,
  \2753(2603)  = ~\2749(2307) ,
  \5492(2402)  = ~\5488(2039) ,
  \393(2937)  = ~\4864(2641)  | ~\4857(2810) ,
  \2571(3018)  = ~\2564(2929) ,
  \5178(399)  = \1198(299) ,
  \1740(2071)  = \1669(904)  & \1630(1824) ,
  \4585(1908)  = ~\7566(1648)  | ~\7559(1340) ,
  \4575(1909)  = ~\7557(1651)  | ~\7554(1011) ,
  \2520(2522)  = \2420(1992)  & (\2481(1721)  & (\2436(1993)  & \2454(1996) )),
  \2800(2530)  = \2724(1722)  & \2701(1995) ,
  \7490(887)  = \4701(765) ,
  \1766(3073)  = \1454(2894)  | (\1450(2996)  | \4091(2899) ),
  \7021(3475)  = ~\7019(3456)  | ~\7016(2249) ,
  \7081(3477)  = ~\7080(3433)  | ~\7079(3459) ,
  \2552(2794)  = ~\5968(2613)  | ~\5961(2617) ,
  \4680(683)  = \4660(581)  & \86(45) ,
  \7256(1022)  = ~\7252(825) ,
  \2085(986)  = \2056(674)  | \2055(785) ,
  \3489(2906)  = ~\3488(2771)  | ~\3487(2574) ,
  \6598(1704)  = ~\6594(1375) ,
  \4368(2855)  = ~\4364(2720) ,
  \6702(1216)  = ~\6698(938) ,
  \363(3380)  = ~\4823(3327)  | ~\4820(2281) ,
  \1336(405)  = \1512(300) ,
  \5967(2796)  = ~\5961(2617) ,
  \1014(560)  = \1519(374)  & \1198(299) ,
  \6856(1327)  = \3838(1004) ,
  \5539(3104)  = ~\5533(3037) ,
  \4745(3222)  = \1973(3167)  | \1929(910) ,
  \5503(3465)  = ~\5501(3441)  | ~\5498(2023) ,
  \3469(2900)  = ~\6645(2762)  | ~\6642(2227) ,
  \4590(2499)  = ~\4586(2182) ,
  \3061(1672)  = ~\6454(1354)  | ~\6447(1335) ,
  \3035(2374)  = \3029(2043)  & \3022(1998) ,
  \3479(2902)  = ~\6669(2767)  | ~\6666(2232) ,
  \3807(834)  = \3786(568)  | \3785(623) ,
  \5599(3107)  = ~\5597(3043)  | ~\5594(2675) ,
  \7396(1045)  = \2316(837) ,
  \1921(1832)  = ~\1920(1544)  | ~\1919(1188) ,
  \6992(3002)  = ~\6990(2904)  | ~\6983(1470) ,
  \7296(811)  = \1364(519)  | \1363(647) ,
  \5924(1382)  = \2323(1038) ,
  \3051(1669)  = ~\6446(1332)  | ~\6439(1333) ,
  \6825(2469)  = ~\6819(2152) ,
  \6658(2233)  = \3295(1965) ,
  \7248(1668)  = ~\7246(1355)  | ~\7239(1005) ,
  \4485(711)  = \4457(583)  & \54(17) ,
  \4149(742)  = \4114(735)  & \4439(209) ,
  \2616(1491)  = ~\6007(453)  | ~\6004(1254) ,
  \3490(3195)  = \2580(3145)  & \3446(2265) ,
  \2124(731)  = ~\2117(577) ,
  \5836(2008)  = \1805(1806) ,
  \4017(2569)  = \4016(2258)  | \3885(1112) ,
  \5761(357)  = \2249(255) ,
  \5447(487)  = ~\5441(367) ,
  \4496(999)  = \4479(694)  | \4478(757) ,
  \7469(1186)  = ~\7463(913) ,
  \5432(1242)  = ~\5428(963) ,
  \3033(2092)  = \2992(1821)  & (\3015(912)  & (\2982(1816)  & (\3001(1823)  & \3009(1828) ))),
  \3527(2160)  = ~\3526(1610)  | ~\3525(1873) ,
  \955(3172)  = ~\1447(3100)  | ~\920(2100) ,
  \7100(3551)  = ~\7098(2581)  | ~\7091(3532) ,
  \1955(2073)  = \1869(1819)  & (\1914(905)  & (\1859(1818)  & \1885(1825) )),
  \5521(3560)  = ~\5515(3539) ,
  \2790(2526)  = \2655(1991)  & (\2724(1722)  & (\2676(1994)  & \2701(1995) )),
  \550(236)  = \3729(191) ,
  \1965(2074)  = \1885(1825)  & \1914(905) ,
  \1436(3029)  = \1788(2375)  & \4091(2899) ,
  \601(422)  = \1206(306) ,
  \6511(429)  = \2883(314) ,
  \4605(2405)  = ~\4602(2041) ,
  \6057(1136)  = ~\2091(969)  & ~\3731(235) ,
  \6941(3141)  = ~\6935(3077) ,
  \7060(3079)  = ~\7058(2912)  | ~\7051(3007) ,
  \989(3676)  = ~\988(3652)  | ~\987(3667) ,
  \4625(2678)  = \4605(2405)  & (\4544(2062)  & \4531(1830) ),
  \5210(1094)  = \2942(859) ,
  \3600(2838)  = ~\3599(2436)  & ~\3598(2692) ,
  \3279(3072)  = \3277(2891)  | (\3274(2999)  | \3468(2898) ),
  \6933(2908)  = ~\6931(1471)  | ~\6928(2770) ,
  \375(3090)  = \2543(3009)  & \2564(2929) ,
  \4567(2501)  = ~\4563(2184) ,
  \4258(2716)  = ~\4255(2488) ,
  \2272(594)  = \1507(418) ,
  \5175(372)  = \1541(275) ,
  \6788(1719)  = ~\6784(1396) ,
  \5641(3583)  = ~\5640(3541)  | ~\5639(3564) ,
  \2749(2307)  = \2589(1981)  & (\2600(1984)  & (\2618(1985)  & \2734(1987) )),
  \2144(663)  = \2117(577)  & \115(60) ,
  \2971(1744)  = ~\6389(1154)  | ~\6386(1069) ,
  \2058(654)  = \2032(592)  & \130(65) ,
  \3130(2513)  = \3062(2194)  & (\3079(1370)  & (\3052(2192)  & \3071(2195) )),
  \5563(3481)  = ~\5562(3439)  | ~\5561(3466) ,
  \1170(3367)  = \1166(3292)  & \1158(1927) ,
  \4832(2597)  = ~\4828(2293) ,
  \4919(605)  = ~\4913(497) ,
  \3658(681)  = \3642(579)  & \88(47) ,
  \5482(2661)  = ~\5478(2388) ,
  \1982(2816)  = \1981(2655)  | \1941(2379) ,
  \3695(1050)  = \2305(826)  & \1535(302) ,
  \7433(2949)  = ~\4624(2829)  | ~\4627(2827) ,
  \6241(3646)  = ~\6239(3633)  | ~\6236(2360) ,
  \1544(1148)  = ~\5399(466)  | ~\5396(1084) ,
  \6567(319)  = \4439(209) ,
  \2143(806)  = \2124(731)  & \197(120) ,
  \323(3238)  = ~\4760(2455)  | ~\4753(3158) ,
  \6973(3531)  = ~\6971(3513)  | ~\6968(2226) ,
  \3142(2478)  = \3093(2156)  & (\3116(1271)  & (\3082(2179)  & (\3102(2177)  & \3110(2175) ))),
  \1960(2059)  = \1897(900)  & \1869(1819) ,
  \3620(3117)  = ~\6852(2965)  | ~\6845(3058) ,
  \1503(303)  = \18(5) ,
  \5840(2386)  = ~\5836(2008) ,
  \7159(3377)  = ~\7158(3251)  | ~\7157(3322) ,
  \7172(2291)  = \3957(1977) ,
  \2063(789)  = \2039(737)  & \231(154) ,
  \5119(3175)  = ~\5118(3050)  | ~\5117(3113) ,
  \5952(2607)  = ~\5948(2311) ,
  \1945(2019)  = \1834(878)  & \1805(1806) ,
  \2296(715)  = \2272(594)  & \44(13) ,
  \917(1190)  = \916(1030)  | \777(370) ,
  \1281(1859)  = ~\1280(1751)  | ~\1279(1585) ,
  \2371(1788)  = ~\5888(1593)  | ~\5881(341) ,
  \7145(3080)  = ~\7139(3006) ,
  \7003(3247)  = ~\7002(3138)  | ~\7001(3193) ,
  \624(635)  = \623(533)  | \611(573) ,
  \3168(828)  = ~\6517(598)  | ~\6514(397) ,
  \3207(936)  = \633(843)  & \3670(778) ,
  \710(642)  = \709(545)  | \685(588) ,
  \6070(2612)  = \2764(2319)  | (\2763(2338)  | (\2762(2326)  | \2612(1131) )),
  \7221(1020)  = \3801(824) ,
  \926(2163)  = \845(980)  & (\792(1841)  & \805(1844) ),
  \6251(3634)  = ~\6327(3612)  | ~\6324(2359) ,
  \997(2432)  = \920(2100)  & \902(1199) ,
  \4278(2739)  = \4255(2488)  & (\4203(1923)  & \4212(1937) ),
  \6853(318)  = \4439(209) ,
  \1024(1209)  = ~\5197(501)  | ~\5194(1106) ,
  \2946(858)  = \2886(425)  & \2926(611) ,
  \5021(2960)  = ~\5020(2844)  | ~\5019(2691) ,
  \5112(2687)  = ~\950(2448) ,
  \2384(1132)  = \2099(970)  & \3739(233) ,
  \2005(2824)  = ~\2004(2666)  | ~\2003(2399) ,
  \5566(2000)  = \1546(1803) ,
  \3559(2205)  = ~\3558(1938)  | ~\3557(1935) ,
  \3245(3230)  = \3243(3171)  & \3238(2684) ,
  \5570(2376)  = ~\5566(2000) ,
  \707(544)  = \678(414)  & \154(77) ,
  \3548(1924)  = ~\6771(1697)  | ~\6768(1023) ,
  \3473(2759)  = ~\6654(2557)  | ~\6647(2559) ,
  \4520(3243)  = ~\4519(3124)  | ~\4518(3183) ,
  \3614(3044)  = ~\6836(1833)  | ~\6829(2957) ,
  \2819(3610)  = ~\2818(3575)  | ~\2817(3590) ,
  \711(852)  = \650(423)  & \692(626) ,
  \1992(2820)  = ~\5839(2664)  | ~\5836(2008) ,
  \2676(1994)  = ~\2675(1798)  | ~\2674(1504) ,
  \4276(2967)  = ~\4275(2707)  & ~\4274(2852) ,
  \5017(1219)  = ~\5011(941) ,
  \4058(3569)  = ~\6982(2565)  | ~\6975(3549) ,
  \4935(722)  = ~\4929(564) ,
  \7047(1485)  = ~\7041(1127) ,
  \5420(1082)  = \731(855) ,
  \1530(411)  = ~\1524(301) ,
  \4908(1096)  = \2938(860) ,
  \2286(554)  = \2259(413)  & \44(13) ,
  \6083(3332)  = ~\6077(3261) ,
  \1418(819)  = \1382(540)  | \1381(651) ,
  \4007(2231)  = \3868(1110)  & \3845(1963) ,
  \2158(677)  = \2130(593)  & \97(50) ,
  \1157(1699)  = ~\5246(1194)  | ~\5239(719) ,
  \5491(3269)  = ~\5485(3213) ,
  \6514(397)  = \1210(298) ,
  \5892(1250)  = \2091(969) ,
  \984(3668)  = ~\5087(3655)  | ~\5084(2108) ,
  \6851(3120)  = ~\6845(3058) ,
  \478(269)  = \2211(176) ,
  \270(3109)  = \[60] ,
  \3926(1120)  = \2198(974)  & \4412(219) ,
  \2452(1506)  = ~\5927(464)  | ~\5924(1382) ,
  \3854(1466)  = ~\6867(434)  | ~\6864(1352) ,
  \337(3712)  = ~\1004(3708)  | ~\1003(3702) ,
  \7423(1687)  = ~\7417(1349) ,
  \3909(1478)  = ~\6891(442)  | ~\6888(1267) ,
  \6534(1408)  = ~\6530(1053) ,
  \450(288)  = \1459(167) ,
  \5576(2013)  = \1556(1807) ,
  \6362(2849)  = ~\6361(2702)  | ~\6360(2697) ,
  \3558(1938)  = ~\6780(1711)  | ~\6773(1388) ,
  \7058(2912)  = ~\7054(2779) ,
  \5425(363)  = \2232(262) ,
  \4255(2488)  = \4221(2171) ,
  \3503(1221)  = ~\6694(945)  | ~\6687(943) ,
  \3465(3201)  = \3417(1979)  & \2580(3145) ,
  \1380(539)  = \1350(415)  & \159(82) ,
  \7376(1599)  = ~\7372(1263) ,
  \6953(3374)  = ~\6951(3313)  | ~\6948(2260) ,
  \6360(2697)  = ~\7351(2471)  | ~\7348(2148) ,
  \1234(1760)  = ~\5270(1446)  | ~\5263(1104) ,
  \1971(3165)  = \1903(1826)  & (\1921(1832)  & \3279(3072) ),
  \5061(3527)  = ~\5060(3486)  | ~\5059(3507) ,
  \6558(556)  = ~\6554(396) ,
  \3796(725)  = \3768(595)  & \32(9) ,
  \3804(833)  = \3784(567)  | \3783(622) ,
  \3210(1026)  = ~\6557(741)  | ~\6554(396) ,
  \7000(2763)  = ~\6996(2561) ,
  \6479(1339)  = \4157(1010) ,
  \2220(266)  = ~\2218(177) ,
  \6223(3557)  = ~\6222(3521)  | ~\6221(3536) ,
  \5560(2396)  = ~\5556(2024) ,
  \7383(1685)  = ~\7377(1347) ,
  \5556(2024)  = \1573(1810) ,
  \6439(1333)  = \4175(1007) ,
  \5743(3647)  = ~\5737(3636) ,
  \633(843)  = \581(421)  & \618(632) ,
  \4839(316)  = ~\4833(207) ,
  \6378(1066)  = \723(849) ,
  \2863(3127)  = ~\6356(2869)  | ~\6347(3057) ,
  \4189(2176)  = ~\4188(1887)  | ~\4187(1884) ,
  \4764(2102)  = \1026(1842) ,
  \528(214)  = \4427(202) ,
  \6113(3574)  = ~\6107(3555) ,
  \3786(568)  = \3755(412)  & \32(9) ,
  \3799(799)  = \3775(740)  & \219(142) ,
  \4146(743)  = \4114(735)  & \4434(211) ,
  \7618(2498)  = ~\7614(2181) ,
  \5580(2390)  = ~\5576(2013) ,
  \958(3228)  = \955(3172)  & \933(2683) ,
  \4493(998)  = \4477(693)  | \4476(758) ,
  \5855(1161)  = ~\5849(884) ,
  \5549(3268)  = ~\5543(3212) ,
  \6768(1023)  = \2296(715)  | \2295(781) ,
  \5300(1052)  = \641(841) ,
  \4141(690)  = \4107(585)  & \79(38) ,
  \3855(1765)  = ~\6868(1690)  | ~\6861(321) ,
  \7158(3251)  = ~\7156(2774)  | ~\7149(3198) ,
  \3449(2267)  = \3376(1119)  & \3353(1972) ,
  \4812(2269)  = \3365(1973) ,
  \5546(2038)  = \1687(1813) ,
  \4823(3327)  = ~\4817(3254) ,
  \7506(1507)  = ~\7504(1150)  | ~\7497(868) ,
  \1495(276)  = ~\1492(172) ,
  \6477(1639)  = ~\6471(1307) ,
  \4488(752)  = \4464(733)  & \3751(229) ,
  \1224(1756)  = ~\5261(1447)  | ~\5258(1097) ,
  \3439(2252)  = \3295(1965)  & (\3335(1113)  & \3314(1967) ),
  \7245(1331)  = ~\7239(1005) ,
  \1377(649)  = \1357(589)  & \138(69) ,
  \346(3311)  = \3471(2997)  & \3491(3249) ,
  \1154(1928)  = ~\1153(1700)  | ~\1152(1369) ,
  \6655(2568)  = \3444(2246)  | (\3443(2253)  | \3327(1111) ),
  \2844(3625)  = \2833(317)  & (\2784(2802)  & \2824(3611) ),
  \5197(501)  = ~\5191(376) ,
  \4086(3630)  = \4067(3144)  & (\4056(3005)  & \4059(3604) ),
  \5791(480)  = ~\5785(362) ,
  \5027(3053)  = ~\5021(2960) ,
  \5672(2418)  = ~\1744(2085)  & (~\1743(2070)  & ~\1647(899) ),
  \2775(2803)  = ~\2771(2634) ,
  \902(1199)  = \765(774)  & \887(922) ,
  \1867(1170)  = ~\5791(480)  | ~\5788(964) ,
  \6845(3058)  = ~\3609(2984)  | ~\3612(2970) ,
  \946(2122)  = \853(1849)  & (\827(1874)  & \895(1850) ),
  \7385(1324)  = \4499(1001) ,
  \6597(438)  = ~\6591(325) ,
  \296(3340)  = \2014(3274)  & \1991(3031) ,
  \7494(1164)  = ~\7490(887) ,
  \1999(2400)  = ~\5855(1161)  | ~\5852(2026) ,
  \4683(468)  = \4653(410)  & \2255(252) ,
  \7195(3606)  = ~\7189(3588) ,
  \4720(2430)  = ~\4716(2094) ,
  \5692(2413)  = ~\1739(2082)  & (~\1738(2067)  & (~\1737(2056)  & ~\1624(894) )),
  \5465(885)  = ~\737(854)  & ~\2241(257) ,
  \5748(1085)  = \757(856) ,
  \2599(1786)  = ~\6000(1597)  | ~\5993(339) ,
  \696(628)  = \695(525)  | \664(574) ,
  \419(3444)  = \1175(3403) ,
  \1857(1169)  = ~\5783(479)  | ~\5780(1081) ,
  \7573(1643)  = ~\7567(1310) ,
  \5804(958)  = \1406(817) ,
  \941(2161)  = \845(980)  & \805(1844) ,
  \3353(1972)  = ~\3352(1773)  | ~\3351(1476) ,
  \2878(386)  = \1501(291)  & \4442(290) ,
  \3283(1964)  = ~\3282(1763)  | ~\3281(1464) ,
  \4063(3570)  = ~\7040(2566)  | ~\7033(3548) ,
  \7182(2262)  = \3899(1971) ,
  \1705(2010)  = \1567(876)  & \1546(1803) ,
  \7299(1232)  = ~\7293(953) ,
  \956(2124)  = \853(1849)  & \895(1850) ,
  \1363(647)  = \1343(575)  & \141(70) ,
  \5609(3277)  = ~\5607(3221)  | ~\5604(2414) ,
  \1156(1368)  = ~\5245(830)  | ~\5242(917) ,
  \6836(1833)  = ~\6832(1546) ,
  \5071(3585)  = ~\5070(3545)  | ~\5069(3566) ,
  \4270(2459)  = ~\4267(2143) ,
  \263(2858)  = \3249(2223)  & (\3035(2374)  & (\3156(2706)  & (\4386(2698)  & \89(48) ))),
  \1175(3403)  = \1174(3290)  | \1173(3357) ,
  \2824(3611)  = ~\2823(3576)  | ~\2822(3591) ,
  \6017(346)  = \3719(239) ,
  \380(3086)  = \2571(3018)  & \2561(2925) ,
  \4474(759)  = \4451(732)  & \3707(243) ,
  \3214(1571)  = ~\6566(1414)  | ~\6559(944) ,
  \3274(2999)  = \3466(2558)  & \2537(2915) ,
  \6883(439)  = ~\6877(326) ,
  \7192(2278)  = \3932(1975) ,
  \3150(3241)  = ~\3149(3182)  | ~\3136(2475) ,
  \385(3151)  = \[68] ,
  \1940(2032)  = \1805(1806)  & (\1841(883)  & (\1795(1804)  & \1822(1811) )),
  \7451(3123)  = ~\7443(3061) ,
  \1607(1171)  = ~\5431(481)  | ~\5428(963) ,
  \5186(398)  = \1198(299) ,
  \7461(3125)  = ~\7453(3062) ,
  \991(3405)  = \980(3210)  & (\933(2683)  & \971(3356) ),
  \3666(698)  = \3642(579)  & \70(31) ,
  \6610(1266)  = \2198(974) ,
  \907(1028)  = \784(559)  & \765(774) ,
  \5455(475)  = ~\5449(359) ,
  \3092(1888)  = ~\6478(1604)  | ~\6471(1307) ,
  \2701(1995)  = ~\2700(1799)  | ~\2699(1505) ,
  \1935(2004)  = \1795(1804)  & (\1822(1811)  & (\1850(1812)  & \1805(1806) )),
  \1136(3174)  = \1038(1843)  & (\1074(1846)  & (\1055(1875)  & (\1093(1853)  & \3271(3101) ))),
  \6437(1187)  = ~\6431(914) ,
  \373(2994)  = \[56] ,
  \4743(3282)  = ~\4737(3220) ,
  \5102(2481)  = ~\948(2130)  & (~\947(2113)  & ~\845(980) ),
  \616(729)  = \587(402)  | \594(572) ,
  \1993(2659)  = ~\5840(2386)  | ~\5833(2393) ,
  \3971(1124)  = \2186(989)  & \4402(223) ,
  \3194(1617)  = ~\6542(1410)  | ~\6535(984) ,
  \5679(2951)  = ~\5678(2832)  | ~\5677(2676) ,
  \2972(1515)  = ~\6390(1424)  | ~\6383(880) ,
  \6917(335)  = \4396(225) ,
  \2436(1993)  = ~\2435(1797)  | ~\2434(1503) ,
  \1950(2047)  = \1903(1826)  & (\1859(1818)  & (\1885(1825)  & (\1921(1832)  & \1869(1819) ))),
  \3549(1696)  = ~\6772(1363)  | ~\6765(1365) ,
  \249(3418)  = \[72] ,
  \2554(3085)  = ~\2553(3012) ,
  \3755(412)  = \1535(302) ,
  \5148(3487)  = ~\5146(2452)  | ~\5139(3470) ,
  \1192(251)  = ~\2256(184) ,
  \6961(3457)  = ~\6955(3423) ,
  \3235(2435)  = \3234(2137)  | (\3233(2119)  | (\3232(2169)  | (\3231(2109)  | \3183(926) ))),
  \6318(2632)  = ~\6314(2346) ,
  \7479(890)  = \4698(766) ,
  \5940(2310)  = \2343(1982) ,
  \4344(2188)  = ~\4343(1658)  | ~\4342(1936) ,
  \7617(2506)  = ~\7611(2193) ,
  \268(3028)  = \997(2432)  & (\1788(2375)  & (\4089(2553)  & \2854(2916) )),
  \2299(782)  = \2279(739)  & \238(161) ,
  \318(3283)  = ~\4752(2425)  | ~\4745(3222) ,
  \6128(2611)  = ~\2766(2340)  & (~\2765(2324)  & ~\2612(1131) ),
  \2764(2319)  = \2600(1984)  & (\2618(1985)  & \2734(1987) ),
  \3474(2998)  = ~\3473(2759)  | ~\3472(2901) ,
  \2504(2334)  = \2354(1983)  & (\2372(1986)  & \2391(1134) ),
  \5511(3503)  = ~\5505(3480) ,
  \6935(3077)  = ~\6934(3003)  | ~\6933(2908) ,
  \4666(687)  = \4647(580)  & \82(41) ,
  \5213(672)  = ~\5207(549) ,
  \5424(1437)  = ~\5420(1082) ,
  \359(3426)  = \[96] ,
  \5009(3225)  = ~\5007(1201)  | ~\5000(3169) ,
  \2804(2327)  = \2618(1985)  & \2734(1987) ,
  \4076(3670)  = ~\7117(3661)  | ~\7114(2272) ,
  \6328(2642)  = ~\6324(2359) ,
  \311(3349)  = ~\4735(3280)  | ~\4732(2051) ,
  \2754(2314)  = \2612(1131)  & \2589(1981) ,
  \6740(1265)  = \2198(974) ,
  \3026(2020)  = \2977(879)  & (\2956(1802)  & \2965(1805) ),
  \763(723)  = ~\4879(495)  | ~\4876(401) ,
  \5314(1415)  = ~\5312(1061)  | ~\5305(845) ,
  \6762(1689)  = ~\6758(1351) ,
  \4966(1198)  = ~\4962(919) ,
  \2883(314)  = ~\2207(272)  | ~\4528(206) ,
  \7345(2154)  = ~\7292(1881)  | ~\7291(1868) ,
  \4889(378)  = \1482(281) ,
  \5173(3469)  = ~\5167(3446) ,
  \6397(1167)  = ~\6391(891) ,
  \5631(3525)  = ~\5630(3482)  | ~\5629(3505) ,
  \3468(2898)  = \3467(2760)  | \3437(2551) ,
  \2002(2947)  = ~\2001(2825) ,
  \4203(1923)  = ~\4202(1362)  | ~\4201(1695) ,
  \5368(2541)  = ~\5366(2217)  | ~\5359(1957) ,
  \6308(2647)  = ~\6304(2370) ,
  \1230(2221)  = ~\1226(1959) ,
  \2905(426)  = \1207(307) ,
  \1324(2461)  = \1304(2147)  & (\1267(2144)  & \1276(2145) ),
  \6106(3518)  = ~\6104(2605)  | ~\6097(3498) ,
  \1771(3137)  = ~\1766(3073) ,
  \5597(3043)  = ~\5591(2952) ,
  \4976(829)  = ~\4970(718) ,
  \3379(1480)  = ~\6621(444)  | ~\6618(1303) ,
  \6594(1375)  = \3821(1034) ,
  \4360(2699)  = ~\4356(2466) ,
  \4143(744)  = \4114(735)  & \4429(213) ,
  \825(1279)  = ~\4903(671)  | ~\4900(1093) ,
  \1138(2134)  = \1102(940)  & (\1055(1875)  & \1074(1846) ),
  \5214(1449)  = ~\5210(1094) ,
  \5904(1623)  = ~\5900(1288) ,
  \6575(320)  = \4434(211) ,
  \1128(2132)  = \1038(1843)  & (\1102(940)  & (\1026(1842)  & (\1055(1875)  & \1074(1846) ))),
  \6340(2539)  = ~\7359(2215)  | ~\7356(1955) ,
  \7237(1701)  = ~\7235(1381)  | ~\7232(1033) ,
  \4132(707)  = \4094(584)  & \59(22) ,
  \2152(660)  = \2117(577)  & \121(62) ,
  \4381(2964)  = ~\4360(2699)  | ~\4368(2855) ,
  \1929(910)  = \1399(820)  & \2213(268) ,
  \6074(2793)  = ~\6070(2612) ,
  \7432(1724)  = ~\7428(1404) ,
  \5919(461)  = ~\5913(348) ,
  \2051(804)  = \2026(730)  & \201(124) ,
  \5117(3113)  = ~\5115(3052)  | ~\5112(2687) ,
  \6670(2563)  = ~\6666(2232) ,
  \5474(2948)  = ~\5472(2822)  | ~\5465(885) ,
  \4570(1896)  = ~\7529(1661)  | ~\7526(1320) ,
  \2837(3682)  = ~\6249(3673)  | ~\6246(2351) ,
  \5980(2330)  = \2372(1986) ,
  \6096(3460)  = ~\6094(2620)  | ~\6087(3435) ,
  \6407(903)  = \4692(768) ,
  \4042(2289)  = \3971(1124)  & \3932(1975) ,
  \292(392)  = \[51] ,
  \4638(2723)  = \4618(2496)  & (\4581(2500)  & \4590(2499) ),
  \5540(2660)  = ~\5536(2387) ,
  \3703(245)  = ~\3701(186) ,
  \1590(882)  = \737(854)  & \2241(257) ,
  \3517(2120)  = ~\3513(1848) ,
  \4647(580)  = ~\4640(409) ,
  \7033(3548)  = ~\7032(3511)  | ~\7031(3530) ,
  \3082(2179)  = ~\3081(1641)  | ~\3080(1920) ,
  \3267(3035)  = \1974(2382)  & (\3466(2558)  & \2537(2915) ),
  \7120(3608)  = ~\7196(2591)  | ~\7189(3588) ,
  \7110(3609)  = ~\7108(2592)  | ~\7101(3589) ,
  \2151(809)  = \2124(731)  & \194(117) ,
  \6864(1352)  = \3833(1016) ,
  \6134(3146)  = ~\6132(2792)  | ~\6125(3087) ,
  \3107(1305)  = \2171(992)  & \4157(1010) ,
  \6861(321)  = \4434(211) ,
  \361(3324)  = ~\4816(2586)  | ~\4809(3253) ,
  \4710(762)  = \4685(465)  | \4684(669) ,
  \1074(1846)  = ~\1073(1565)  | ~\1072(1214) ,
  \4631(2866)  = \4613(2728)  & (\4567(2501)  & \4554(1900) ),
  \4442(290)  = \186(109)  & (\185(108)  & (\182(105)  & \183(106) )),
  \2629(1133)  = \2099(970)  & \3739(233) ,
  \6582(1688)  = ~\6578(1350) ,
  \3571(2096)  = \3522(1839) ,
  \971(3356)  = ~\5009(3225)  | ~\5008(3289) ,
  \1331(3188)  = ~\1330(3067)  | ~\1329(3132) ,
  \2052(658)  = \2019(576)  & \124(63) ,
  \2341(1488)  = ~\5871(450)  | ~\5868(1291) ,
  \2560(2800)  = ~\5984(2622)  | ~\5977(1493) ,
  \4544(2062)  = ~\4540(1822) ,
  \5571(3523)  = ~\5569(3504)  | ~\5566(2000) ,
  \5315(965)  = \1399(820) ,
  \4968(3224)  = ~\4966(1198)  | ~\4959(3170) ,
  \6143(3383)  = ~\6141(3331)  | ~\6138(2342) ,
  \4094(584)  = \1530(411) ,
  \4417(217)  = ~\4415(200) ,
  \303(3271)  = \2002(2947)  & \2008(3214) ,
  \1991(3031)  = ~\1990(2943) ,
  \1117(1193)  = \1116(1031)  | \1115(371) ,
  \7157(3322)  = ~\7155(3255)  | ~\7152(2584) ,
  \1387(812)  = \1368(520)  | \1367(650) ,
  \258(3122)  = \[58] ,
  \2579(3011)  = \2564(2929)  & \2577(2920) ,
  \4783(3299)  = ~\4777(3235) ,
  \6729(1301)  = \2192(991) ,
  \406(388)  = \[43] ,
  \6543(937)  = \3670(778) ,
  \3801(824)  = \3782(553)  | \3781(621) ,
  \1025(1560)  = ~\5198(1461)  | ~\5191(376) ,
  \5792(1243)  = ~\5788(964) ,
  \2812(2995)  = ~\2809(2893) ,
  \6350(2514)  = ~\7343(2191)  | ~\7340(1931) ,
  \5889(343)  = \3731(235) ,
  \5639(3564)  = ~\5637(3542)  | ~\5634(2045) ,
  \4639(2973)  = ~\4638(2723)  & ~\4637(2864) ,
  \1329(3132)  = ~\5383(3066)  | ~\5380(1736) ,
  \5059(3507)  = ~\5057(3489)  | ~\5054(2121) ,
  \5579(3559)  = ~\5573(3538) ,
  \4477(693)  = \4444(582)  & \76(35) ,
  \3910(1775)  = ~\6892(1603)  | ~\6885(329) ,
  \1710(2028)  = \1556(1807)  & (\1590(882)  & \1573(1810) ),
  \7200(3699)  = \4088(3688)  | \4087(3695) ,
  \1133(2115)  = \1038(1843)  & (\1086(935)  & \1055(1875) ),
  \4860(2358)  = \2436(1993) ,
  \3131(2733)  = \3130(2513)  | (\3129(2516)  | (\3128(2509)  | \3059(1330) )),
  \1155(2201)  = ~\1154(1928) ,
  \2537(2915)  = \2536(2789)  | \2495(2601) ,
  \4912(1451)  = ~\4908(1096) ,
  \1249(1952)  = ~\1248(1730)  | ~\1247(1732) ,
  \5304(1407)  = ~\5300(1052) ,
  \5250(1101)  = ~\4525(862) ,
  \2919(518)  = \2892(416)  & \209(132) ,
  \3015(912)  = \1383(815)  & \4686(770) ,
  \701(541)  = \678(414)  & \157(80) ,
  \1291(2543)  = ~\1288(2219) ,
  \3156(2706)  = \3136(2475)  & \3123(2497) ,
  \4081(3679)  = ~\4080(3658)  | ~\4079(3669) ,
  \6920(1276)  = \2179(977) ,
  \3652(668)  = \3629(578)  & \111(56) ,
  \1323(2695)  = \1307(2463)  & (\1276(2145)  & \1263(1857) ),
  \4012(2255)  = \3856(1966)  & (\3891(1114)  & \3874(1968) ),
  \5433(364)  = \2226(264) ,
  \6033(350)  = \3707(243) ,
  \6815(2504)  = ~\6809(2190) ,
  \2654(1795)  = ~\6024(1718)  | ~\6017(346) ,
  \7487(881)  = \4704(764) ,
  \3660(608)  = \3642(579)  & \1455(166) ,
  \2924(610)  = \2923(513)  | \2899(590) ,
  \2833(317)  = ~\2828(208) ,
  \2285(616)  = \2266(587)  & \208(131) ,
  \3(312)  = \1(0) ,
  \536(222)  = \4405(198) ,
  \4949(2954)  = ~\4948(2680)  | ~\4947(2836) ,
  \4037(2298)  = \3911(1974)  & (\3979(1126)  & (\3932(1975)  & \3957(1977) )),
  \3164(2980)  = \3163(2861)  | \3131(2733) ,
  \2399(1792)  = ~\5896(1588)  | ~\5889(343) ,
  \3891(1114)  = \3821(1034)  & \4422(215) ,
  \6546(1057)  = \633(843) ,
  \4027(2299)  = \3911(1974)  & (\3979(1126)  & (\3899(1971)  & (\3932(1975)  & \3957(1977) ))),
  \1325(2848)  = ~\1324(2461)  & ~\1323(2695) ,
  \4154(996)  = \4129(691)  | \4128(749) ,
  \1257(1737)  = ~\5304(1407)  | ~\5297(1062) ,
  \6784(1396)  = \2335(1044) ,
  \5729(3582)  = ~\5728(3540)  | ~\5727(3563) ,
  \615(529)  = \587(402)  & \170(93) ,
  \1247(1732)  = ~\5295(1409)  | ~\5292(1056) ,
  \6211(3491)  = ~\6209(3464)  | ~\6206(2747) ,
  \522(226)  = \4394(196) ,
  \1545(1509)  = ~\5400(1439)  | ~\5393(352) ,
  \6525(1207)  = ~\6519(928) ,
  \3522(1839)  = ~\3521(1557)  | ~\3520(1564) ,
  \5644(2064)  = \1630(1824) ,
  \316(3397)  = \[79] ,
  \3540(2491)  = ~\3536(2174) ,
  \6329(3641)  = \2847(3624)  | (\2846(3623)  | (\2845(3626)  | \2844(3625) )),
  \575(309)  = ~\5(1) ,
  \7521(1652)  = ~\7515(1317) ,
  \1412(818)  = \1380(539)  | \1379(645) ,
  \2861(3189)  = ~\2860(3068)  | ~\2859(3133) ,
  \6690(780)  = \3649(511)  | \3648(665) ,
  \581(421)  = \1206(306) ,
  \7079(3459)  = ~\7077(3428)  | ~\7074(2306) ,
  \2557(2928)  = ~\2556(2801)  | ~\2555(2627) ,
  \486(258)  = \2239(181) ,
  \4618(2496)  = \4595(2178) ,
  \2130(593)  = \1507(418) ,
  \1791(3701)  = ~\5743(3647)  | ~\5740(3694) ,
  \5258(1097)  = \2938(860) ,
  \641(841)  = \581(421)  & \622(634) ,
  \6677(1474)  = ~\6671(1116) ,
  \4978(1926)  = ~\4976(829)  | ~\4973(1548) ,
  \4508(1013)  = \4487(710)  | \4486(753) ,
  \6301(3490)  = ~\6300(3453)  | ~\6299(3472) ,
  \5218(1095)  = \2938(860) ,
  \5149(3528)  = ~\5148(3487)  | ~\5147(3508) ,
  \7271(1620)  = ~\7265(1285) ,
  \2577(2920)  = ~\2491(2608)  | ~\2499(2782) ,
  \7188(3550)  = ~\7186(2580)  | ~\7179(3533) ,
  \5041(3360)  = ~\5040(3232)  | ~\5039(3296) ,
  \293(3285)  = ~\4719(3192)  | ~\4716(2094) ,
  \400(297)  = ~\57(20) ,
  \6311(3537)  = ~\6310(3500)  | ~\6309(3522) ,
  \3856(1966)  = ~\3855(1765)  | ~\3854(1466) ,
  \7019(3456)  = ~\7013(3422) ,
  \1366(528)  = \1336(405)  & \171(94) ,
  \5848(2385)  = ~\5844(2007) ,
  \2419(1796)  = ~\5912(1717)  | ~\5905(347) ,
  \343(3258)  = ~\4800(2598)  | ~\4793(3203) ,
  \5318(816)  = \1374(537)  | \1373(648) ,
  \6835(3049)  = ~\6829(2957) ,
  \6999(3140)  = ~\6993(3076) ,
  \7515(1317)  = \4493(998) ,
  \4315(1877)  = ~\7391(1662)  | ~\7388(1283) ,
  \4880(566)  = ~\4876(401) ,
  \1555(1514)  = ~\5408(1442)  | ~\5401(355) ,
  \7255(1364)  = ~\7249(1024) ,
  \3232(2169)  = \3200(982)  & (\3176(1840)  & \3186(1845) ),
  \2294(571)  = \2259(413)  & \23(6) ,
  \1161(3229)  = \1160(3173)  | \1129(2434) ,
  \3595(2688)  = \3574(2438)  & (\3513(1848)  & \3508(2138) ),
  \3122(2158)  = ~\3121(1894)  | ~\3120(1871) ,
  \1609(1820)  = ~\1608(1530)  | ~\1607(1171) ,
  \2491(2608)  = ~\2487(2312) ,
  \4235(1855)  = ~\4234(1577)  | ~\4233(1576) ,
  \2842(3681)  = ~\2841(3662)  | ~\2840(3671) ,
  \4375(2521)  = \4327(2186)  & (\4349(1400)  & (\4317(2170)  & (\4336(2185)  & \4344(2188) ))),
  \4962(919)  = \765(774) ,
  \1738(2067)  = \1609(1820)  & (\1669(904)  & \1630(1824) ),
  \2545(2787)  = ~\5952(2607)  | ~\5945(2609) ,
  \3785(623)  = \3762(586)  & \191(114) ,
  \6161(3520)  = ~\6155(3499) ,
  \5664(2052)  = \1609(1820) ,
  \436(286)  = \1462(168) ,
  \6280(3096)  = ~\6278(2940)  | ~\6271(3064) ,
  \5654(2054)  = \1609(1820) ,
  \1068(981)  = \2942(859)  & \1477(394) ,
  \6239(3633)  = ~\6233(3613) ,
  \6565(1223)  = ~\6559(944) ,
  \6466(1019)  = \3801(824) ,
  \3793(796)  = \3775(740)  & \222(145) ,
  \2335(1044)  = \2304(728)  | \2303(784) ,
  \7249(1024)  = \2305(826) ,
  \4669(490)  = \4640(409)  & \2213(268) ,
  \2777(2357)  = \2693(1143)  & (\2643(1990)  & \2655(1991) ),
  \4793(3203)  = \2580(3145) ,
  \4140(745)  = \4114(735)  & \4422(215) ,
  \243(3032)  = \1146(2431)  & (\1974(2382)  & \3468(2898) ),
  \1779(3648)  = ~\5668(2416)  | ~\5661(3637) ,
  \3700(247)  = ~\3698(185) ,
  \5279(1458)  = ~\5277(1102)  | ~\5274(864) ,
  \7581(1677)  = ~\7575(1338) ,
  \4613(2728)  = ~\4610(2502) ,
  \7575(1338)  = \4169(1009) ,
  \6345(3054)  = ~\6337(2961) ,
  \5269(1459)  = ~\5263(1104) ,
  \5326(956)  = \1406(817) ,
  \4444(582)  = \1530(411) ,
  \4482(755)  = \4464(733)  & \3731(235) ,
  \1743(2070)  = \1669(904)  & \1630(1824) ,
  \2979(886)  = \715(851)  & \4701(765) ,
  \7235(1381)  = ~\7229(1037) ,
  \4267(2143)  = \4244(1856) ,
  \7348(2148)  = ~\7282(1865)  | ~\7281(1860) ,
  \3017(1524)  = ~\6430(1425)  | ~\6423(888) ,
  \6025(349)  = \3713(241) ,
  \366(3381)  = ~\4831(3329)  | ~\4828(2293) ,
  \3102(2177)  = ~\3101(1907)  | ~\3100(1886) ,
  \3258(2546)  = \3235(2435)  & \3216(1462) ,
  \6279(3155)  = ~\6277(3130)  | ~\6274(2812) ,
  \3163(2861)  = \3143(2738)  & \3123(2497) ,
  \4552(1664)  = ~\7513(1325)  | ~\7510(1003) ,
  \7591(1671)  = ~\7585(1334) ,
  \3673(821)  = \3655(550)  | \3654(682) ,
  \7585(1334)  = \4175(1007) ,
  \6891(442)  = ~\6885(329) ,
  \6110(2318)  = \2600(1984) ,
  \7169(3476)  = ~\7168(3432)  | ~\7167(3458) ,
  \2312(836)  = \2292(570)  | \2291(618) ,
  \6892(1603)  = ~\6888(1267) ,
  \4539(1533)  = ~\7478(1181)  | ~\7471(902) ,
  \3613(3108)  = ~\6835(3049)  | ~\6832(1546) ,
  \7436(2394)  = ~\7601(1997)  | ~\7598(1809) ,
  \3502(1573)  = ~\6693(1222)  | ~\6690(780) ,
  \7602(2021)  = ~\7598(1809) ,
  \1757(3594)  = ~\1756(3561)  | ~\1755(3580) ,
  \3028(2372)  = \3027(2040)  | (\3026(2020)  | (\3025(2005)  | \2962(867) )),
  \5991(449)  = ~\5985(336) ,
  \7570(1308)  = \4160(993) ,
  \5812(966)  = \1399(820) ,
  \6876(1706)  = ~\6872(1377) ,
  \5624(2076)  = \1655(1827) ,
  \4577(2183)  = ~\4576(1650)  | ~\4575(1909) ,
  \2487(2312)  = \2343(1982)  & (\2372(1986)  & (\2400(1988)  & \2354(1983) )),
  \1920(1544)  = ~\5816(1245)  | ~\5809(369) ,
  \6221(3536)  = ~\6219(3529)  | ~\6216(2369) ,
  \3140(2494)  = \3107(1305)  & (\3082(2179)  & \3093(2156) ),
  \6718(921)  = ~\6714(775) ,
  \6125(3087)  = ~\6124(3014)  | ~\6123(2926) ,
  \396(2941)  = ~\4872(2649)  | ~\4865(2877) ,
  \3031(2061)  = \3006(901)  & (\2982(1816)  & \2992(1821) ),
  \3052(2192)  = ~\3051(1669)  | ~\3050(1903) ,
  \4052(2292)  = \3957(1977)  & \3997(1980) ,
  \6490(1299)  = \2167(990) ,
  \7132(2589)  = ~\4046(2303)  & (~\4045(2288)  & ~\3949(1122) ),
  \416(3368)  = \[71] ,
  \7152(2584)  = ~\4041(2300)  & (~\4040(2285)  & (~\4039(2275)  & ~\3926(1120) )),
  \3739(233)  = ~\3737(192) ,
  \2157(792)  = \2137(738)  & \226(149) ,
  \6151(3462)  = ~\6145(3434) ,
  \7400(1398)  = ~\7396(1045) ,
  \3062(2194)  = ~\3061(1672)  | ~\3060(1919) ,
  \827(1874)  = ~\826(1614)  | ~\825(1279) ,
  \3586(2704)  = ~\3583(2472) ,
  \6189(3187)  = ~\6183(3131) ,
  \7360(2216)  = ~\7356(1955) ,
  \1869(1819)  = ~\1868(1529)  | ~\1867(1170) ,
  \1859(1818)  = ~\1858(1528)  | ~\1857(1169) ,
  \4529(1545)  = ~\7469(1186)  | ~\7466(771) ,
  \6944(3139)  = ~\6942(2764)  | ~\6935(3077) ,
  \4668(701)  = \4647(580)  & \65(28) ,
  \3169(597)  = ~\6518(558)  | ~\6511(429) ,
  \7068(2775)  = ~\7064(2585) ,
  \7048(2777)  = ~\7044(2590) ,
  \7364(1292)  = \2081(988) ,
  \2512(2354)  = \2448(1142)  & (\2409(1989)  & \2420(1992) ),
  \1166(3292)  = ~\1161(3229) ,
  \3725(237)  = ~\3723(190) ,
  \5081(3640)  = ~\5080(3603)  | ~\5079(3622) ,
  \6382(1421)  = ~\6378(1066) ,
  \7312(952)  = \1395(814) ,
  \6727(1611)  = ~\6721(1274) ,
  \1173(3357)  = \1166(3292)  & \1019(923) ,
  \5960(2614)  = ~\5956(2316) ,
  \3380(1777)  = ~\6622(1636)  | ~\6615(331) ,
  \2828(208)  = \4526(205) ,
  \5109(2959)  = ~\5108(2843)  | ~\5107(2690) ,
  \4841(2804)  = \2522(2550)  | (\2520(2522)  | (\2519(2361)  | (\2518(2353)  | \2431(1140) ))),
  \6366(2963)  = ~\6362(2849) ,
  \5039(3296)  = ~\5037(3236)  | ~\5034(2444) ,
  \3220(1761)  = ~\3216(1462) ,
  \4314(1248)  = \2069(968)  & \4502(1015) ,
  \378(3091)  = \2550(3013)  & \2564(2929) ,
  \1733(2057)  = \1647(899)  & \1609(1820) ,
  \1723(2058)  = \1647(899)  & (\1598(1817)  & \1609(1820) ),
  \6981(3568)  = ~\6975(3549) ,
  \6352(2734)  = ~\6351(2505)  | ~\6350(2514) ,
  \5475(3038)  = ~\5474(2948)  | ~\5473(2826) ,
  \2954(1740)  = ~\6373(1147)  | ~\6370(1065) ,
  \4916(400)  = \1198(299) ,
  \5463(489)  = ~\5457(368) ,
  \5611(3348)  = ~\5610(3216)  | ~\5609(3277) ,
  \388(3093)  = \[61] ,
  \5614(2091)  = \1695(1829) ,
  \4151(997)  = \4126(692)  | \4125(750) ,
  \2589(1981)  = ~\2588(1783)  | ~\2587(1487) ,
  \5369(2989)  = ~\1310(2887)  | ~\1313(2886) ,
  \5091(3639)  = ~\5090(3602)  | ~\5089(3621) ,
  \4352(2149)  = ~\4351(1917)  | ~\4350(1861) ,
  \7146(2911)  = ~\7142(2778) ,
  \7061(3199)  = ~\7060(3079)  | ~\7059(3143) ,
  \7340(1931)  = ~\7238(1708)  | ~\7237(1701) ,
  \7229(1037)  = \3807(834) ,
  \5784(1436)  = ~\5780(1081) ,
  \6787(1621)  = ~\6781(1286) ,
  \7001(3193)  = ~\6999(3140)  | ~\6996(2561) ,
  \4540(1822)  = ~\4539(1533)  | ~\4538(1540) ,
  \4515(3099)  = ~\7441(3039)  | ~\7438(2650) ,
  \1985(2817)  = ~\5823(2657)  | ~\5820(2002) ,
  \3007(1575)  = ~\6421(1180)  | ~\6418(947) ,
  \2304(728)  = \2272(594)  & \23(6) ,
  \4059(3604)  = ~\4058(3569)  | ~\4057(3586) ,
  \7148(3078)  = ~\7146(2911)  | ~\7139(3006) ,
  \7304(948)  = \1387(812) ,
  \6418(947)  = \1387(812) ,
  \4674(684)  = \4647(580)  & \85(44) ,
  \3525(1873)  = ~\6727(1611)  | ~\6724(979) ,
  \1995(2819)  = ~\5847(2663)  | ~\5844(2007) ,
  \5551(3344)  = ~\5549(3268)  | ~\5546(2038) ,
  \5769(358)  = \2241(257) ,
  \351(3372)  = \3497(3319)  & \3489(2906) ,
  \606(403)  = \1512(300) ,
  \5927(464)  = ~\5921(351) ,
  \5254(1456)  = ~\5250(1101) ,
  \251(3365)  = \3131(2733)  & \3152(3305) ,
  \6423(888)  = \4701(765) ,
  \6710(1213)  = ~\6706(933) ,
  \558(244)  = \3705(187) ,
  \1953(2050)  = \1880(895)  & \1859(1818) ,
  \2065(985)  = \2046(673)  | \2045(801) ,
  \6583(322)  = \4429(213) ,
  \7404(1042)  = \2312(836) ,
  \289(383)  = \[50] ,
  \5687(3106)  = ~\5685(3042)  | ~\5682(2674) ,
  \5191(376)  = \1488(279) ,
  \2792(2355)  = \2693(1143)  & \2655(1991) ,
  \7211(1609)  = ~\7205(1273) ,
  \6080(2343)  = \2734(1987) ,
  \241(2837)  = \1151(2681)  | \1117(1193) ,
  \5494(3273)  = ~\5492(2402)  | ~\5485(3213) ,
  \5945(2609)  = ~\2504(2334)  & (~\2503(2323)  & ~\2366(1130) ),
  \4518(3183)  = ~\7451(3123)  | ~\7448(2862) ,
  \5472(2822)  = ~\5468(2665) ,
  \2179(977)  = \2156(662)  | \2155(800) ,
  \2962(867)  = \727(848)  & \4710(762) ,
  \301(3388)  = \[88] ,
  \6077(3261)  = ~\6076(3147)  | ~\6075(3205) ,
  \3535(1885)  = ~\6736(1629)  | ~\6729(1301) ,
  \2918(736)  = \2892(416)  | \2899(590) ,
  \5621(3468)  = ~\5620(3400)  | ~\5619(3443) ,
  \3545(2155)  = ~\3544(1922)  | ~\3543(1869) ,
  \271(3354)  = \1166(3292)  & \1117(1193) ,
  \4572(2187)  = ~\4571(1898)  | ~\4570(1896) ,
  \4193(2493)  = ~\4189(2176) ,
  \5561(3466)  = ~\5559(3440)  | ~\5556(2024) ,
  \3212(1367)  = ~\3211(827)  | ~\3210(1026) ,
  \3222(1366)  = \3173(717)  & \3170(866) ,
  \1270(1583)  = ~\5329(1238)  | ~\5326(956) ,
  \1948(2027)  = \1822(1811)  & \1850(1812) ,
  \4451(732)  = ~\4444(582) ,
  \826(1614)  = ~\4904(1448)  | ~\4897(548) ,
  \2060(655)  = \2032(592)  & \127(64) ,
  \1784(3617)  = \1766(3073)  & (\1751(2828)  & \1762(3595) ),
  \3242(3098)  = \3241(2859)  | (\3240(3026)  | (\3239(3025)  | \3046(2813) )),
  \3243(3171)  = ~\3242(3098)  | ~\3228(2097) ,
  \1178(261)  = ~\2236(180) ,
  \6415(907)  = \4689(769) ,
  \6086(3334)  = ~\6084(2626)  | ~\6077(3261) ,
  \5323(959)  = \1412(818) ,
  \2492(2313)  = \2366(1130)  & \2343(1982) ,
  \3979(1126)  = \2179(977)  & \4396(225) ,
  \1475(295)  = \106(53) ,
  \3949(1122)  = \2192(991)  & \4407(221) ,
  \1762(3595)  = ~\1761(3562)  | ~\1760(3581) ,
  \3897(1475)  = ~\6883(439)  | ~\6880(1361) ,
  \4439(209)  = ~\4437(204) ,
  \7239(1005)  = \3813(822) ,
  \7315(1427)  = ~\7309(1072) ,
  \2279(739)  = ~\2272(594) ,
  \469(3452)  = \1172(3419) ,
  \2417(1138)  = \2085(986)  & \3725(237) ,
  \987(3667)  = ~\5097(3654)  | ~\5094(2106) ,
  \4948(2680)  = ~\4946(1837)  | ~\4939(2512) ,
  \6666(2232)  = \3295(1965) ,
  \6728(1278)  = ~\6724(979) ,
  \7012(3315)  = ~\7010(2575)  | ~\7003(3247) ,
  \6827(2700)  = ~\6825(2469)  | ~\6822(2150) ,
  \4768(2442)  = ~\4764(2102) ,
  \4523(3246)  = ~\4522(3128)  | ~\4521(3186) ,
  \2734(1987)  = ~\2733(1791)  | ~\2732(1496) ,
  \4350(1861)  = ~\7423(1687)  | ~\7420(1249) ,
  \790(1208)  = ~\4887(500)  | ~\4884(1105) ,
  \1395(814)  = \1372(522)  | \1371(652) ,
  \6121(1790)  = ~\6115(1494) ,
  \6438(1233)  = ~\6434(954) ,
  \1957(2411)  = \1956(2087)  | (\1955(2073)  | (\1954(2060)  | (\1953(2050)  | \1866(893) ))),
  \2320(1025)  = \2298(716)  | \2297(790) ,
  \4728(2412)  = ~\4724(2048) ,
  \7279(1595)  = ~\7273(1258) ,
  \544(230)  = \3749(194) ,
  \6090(2328)  = \2618(1985) ,
  \2724(1722)  = \4389(1405)  & \3682(839) ,
  \331(3364)  = ~\4783(3299)  | ~\4780(2168) ,
  \6141(3331)  = ~\6135(3260) ,
  \5330(1235)  = ~\5326(956) ,
  \5897(344)  = \3725(237) ,
  \4224(1574)  = ~\7299(1232)  | ~\7296(811) ,
  \6181(2987)  = ~\6179(1946)  | ~\6176(2809) ,
  \5069(3566)  = ~\5067(3546)  | ~\5064(2099) ,
  \3128(2509)  = \3068(1353)  & \3052(2192) ,
  \1445(2895)  = \1788(2375)  & (\4089(2553)  & (\2852(2785)  & \4526(205) )),
  \3898(1772)  = ~\6884(1694)  | ~\6877(326) ,
  \5844(2007)  = \1805(1806) ,
  \5629(3505)  = ~\5627(3485)  | ~\5624(2076) ,
  \1964(3162)  = \1869(1819)  & (\1903(1826)  & (\1885(1825)  & (\1921(1832)  & \3279(3072) ))),
  \5440(1240)  = ~\5436(961) ,
  \1500(296)  = ~\106(53) ,
  \6991(2907)  = ~\6989(1769)  | ~\6986(2769) ,
  \6971(3513)  = ~\6965(3492) ,
  \7224(1270)  = \2175(975) ,
  \3045(2651)  = \3034(2403)  & \3022(1998) ,
  \2801(2645)  = \2800(2530)  | \2715(1145) ,
  \5948(2311)  = \2343(1982) ,
  \2791(2637)  = \2701(1995)  & (\2655(1991)  & (\2676(1994)  & \2742(2533) )),
  \6231(3593)  = ~\6229(3579)  | ~\6226(2347) ,
  \2982(1816)  = ~\2981(1526)  | ~\2980(1748) ,
  \6942(2764)  = ~\6938(2562) ,
  \3655(550)  = \3622(407)  & \1500(296) ,
  \3911(1974)  = ~\3910(1775)  | ~\3909(1478) ,
  \494(267)  = \2218(177) ,
  \2932(614)  = \2931(517)  | \2914(591) ,
  \4207(2198)  = ~\4203(1923) ,
  \6888(1267)  = \2198(974) ,
  \6454(1354)  = ~\6450(1017) ,
  \6287(3264)  = ~\6281(3209) ,
  \719(850)  = \650(423)  & \696(628) ,
  \4138(689)  = \4107(585)  & \80(39) ,
  \4234(1577)  = ~\7308(1227)  | ~\7301(949) ,
  \623(533)  = \606(403)  & \166(89) ,
  \2771(2634)  = \2643(1990)  & (\2655(1991)  & (\2676(1994)  & (\2701(1995)  & \2742(2533) ))),
  \4210(1712)  = ~\7263(1393)  | ~\7260(1040) ,
  \6100(2309)  = \2589(1981) ,
  \2293(619)  = \2266(587)  & \205(128) ,
  \2927(515)  = \2909(417)  & \213(136) ,
  \4800(2598)  = ~\4796(2304) ,
  \7204(3706)  = ~\7200(3699) ,
  \6557(741)  = ~\6551(599) ,
  \2057(786)  = \2039(737)  & \234(157) ,
  \618(632)  = \617(530)  | \594(572) ,
  \7059(3143)  = ~\7057(3081)  | ~\7054(2779) ,
  \5999(452)  = ~\5993(339) ,
  \7443(3061)  = ~\4636(2976)  | ~\4639(2973) ,
  \4791(3301)  = ~\4785(3237) ,
  \6751(1705)  = ~\6745(1376) ,
  \1450(2996)  = \4089(2553)  & \2854(2916) ,
  \4271(2857)  = \4250(2709)  & (\4189(2176)  & \4184(2479) ),
  \3116(1271)  = \2163(976)  & \4151(997) ,
  \6321(3592)  = ~\6320(3556)  | ~\6319(3577) ,
  \1004(3708)  = ~\5174(3700)  | ~\5167(3446) ,
  \5205(502)  = ~\5199(377) ,
  \2856(3709)  = ~\6336(3704)  | ~\6329(3641) ,
  \704(639)  = \703(542)  | \685(588) ,
  \961(3291)  = ~\958(3228) ,
  \2160(679)  = \2130(593)  & \94(49) ,
  \376(3206)  = \[65] ,
  \349(3314)  = \3478(3001)  & \3491(3249) ,
  \4279(2982)  = ~\4278(2739)  & ~\4277(2876) ,
  \4064(3605)  = ~\4063(3570)  | ~\4062(3587) ,
  \1464(285)  = ~\1462(168) ,
  \5441(367)  = \2220(266) ,
  \5366(2217)  = ~\5362(1956) ,
  \7477(1174)  = ~\7471(902) ,
  \7453(3062)  = ~\4630(2977)  | ~\4633(2978) ,
  \6622(1636)  = ~\6618(1303) ,
  \6720(1189)  = ~\6718(921)  | ~\6711(772) ,
  \6605(440)  = ~\6599(327) ,
  \1990(2943)  = ~\1989(2654)  | ~\1988(2818) ,
  \4471(699)  = \4444(582)  & \69(30) ,
  \4753(3158)  = \3271(3101) ,
  \5569(3504)  = ~\5563(3481) ,
  \4724(2048)  = \1859(1818) ,
  \6916(1703)  = ~\6912(1374) ,
  \2847(3624)  = \2828(208)  & (\2816(3019)  & \2819(3610) ),
  \4980(2511)  = ~\4979(2200)  | ~\4978(1926) ,
  \3611(2718)  = \3591(2490)  & (\3554(2510)  & \3563(2517) ),
  \7566(1648)  = ~\7562(1314) ,
  \3612(2970)  = ~\3611(2718)  & ~\3610(2873) ,
  \3101(1907)  = ~\6486(1637)  | ~\6479(1339) ,
  \480(250)  = \2256(184) ,
  \939(2125)  = \805(1844)  & (\877(939)  & (\827(1874)  & \853(1849) )),
  \1371(652)  = \1343(575)  & \135(68) ,
  \7603(2196)  = ~\7550(1910)  | ~\7549(1913) ,
  \2992(1821)  = ~\2991(1531)  | ~\2990(1579) ,
  \530(216)  = \4420(201) ,
  \444(282)  = \1480(170) ,
  \4376(2714)  = \4375(2521)  | (\4374(2518)  | (\4373(2519)  | (\4372(2520)  | \4324(1284) ))),
  \299(3341)  = \2014(3274)  & \1998(3036) ,
  \5399(466)  = ~\5393(352) ,
  \4623(2420)  = \4598(2042)  & (\4531(1830)  & \4540(1822) ),
  \1718(2046)  = \1598(1817)  & (\1609(1820)  & (\1630(1824)  & (\1655(1827)  & \1695(1829) ))),
  \2866(3115)  = ~\6366(2963)  | ~\6357(3063) ,
  \1288(2219)  = \1235(1958) ,
  \6259(3663)  = ~\6253(3645) ,
  \4514(292)  = \230(153)  & (\218(141)  & (\152(75)  & \210(133) )),
  \3482(3075)  = ~\3481(3000) ,
  \949(2129)  = \877(939)  & \853(1849) ,
  \256(2991)  = \3249(2223)  & (\3035(2374)  & (\3156(2706)  & \4388(2971) )),
  \7301(949)  = \1391(813) ,
  \383(3089)  = \2571(3018)  & \2400(1988) ,
  \4101(734)  = ~\4094(584) ,
  \4955(3046)  = ~\4949(2954) ,
  \6817(2744)  = ~\6815(2504)  | ~\6812(2204) ,
  \2998(896)  = \1395(814)  & \4695(767) ,
  \3472(2901)  = ~\6653(2761)  | ~\6650(2228) ,
  \994(3407)  = \975(3157)  & (\965(2958)  & \967(3355) ),
  \727(848)  = \650(423)  & \700(630) ,
  \6829(2957)  = ~\3597(2841)  | ~\3600(2838) ,
  \3838(1004)  = \3800(700)  | \3799(799) ,
  \4868(2371)  = \2454(1996) ,
  \4820(2281)  = \3381(1976) ,
  \1943(2034)  = \1805(1806)  & (\1841(883)  & \1822(1811) ),
  \1374(537)  = \1350(415)  & \161(84) ,
  \4610(2502)  = \4572(2187) ,
  \5871(450)  = ~\5865(337) ,
  \4317(2170)  = ~\4316(1899)  | ~\4315(1877) ,
  \2014(3274)  = ~\2008(3214) ,
  \5542(3102)  = ~\5540(2660)  | ~\5533(3037) ,
  \2868(3308)  = \2867(3239)  & (\2864(3245)  & (\2861(3189)  & \1331(3188) )),
  \6426(1070)  = \715(851) ,
  \4091(2899)  = \4090(2757)  | \4010(2552) ,
  \3663(493)  = \3635(408)  & \1499(273) ,
  \3029(2043)  = \2982(1816)  & (\2992(1821)  & (\3001(1823)  & (\3009(1828)  & \3021(1831) ))),
  \6925(1115)  = ~\3821(1034)  & ~\4422(215) ,
  \6132(2792)  = ~\6128(2611) ,
  \4355(2207)  = ~\4354(1943)  | ~\4353(1720) ,
  \4927(508)  = ~\4921(381) ,
  \2547(3084)  = ~\2546(3010) ,
  \5833(2393)  = \1948(2027)  | (\1947(2035)  | \1834(878) ),
  \6434(954)  = \1383(815) ,
  \3457(2282)  = \3365(1973)  & (\3410(1123)  & \3381(1976) ),
  \5334(962)  = \1418(819) ,
  \5523(1158)  = \1590(882) ,
  \3872(1468)  = ~\6875(436)  | ~\6872(1377) ,
  \906(1554)  = ~\902(1199) ,
  \1787(3678)  = \1777(3675)  & \1766(3073) ,
  \5337(1435)  = ~\5331(1080) ,
  \1309(2545)  = \1284(2220)  & (\1217(1960)  & \1226(1959) ),
  \1996(2658)  = ~\5848(2385)  | ~\5841(2392) ,
  \5478(2388)  = \1711(2012)  | (\1710(2028)  | (\1709(2016)  | \1567(876) )),
  \4422(215)  = ~\4420(201) ,
  \4998(3111)  = ~\4996(3045)  | ~\4993(1203) ,
  \957(1836)  = ~\906(1554)  | ~\912(1550) ,
  \3248(3293)  = ~\3245(3230) ,
  \3987(1472)  = ~\6915(437)  | ~\6912(1374) ,
  \4010(2552)  = \4009(2256)  | (\4008(2242)  | (\4007(2231)  | \3853(1108) )),
  \5799(485)  = ~\5793(365) ,
  \1986(2653)  = ~\5824(2380)  | ~\5817(2384) ,
  \1334(3190)  = ~\1333(3069)  | ~\1332(3134) ,
  \6542(1410)  = ~\6538(1055) ,
  \5588(2672)  = ~\5584(2419) ,
  \4677(477)  = \4653(410)  & \2238(259) ,
  \1777(3675)  = ~\1776(3649)  | ~\1775(3666) ,
  \2767(2341)  = \2635(1135)  & \2618(1985) ,
  \5608(2670)  = ~\5604(2414) ,
  \1938(2006)  = \1816(875)  & \1795(1804) ,
  \5977(1493)  = \2391(1134) ,
  \2019(576)  = \1514(406) ,
  \4327(2186)  = ~\4326(1655)  | ~\4325(1941) ,
  \6447(1335)  = \4172(1008) ,
  \3616(3184)  = ~\6843(3118)  | ~\6840(2867) ,
  \3202(1566)  = ~\6550(1412)  | ~\6543(937) ,
  \1715(2391)  = \1714(2031)  | \1584(877) ,
  \6249(3673)  = ~\6243(3664) ,
  \6386(1069)  = \719(850) ,
  \3988(1770)  = ~\6916(1703)  | ~\6909(324) ,
  \2266(587)  = ~\2259(413) ,
  \5550(2401)  = ~\5546(2038) ,
  \3873(1767)  = ~\6876(1706)  | ~\6869(323) ,
  \7149(3198)  = ~\7148(3078)  | ~\7147(3142) ,
  \1007(773)  = ~\1006(602)  | ~\1005(721) ,
  \7384(1594)  = ~\7380(1257) ,
  \5634(2045)  = \1598(1817) ,
  \6678(2571)  = ~\6674(2245) ,
  \4772(2105)  = \1038(1843) ,
  \5514(3502)  = ~\5512(2377)  | ~\5505(3480) ,
  \4848(2631)  = ~\4844(2345) ,
  \7393(1319)  = \4496(999) ,
  \2145(810)  = \2124(731)  & \187(110) ,
  \281(547)  = \[53] ,
  \5278(1103)  = ~\5274(864) ,
  \6695(983)  = \3673(821) ,
  \7309(1072)  = \711(852) ,
  \944(2114)  = \868(934)  & \827(1874) ,
  \2409(1989)  = ~\2408(1793)  | ~\2407(1499) ,
  \5719(3526)  = ~\5718(3483)  | ~\5717(3506) ,
  \6964(3454)  = ~\6962(2572)  | ~\6955(3423) ,
  \2507(2337)  = \2391(1134)  & \2372(1986) ,
  \1713(2030)  = \1556(1807)  & (\1590(882)  & \1573(1810) ),
  \6844(2979)  = ~\6840(2867) ,
  \3566(1940)  = ~\6787(1621)  | ~\6784(1396) ,
  \4707(763)  = \4683(468)  | \4682(670) ,
  \3601(2856)  = \3582(2705)  & (\3536(2174)  & \3531(2480) ),
  \5287(1413)  = ~\5281(1058) ,
  \5159(3584)  = ~\5158(3544)  | ~\5157(3565) ,
  \4676(702)  = \4660(581)  & \64(27) ,
  \414(3338)  = \[70] ,
  \1262(1234)  = ~\5322(955)  | ~\5315(965) ,
  \1685(1163)  = ~\5455(475)  | ~\5452(1077) ,
  \3193(1731)  = ~\6541(1282)  | ~\6538(1055) ,
  \6840(2867)  = ~\6818(2732)  | ~\6817(2744) ,
  \4363(2465)  = \4300(2153)  & (\4314(1248)  & (\4291(2173)  & \4308(2151) )),
  \1299(2536)  = ~\1296(2212) ,
  \7289(1628)  = ~\7283(1294) ,
  \4831(3329)  = ~\4825(3257) ,
  \6663(2567)  = ~\3445(2254)  & ~\3327(1111) ,
  \7335(1742)  = ~\7333(1419)  | ~\7330(1067) ,
  \3213(1735)  = ~\6565(1223)  | ~\6562(1059) ,
  \784(559)  = \1198(299)  & \1519(374) ,
  \6171(3573)  = ~\6165(3554) ,
  \5661(3637)  = ~\5660(3598)  | ~\5659(3619) ,
  \4135(688)  = \4094(584)  & \81(40) ,
  \2990(1579)  = ~\6405(1172)  | ~\6402(951) ,
  \266(2956)  = \997(2432)  & \1790(2815) ,
  \5064(2099)  = \792(1841) ,
  \4283(2694)  = \4266(2458)  & (\4235(1855)  & \4230(2140) ),
  \5651(3638)  = ~\5650(3599)  | ~\5649(3620) ,
  \4043(2301)  = \3979(1126)  & (\3932(1975)  & \3957(1977) ),
  \4593(1889)  = ~\7573(1643)  | ~\7570(1308) ,
  \4079(3669)  = ~\7127(3660)  | ~\7124(2270) ,
  \1307(2463)  = ~\1304(2147) ,
  \6951(3313)  = ~\6945(3248) ,
  \791(1559)  = ~\4888(1460)  | ~\4881(375) ,
  \695(525)  = \657(404)  & \175(98) ,
  \1308(2752)  = \1287(2544)  & (\1226(1959)  & \1221(2222) ),
  \326(3294)  = ~\4768(2442)  | ~\4761(3233) ,
  \4281(2740)  = \4259(2487)  & (\4207(2198)  & \4216(2206) ),
  \3381(1976)  = ~\3380(1777)  | ~\3379(1480) ,
  \2617(1787)  = ~\6008(1592)  | ~\6001(340) ,
  \3046(2813)  = \3045(2651)  | \3028(2372) ,
  \7391(1662)  = ~\7385(1324) ,
  \7343(2191)  = ~\7337(1902) ,
  \7325(1746)  = ~\7323(1423)  | ~\7320(1071) ,
  \6938(2562)  = \4013(2236)  | (\4012(2255)  | (\4011(2243)  | \3868(1110) )),
  \6219(3529)  = ~\6213(3510) ,
  \4084(3627)  = \4072(3202)  & (\4028(2579)  & \4059(3604) ),
  \364(3326)  = ~\4824(2593)  | ~\4817(3254) ,
  \5756(1086)  = \751(857) ,
  \5697(3276)  = ~\5695(3219)  | ~\5692(2413) ,
  \7424(1587)  = ~\7420(1249) ,
  \6737(1360)  = \3816(1021) ,
  \3550(2199)  = ~\3549(1696)  | ~\3548(1924) ,
  \2864(3245)  = ~\2863(3127)  | ~\2862(3185) ,
  \5084(2108)  = \805(1844) ,
  \1310(2887)  = ~\1309(2545)  & ~\1308(2752) ,
  \7074(2306)  = \3997(1980) ,
  \7529(1661)  = ~\7523(1323) ,
  \5051(3471)  = ~\5050(3414)  | ~\5049(3448) ,
  \4634(2863)  = \4617(2722)  & (\4586(2182)  & \4581(2500) ),
  \6277(3130)  = ~\6271(3064) ,
  \5115(3052)  = ~\5109(2959) ,
  \5900(1288)  = \2085(986) ,
  \4045(2288)  = \3971(1124)  & \3932(1975) ,
  \5094(2106)  = \805(1844) ,
  \3452(2295)  = \3365(1973)  & (\3425(1125)  & (\3353(1972)  & (\3381(1976)  & \3399(1978) ))),
  \3679(776)  = \3659(499)  | \3658(681) ,
  \6687(943)  = \3667(779) ,
  \7307(1228)  = ~\7301(949) ,
  \261(2992)  = \3249(2223)  & (\3035(2374)  & \3164(2980) ),
  \4324(1284)  = \2065(985)  & \4499(1001) ,
  \5238(1195)  = ~\5234(918) ,
  \950(2448)  = \949(2129)  | \868(934) ,
  \4385(3060)  = ~\4382(2972) ,
  \1186(254)  = ~\2253(183) ,
  \6487(1313)  = \4154(996) ,
  \5375(3070)  = ~\5369(2989) ,
  \1253(2214)  = ~\1249(1952) ,
  \1461(287)  = ~\1459(167) ,
  \2502(2317)  = \2354(1983)  & (\2372(1986)  & \2400(1988) ),
  \1790(2815)  = \1789(2652)  | \1708(2378) ,
  \370(3718)  = \[106] ,
  \4682(670)  = \4660(581)  & \109(54) ,
  \6591(325)  = \4422(215) ,
  \4025(2277)  = \3949(1122)  & (\3899(1971)  & \3911(1974) ),
  \3215(1852)  = ~\3214(1571)  | ~\3213(1735) ,
  \3828(1035)  = \3796(725)  | \3795(797) ,
  \4035(2276)  = \3949(1122)  & \3911(1974) ,
  \2026(730)  = ~\2019(576) ,
  \4808(2583)  = ~\4804(2266) ,
  \4913(497)  = \1519(374) ,
  \915(1029)  = \784(559)  & \765(774) ,
  \306(3270)  = \1856(2037)  & \2008(3214) ,
  \3563(2517)  = ~\3559(2205) ,
  \2454(1996)  = ~\2453(1800)  | ~\2452(1506) ,
  \4997(1555)  = ~\4993(1203) ,
  \320(3711)  = ~\1792(3707)  | ~\1791(3701) ,
  \6209(3464)  = ~\6203(3437) ,
  \7540(1914)  = ~\7538(1686)  | ~\7531(1346) ,
  \2073(971)  = \2050(656)  | \2049(803) ,
  \4487(710)  = \4457(583)  & \55(18) ,
  \1981(2655)  = \1935(2004)  & \1957(2411) ,
  \3192(931)  = \641(841)  & \3676(777) ,
  \6405(1172)  = ~\6399(897) ,
  \4092(3705)  = ~\7203(3657)  | ~\7200(3699) ,
  \3583(2472)  = \3545(2155) ,
  \4751(3284)  = ~\4745(3222) ,
  \6993(3076)  = ~\6992(3002)  | ~\6991(2907) ,
  \1584(877)  = \745(853)  & \2249(255) ,
  \5392(2885)  = ~\5388(2751) ,
  \5129(3359)  = ~\5128(3231)  | ~\5127(3295) ,
  \5777(361)  = \1178(261) ,
  \7550(1910)  = ~\7548(1683)  | ~\7541(1342) ,
  \6309(3522)  = ~\6307(3509)  | ~\6304(2370) ,
  \552(238)  = \3723(190) ,
  \3618(3244)  = ~\3617(3126)  | ~\3616(3184) ,
  \3173(717)  = \1210(298)  & \2872(430) ,
  \678(414)  = \1503(303) ,
  \6872(1377)  = \3828(1035) ,
  \7408(1391)  = ~\7404(1042) ,
  \1072(1214)  = ~\5221(505)  | ~\5218(1095) ,
  \3483(2577)  = ~\6677(1474)  | ~\6674(2245) ,
  \3453(2578)  = \3452(2295)  | (\3451(2283)  | (\3450(2274)  | (\3449(2267)  | \3362(1117) ))),
  \3195(1876)  = ~\3194(1617)  | ~\3193(1731) ,
  \7213(1306)  = \2171(992) ,
  \5037(3236)  = ~\5031(3178) ,
  \4833(207)  = \4526(205) ,
  \6342(2750)  = ~\6341(2538)  | ~\6340(2539) ,
  \6168(2320)  = \2600(1984) ,
  \6602(1359)  = \3816(1021) ,
  \7219(1638)  = ~\7213(1306) ,
  \7077(3428)  = ~\7071(3378) ,
  \6148(2329)  = \2618(1985) ,
  \5823(2657)  = ~\5817(2384) ,
  \5263(1104)  = \2950(865) ,
  \2045(801)  = \2026(730)  & \204(127) ,
  \933(2683)  = ~\929(2433) ,
  \1205(305)  = \15(4) ,
  \417(3415)  = \2881(3339)  & (\2878(386)  & \2876(389) ),
  \7554(1011)  = \4123(708)  | \4122(751) ,
  \7456(2737)  = ~\7609(2507)  | ~\7606(2197) ,
  \4801(3250)  = \3459(3196)  | (\3458(2294)  | (\3457(2282)  | (\3456(2273)  | \3376(1119) ))),
  \6502(1371)  = ~\6498(1032) ,
  \5685(3042)  = ~\5679(2951) ,
  \2146(661)  = \2117(577)  & \118(61) ,
  \6164(3517)  = ~\6162(2604)  | ~\6155(3499) ,
  \347(3420)  = \[100] ,
  \4015(2257)  = \3856(1966)  & (\3891(1114)  & \3874(1968) ),
  \319(3398)  = \[80] ,
  \6869(323)  = \4429(213) ,
  \5968(2613)  = ~\5964(2315) ,
  \626(636)  = \625(534)  | \611(573) ,
  \650(423)  = \1206(306) ,
  \7051(3007)  = ~\7050(2914)  | ~\7049(2781) ,
  \2955(1508)  = ~\6374(1420)  | ~\6367(869) ,
  \2762(2326)  = \2629(1133)  & \2600(1984) ,
  \5038(2686)  = ~\5034(2444) ,
  \5699(3347)  = ~\5698(3215)  | ~\5697(3276) ,
  \4137(746)  = \4114(735)  & \4417(217) ,
  \3442(2251)  = \3295(1965)  & (\3314(1967)  & \3335(1113) ),
  \4298(1867)  = ~\7375(1682)  | ~\7372(1263) ,
  \6064(2924)  = ~\6060(2799) ,
  \885(832)  = ~\4919(605)  | ~\4916(400) ,
  \3649(511)  = \3622(407)  & \1461(287) ,
  \2597(1129)  = \2111(987)  & \3751(229) ,
  \6989(1769)  = ~\6983(1470) ,
  \3398(1779)  = ~\6630(1631)  | ~\6623(333) ,
  \3397(1482)  = ~\6629(446)  | ~\6626(1297) ,
  \4040(2285)  = \3911(1974)  & (\3971(1124)  & \3932(1975) ),
  \5552(3272)  = ~\5550(2401)  | ~\5543(3212) ,
  \3899(1971)  = ~\3898(1772)  | ~\3897(1475) ,
  \5030(3051)  = ~\5028(2842)  | ~\5021(2960) ,
  \4704(764)  = \4681(471)  | \4680(683) ,
  \2817(3590)  = ~\6113(3574)  | ~\6110(2318) ,
  \6138(2342)  = \2734(1987) ,
  \3635(408)  = \1524(301) ,
  \2354(1983)  = ~\2353(1785)  | ~\2352(1489) ,
  \7578(1312)  = \4166(995) ,
  \7518(1322)  = \4490(1000) ,
  \4986(2742)  = ~\4980(2511) ,
  \5992(1625)  = ~\5988(1290) ,
  \3209(942)  = \629(844)  & \3667(779) ,
  \1702(1999)  = \1546(1803)  & (\1556(1807)  & (\1573(1810)  & \1687(1813) )),
  \4849(2807)  = \2526(2549)  | (\2524(2525)  | (\2523(2363)  | \2448(1142) )),
  \5182(563)  = ~\5178(399) ,
  \4836(2745)  = \2472(2532) ,
  \2970(872)  = \723(849)  & \4707(763) ,
  \6613(441)  = ~\6607(328) ,
  \2298(716)  = \2272(594)  & \41(12) ,
  \6299(3472)  = ~\6297(3436)  | ~\6294(2746) ,
  \2258(249)  = ~\2256(184) ,
  \3170(866)  = ~\3169(597)  | ~\3168(828) ,
  \5127(3295)  = ~\5125(3234)  | ~\5122(2443) ,
  \2921(512)  = \2892(416)  & \216(139) ,
  \7020(2573)  = ~\7016(2249) ,
  \1276(2145)  = ~\1272(1858) ,
  \3265(3034)  = \1974(2382)  & \3468(2898) ,
  \709(545)  = \678(414)  & \153(76) ,
  \7446(2726)  = ~\7617(2506)  | ~\7614(2181) ,
  \7441(3039)  = ~\7433(2949) ,
  \6075(3205)  = ~\6073(3150)  | ~\6070(2612) ,
  \7010(2575)  = ~\7006(2259) ,
  \6055(1403)  = ~\6049(1049) ,
  \5088(2447)  = ~\5084(2108) ,
  \6772(1363)  = ~\6768(1023) ,
  \6860(1665)  = ~\6856(1327) ,
  \2198(974)  = \2162(659)  | \2161(794) ,
  \6291(3385)  = ~\6290(3262)  | ~\6289(3335) ,
  \6201(3386)  = ~\6199(3337)  | ~\6196(2806) ,
  \5098(2446)  = ~\5094(2106) ,
  \6698(938)  = \3670(778) ,
  \5089(3621)  = ~\5165(3600)  | ~\5162(2166) ,
  \4713(3136)  = \3279(3072) ,
  \7031(3530)  = ~\7029(3514)  | ~\7026(2225) ,
  \2288(555)  = \2259(413)  & \41(12) ,
  \6753(1932)  = ~\6751(1705)  | ~\6748(1373) ,
  \4351(1917)  = ~\7424(1587)  | ~\7417(1349) ,
  \4942(1551)  = \914(1200)  | (\913(1027)  | \777(370) ),
  \792(1841)  = ~\791(1559)  | ~\790(1208) ,
  \2563(2756)  = \4526(205)  & \2508(2630) ,
  \3598(2692)  = \3578(2437)  & (\3517(2120)  & \3504(1851) ),
  \5501(3441)  = ~\5495(3392) ,
  \1868(1529)  = ~\5792(1243)  | ~\5785(362) ,
  \1858(1528)  = ~\5784(1436)  | ~\5777(361) ,
  \7263(1393)  = ~\7257(1043) ,
  \7588(1336)  = \4172(1008) ,
  \7091(3532)  = ~\7090(3494)  | ~\7089(3515) ,
  \386(3020)  = ~\4847(2932)  | ~\4844(2345) ,
  \5079(3622)  = ~\5077(3601)  | ~\5074(2167) ,
  \5068(2440)  = ~\5064(2099) ,
  \3798(713)  = \3768(595)  & \50(15) ,
  \3676(777)  = \3657(504)  | \3656(667) ,
  \327(3408)  = \[81] ,
  \1755(3580)  = ~\5521(3560)  | ~\5518(2011) ,
  \1217(1960)  = ~\1216(1757)  | ~\1215(1758) ,
  \5044(2136)  = \895(1850) ,
  \6482(1304)  = \2171(992) ,
  \1820(1157)  = ~\5767(473)  | ~\5764(1075) ,
  \4020(2264)  = \3899(1971)  & (\3911(1974)  & (\3932(1975)  & (\3957(1977)  & \3997(1980) ))),
  \2046(673)  = \2019(576)  & \103(52) ,
  \7203(3657)  = ~\7197(3642) ,
  \5800(1239)  = ~\5796(960) ,
  \2642(1794)  = ~\6016(1622)  | ~\6009(345) ,
  \4178(1872)  = ~\7211(1609)  | ~\7208(978) ,
  \2853(2784)  = \2780(2629)  & \2749(2307) ,
  \7470(915)  = ~\7466(771) ,
  \2899(590)  = ~\2892(416) ,
  \3240(3026)  = \3035(2374)  & (\3156(2706)  & \4388(2971) ),
  \1834(878)  = \745(853)  & \2249(255) ,
  \1608(1530)  = ~\5432(1242)  | ~\5425(363) ,
  \4188(1887)  = ~\7220(1633)  | ~\7213(1306) ,
  \246(3110)  = \[57] ,
  \1073(1565)  = ~\5222(1450)  | ~\5215(379) ,
  \2137(738)  = ~\2130(593) ,
  \3271(3101)  = \3270(2892)  | (\3267(3035)  | (\3265(3034)  | \1982(2816) )),
  \4732(2051)  = \1869(1819) ,
  \5600(3041)  = ~\5598(2831)  | ~\5591(2952) ,
  \1406(817)  = \1378(538)  | \1377(649) ,
  \1382(540)  = \1350(415)  & \158(81) ,
  \6367(869)  = \4710(762) ,
  \5054(2121)  = \853(1849) ,
  \7610(2508)  = ~\7606(2197) ,
  \3146(2871)  = ~\3143(2738) ,
  \6049(1049)  = \3682(839) ,
  \6763(1918)  = ~\6761(1666)  | ~\6758(1351) ,
  \7040(2566)  = ~\7036(2237) ,
  \7030(2554)  = ~\7026(2225) ,
  \304(3390)  = \[89] ,
  \3342(1473)  = ~\6597(438)  | ~\6594(1375) ,
  \3989(1969)  = ~\3988(1770)  | ~\3987(1472) ,
  \6041(342)  = \3731(235) ,
  \4660(581)  = ~\4653(410) ,
  \7558(1341)  = ~\7554(1011) ,
  \3120(1871)  = ~\6509(1649)  | ~\6506(1272) ,
  \3788(552)  = \3755(412)  & \50(15) ,
  \5953(2618)  = \2506(2332)  | (\2505(2336)  | \2384(1132) ),
  \4202(1362)  = ~\7256(1022)  | ~\7249(1024) ,
  \1171(3307)  = \1155(2201)  & \1161(3229) ,
  \6912(1374)  = \3821(1034) ,
  \6154(3461)  = ~\6152(2621)  | ~\6145(3434) ,
  \1379(645)  = \1357(589)  & \144(71) ,
  \4373(2519)  = \4341(1392)  & (\4317(2170)  & \4327(2186) ),
  \362(3429)  = \[97] ,
  \1736(2053)  = \1655(1827)  & (\1609(1820)  & (\1630(1824)  & \1695(1829) )),
  \6199(3337)  = ~\6193(3263) ,
  \7282(1865)  = ~\7280(1586)  | ~\7273(1258) ,
  \5936(1949)  = ~\5932(1726) ,
  \6832(1546)  = ~\6720(1189)  | ~\6719(1202) ,
  \6645(2762)  = ~\6639(2560) ,
  \3123(2497)  = \3052(2192)  & (\3062(2194)  & (\3071(2195)  & \3119(2180) )),
  \4987(1549)  = ~\4983(1191) ,
  \4671(488)  = \4640(409)  & \2220(266) ,
  \6533(1212)  = ~\6527(932) ,
  \2796(2529)  = \2724(1722)  & (\2676(1994)  & \2701(1995) ),
  \5988(1290)  = \2111(987) ,
  \3069(1934)  = ~\6461(1676)  | ~\6458(1036) ,
  \3343(1771)  = ~\6598(1704)  | ~\6591(325) ,
  \6158(2308)  = \2589(1981) ,
  \7458(2870)  = ~\7457(2736)  | ~\7456(2737) ,
  \6693(1222)  = ~\6687(943) ,
  \1365(644)  = \1343(575)  & \147(72) ,
  \5712(2077)  = \1655(1827) ,
  \6327(3612)  = ~\6321(3592) ,
  \2526(2549)  = \2454(1996)  & (\2436(1993)  & (\2472(2532)  & \4526(205) )),
  \3100(1886)  = ~\6485(1678)  | ~\6482(1304) ,
  \6899(443)  = ~\6893(330) ,
  \3874(1968)  = ~\3873(1767)  | ~\3872(1468) ,
  \4970(718)  = \784(559) ,
  \3833(1016)  = \3798(713)  | \3797(798) ,
  \2822(3591)  = ~\6171(3573)  | ~\6168(2320) ,
  \5234(918)  = \1007(773) ,
  \5266(1091)  = \2946(858) ,
  \1477(394)  = ~\1475(295) ,
  \1141(2133)  = \1102(940)  & \1074(1846) ,
  \5338(1241)  = ~\5334(962) ,
  \3327(1111)  = \3828(1035)  & \4429(213) ,
  \5607(3221)  = ~\5601(3166) ,
  \877(939)  = \2933(861)  & \1464(285) ,
  \3578(2437)  = ~\3575(2095) ,
  \7448(2862)  = ~\7447(2735)  | ~\7446(2726) ,
  \4123(708)  = \4094(584)  & \58(21) ,
  \7523(1323)  = \4499(1001) ,
  \4905(380)  = \1471(283) ,
  \5709(3467)  = ~\5708(3399)  | ~\5707(3442) ,
  \5872(1626)  = ~\5868(1291) ,
  \7167(3458)  = ~\7165(3427)  | ~\7162(2305) ,
  \6289(3335)  = ~\6287(3264)  | ~\6284(2635) ,
  \698(629)  = \697(526)  | \664(574) ,
  \7513(1325)  = ~\7507(1002) ,
  \6807(1866)  = ~\6805(1624)  | ~\6802(1261) ,
  \1988(2818)  = ~\5831(2656)  | ~\5828(2003) ,
  \2301(783)  = \2279(739)  & \237(160) ,
  \4621(2724)  = ~\4618(2496) ,
  \3099(1268)  = \2175(975)  & \4160(993) ,
  \4134(747)  = \4101(734)  & \4412(219) ,
  \3435(2238)  = \3327(1111)  & (\3283(1964)  & \3295(1965) ),
  \5727(3563)  = ~\5725(3543)  | ~\5722(2044) ,
  \5448(1236)  = ~\5444(957) ,
  \5468(2665)  = \1749(2022)  | \1715(2391) ,
  \5581(911)  = ~\1399(820)  & ~\2213(268) ,
  \2587(1487)  = ~\5991(449)  | ~\5988(1290) ,
  \5880(1596)  = ~\5876(1259) ,
  \2559(2624)  = ~\5983(1789)  | ~\5980(2330) ,
  \4685(465)  = \4653(410)  & \2258(249) ,
  \2323(1038)  = \2300(726)  | \2299(782) ,
  \7351(2471)  = ~\7345(2154) ,
  \4476(758)  = \4451(732)  & \3713(241) ,
  \4701(765)  = \4679(476)  | \4678(703) ,
  \7292(1881)  = ~\7290(1600)  | ~\7283(1294) ,
  \1519(374)  = ~\1518(278) ,
  \5078(2484)  = ~\5074(2167) ,
  \3497(3319)  = ~\3491(3249) ,
  \354(3375)  = \3497(3319)  & \3344(1970) ,
  \4595(2178)  = ~\4594(1890)  | ~\4593(1889) ,
  \6797(1862)  = ~\6795(1591)  | ~\6792(1252) ,
  \6735(1634)  = ~\6729(1301) ,
  \3520(1564)  = ~\6709(1206)  | ~\6706(933) ,
  \2840(3671)  = ~\6259(3663)  | ~\6256(2350) ,
  \2652(1139)  = \2085(986)  & \3725(237) ,
  \5049(3448)  = ~\5047(3410)  | ~\5044(2136) ,
  \344(3382)  = \[91] ,
  \5744(3698)  = ~\5740(3694) ,
  \3110(2175)  = ~\3109(1892)  | ~\3108(1883) ,
  \2612(1131)  = \2105(972)  & \3745(231) ,
  \5074(2167)  = \827(1874) ,
  \1760(3581)  = ~\5579(3559)  | ~\5576(2013) ,
  \6210(2881)  = ~\6206(2747) ,
  \4379(2854)  = ~\4376(2714) ,
  \5067(3546)  = ~\5061(3527) ,
  \2471(2209)  = ~\5936(1949)  | ~\5929(1048) ,
  \3312(1467)  = ~\6589(435)  | ~\6586(1378) ,
  \4220(1619)  = ~\7272(1399)  | ~\7265(1285) ,
  \1447(3100)  = \1445(2895)  | (\1440(3030)  | (\1436(3029)  | \1790(2815) )),
  \1687(1813)  = ~\1686(1522)  | ~\1685(1163) ,
  \3241(2859)  = \3035(2374)  & (\3156(2706)  & (\4386(2698)  & \89(48) )),
  \2192(991)  = \2160(679)  | \2159(793) ,
  \2004(2666)  = ~\5864(2397)  | ~\5857(1159) ,
  \1332(3134)  = ~\5391(3055)  | ~\5388(2751) ,
  \5732(2063)  = \1630(1824) ,
  \274(3353)  = \961(3291)  & \957(1836) ,
  \6430(1425)  = ~\6426(1070) ,
  \2795(2368)  = \2715(1145)  & \2676(1994) ,
  \1741(2083)  = \1677(909)  & (\1630(1824)  & \1655(1827) ),
  \4028(2579)  = \4027(2299)  | (\4026(2287)  | (\4025(2277)  | (\4024(2268)  | \3908(1118) ))),
  \3719(239)  = ~\3717(189) ,
  \6485(1678)  = ~\6479(1339) ,
  \4547(1532)  = ~\7485(1166)  | ~\7482(898) ,
  \3665(600)  = \3642(579)  & \3703(245) ,
  \269(2896)  = \997(2432)  & (\1788(2375)  & (\4089(2553)  & (\2852(2785)  & \4526(205) ))),
  \5649(3620)  = ~\5647(3597)  | ~\5644(2064) ,
  \1708(2378)  = \1707(2029)  | (\1706(2015)  | (\1705(2010)  | \1553(870) )),
  \6024(1718)  = ~\6020(1395) ,
  \6445(1670)  = ~\6439(1333) ,
  \314(3350)  = ~\4743(3282)  | ~\4740(2066) ,
  \5905(347)  = \3719(239) ,
  \6826(2467)  = ~\6822(2150) ,
  \5376(1961)  = ~\5372(1759) ,
  \1788(2375)  = \1718(2046)  & \1702(1999) ,
  \5245(830)  = ~\5239(719) ,
  \2081(988)  = \2054(676)  | \2053(805) ,
  \560(248)  = \3698(185) ,
  \5105(1569)  = ~\5099(1218) ,
  \2418(1502)  = ~\5911(460)  | ~\5908(1394) ,
  \3313(1766)  = ~\6590(1707)  | ~\6583(322) ,
  \802(924)  = \2950(865)  & \1488(279) ,
  \7428(1404)  = \3695(1050) ,
  \6319(3577)  = ~\6317(3558)  | ~\6314(2346) ,
  \995(3691)  = \980(3210)  & \990(3685) ,
  \572(427)  = \573(311) ,
  \1174(3290)  = \1023(1205)  & \1161(3229) ,
  \6144(3333)  = ~\6142(2625)  | ~\6135(3260) ,
  \5638(2409)  = ~\5634(2045) ,
  \324(3363)  = \[74] ,
  \7087(3497)  = ~\7081(3477) ,
  \1018(606)  = ~\5190(562)  | ~\5183(498) ,
  \334(3362)  = ~\4791(3301)  | ~\4788(2118) ,
  \5659(3619)  = ~\5735(3596)  | ~\5732(2063) ,
  \4884(1105)  = \2950(865) ,
  \5048(2454)  = ~\5044(2136) ,
  \6974(3512)  = ~\6972(2555)  | ~\6965(3492) ,
  \3114(1298)  = \2167(990)  & \4154(996) ,
  \4511(1012)  = \4489(709)  | \4488(752) ,
  \6805(1624)  = ~\6799(1289) ,
  \5647(3597)  = ~\5641(3583) ,
  \7022(3455)  = ~\7020(2573)  | ~\7013(3422) ,
  \4626(2404)  = \4602(2041)  & (\4535(2093)  & \4544(2062) ),
  \1017(831)  = ~\5189(607)  | ~\5186(398) ,
  \6390(1424)  = ~\6386(1069) ,
  \5199(377)  = \1482(281) ,
  \1956(2087)  = \1869(1819)  & (\1929(910)  & (\1859(1818)  & (\1885(1825)  & \1903(1826) ))),
  \7257(1043)  = \2312(836) ,
  \286(419)  = \[49] ,
  \6115(1494)  = \2635(1135) ,
  \1966(2089)  = \1929(910)  & (\1885(1825)  & \1903(1826) ),
  \5675(1541)  = ~\5669(1182) ,
  \5536(2387)  = ~\1713(2030)  & (~\1712(2014)  & ~\1567(876) ),
  \3594(2719)  = ~\3591(2490) ,
  \5785(362)  = \2232(262) ,
  \6900(1635)  = ~\6896(1302) ,
  \5396(1084)  = \757(856) ,
  \1507(418)  = ~\1503(303) ,
  \2859(3133)  = ~\6345(3054)  | ~\6342(2750) ,
  \6252(3614)  = ~\6328(2642)  | ~\6321(3592) ,
  \1151(2681)  = \1108(1196)  & \1129(2434) ,
  \5058(2451)  = ~\5054(2121) ,
  \3020(1543)  = ~\6438(1233)  | ~\6431(914) ,
  \6877(326)  = \4417(217) ,
  \3362(1117)  = \3816(1021)  & \4417(217) ,
  \4761(3233)  = \1136(3174)  | (\1134(2131)  | (\1133(2115)  | (\1132(2164)  | \1050(930) ))),
  \2531(2547)  = \2472(2532)  & \4526(205) ,
  \4624(2829)  = ~\4623(2420)  & ~\4622(2673) ,
  \5377(2988)  = ~\1316(2882)  | ~\1319(2883) ,
  \3440(2234)  = \3295(1965)  & (\3314(1967)  & \3344(1970) ),
  \2154(664)  = \2130(593)  & \115(60) ,
  \6373(1147)  = ~\6367(869) ,
  \7399(1656)  = ~\7393(1319) ,
  \4932(1547)  = \953(1197)  | \917(1190) ,
  \7135(1780)  = ~\7129(1483) ,
  \5648(2422)  = ~\5644(2064) ,
  \2053(805)  = \2026(730)  & \200(123) ,
  \3568(2172)  = ~\3567(1878)  | ~\3566(1940) ,
  \294(3223)  = ~\4720(2430)  | ~\4713(3136) ,
  \4023(2582)  = ~\4020(2264) ,
  \2871(315)  = \1458(289)  & \4528(206) ,
  \3090(1356)  = \3801(824)  & \4163(994) ,
  \3543(1869)  = ~\6743(1693)  | ~\6740(1265) ,
  \379(3207)  = \[66] ,
  \5702(2090)  = \1695(1829) ,
  \6242(3635)  = ~\6240(2643)  | ~\6233(3613) ,
  \6779(1713)  = ~\6773(1388) ,
  \6192(3154)  = ~\6190(2939)  | ~\6183(3131) ,
  \5628(2426)  = ~\5624(2076) ,
  \6848(2851)  = ~\6828(2701)  | ~\6827(2700) ,
  \6007(453)  = ~\6001(340) ,
  \6559(944)  = \3667(779) ,
  \6462(1380)  = ~\6458(1036) ,
  \4274(2852)  = \4254(2708)  & (\4193(2493)  & \4180(2159) ),
  \5618(2429)  = ~\5614(2091) ,
  \3512(1616)  = ~\6702(1216)  | ~\6695(983) ,
  \3484(2772)  = ~\6678(2571)  | ~\6671(1116) ,
  \3006(901)  = \1391(813)  & \4692(768) ,
  \3000(1534)  = ~\6414(1229)  | ~\6407(903) ,
  \5668(2416)  = ~\5664(2052) ,
  \5658(2417)  = ~\5654(2054) ,
  \6510(1607)  = ~\6506(1272) ,
  \5147(3508)  = ~\5145(3488)  | ~\5142(2123) ,
  \4230(2140)  = ~\4226(1854) ,
  \7606(2197)  = ~\7540(1914)  | ~\7539(1916) ,
  \908(1192)  = \907(1028)  | \777(370) ,
  \1272(1858)  = ~\1271(1584)  | ~\1270(1583) ,
  \2342(1784)  = ~\5872(1626)  | ~\5865(337) ,
  \6431(914)  = \4686(770) ,
  \408(385)  = \[44] ,
  \3399(1978)  = ~\3398(1779)  | ~\3397(1482) ,
  \3203(1847)  = ~\3202(1566)  | ~\3201(1733) ,
  \5221(505)  = ~\5215(379) ,
  \895(1850)  = ~\894(1570)  | ~\893(1220) ,
  \3018(1814)  = ~\3017(1524)  | ~\3016(1745) ,
  \5190(562)  = ~\5186(398) ,
  \1789(2652)  = \1726(2407)  & \1702(1999) ,
  \6819(2152)  = ~\6808(1879)  | ~\6807(1866) ,
  \5222(1450)  = ~\5218(1095) ,
  \1606(892)  = \731(855)  & \1178(261) ,
  \7333(1419)  = ~\7327(1064) ,
  \937(2162)  = \845(980)  & \805(1844) ,
  \6229(3579)  = ~\6223(3557) ,
  \3485(2909)  = ~\3484(2772)  | ~\3483(2577) ,
  \3654(682)  = \3629(578)  & \87(46) ,
  \4243(1747)  = ~\7316(1231)  | ~\7309(1072) ,
  \5449(359)  = \2241(257) ,
  \5407(470)  = ~\5401(355) ,
  \3475(3074)  = ~\3474(2998) ,
  \2287(620)  = \2266(587)  & \198(121) ,
  \5752(1440)  = ~\5748(1085) ,
  \2465(1144)  = \2323(1038)  & \3707(243) ,
  \7323(1423)  = ~\7317(1068) ,
  \6674(2245)  = \3314(1967) ,
  \4721(3217)  = \1964(3162)  | (\1962(2086)  | (\1961(2072)  | (\1960(2059)  | \1880(895) ))),
  \4131(748)  = \4101(734)  & \4407(221) ,
  \4780(2168)  = \1055(1875) ,
  \3238(2684)  = ~\3235(2435) ,
  \5262(1452)  = ~\5258(1097) ,
  \4008(2242)  = \3885(1112)  & (\3845(1963)  & \3856(1966) ),
  \5868(1291)  = \2111(987) ,
  \280(391)  = \575(309)  & \1184(294) ,
  \6621(444)  = ~\6615(331) ,
  \765(774)  = ~\764(603)  | ~\763(723) ,
  \1126(2165)  = \1068(981)  & (\1026(1842)  & \1038(1843) ),
  \5943(2791)  = ~\5937(2610) ,
  \620(633)  = \619(531)  | \594(572) ,
  \4958(3048)  = ~\4956(1556)  | ~\4949(2954) ,
  \4266(2458)  = ~\4263(2142) ,
  \4479(694)  = \4444(582)  & \75(34) ,
  \1782(3616)  = \1771(3137)  & (\1730(2668)  & \1762(3595) ),
  \488(260)  = \2236(180) ,
  \1946(2033)  = \1805(1806)  & (\1822(1811)  & \1841(883) ),
  \4353(1720)  = ~\7431(1401)  | ~\7428(1404) ,
  \4242(1580)  = ~\7315(1427)  | ~\7312(952) ,
  \985(3653)  = ~\5088(2447)  | ~\5081(3640) ,
  \7101(3589)  = ~\7100(3551)  | ~\7099(3572) ,
  \5856(2398)  = ~\5852(2026) ,
  \5807(486)  = ~\5801(366) ,
  \5152(2098)  = \792(1841) ,
  \7242(1018)  = \3810(823) ,
  \6056(1948)  = ~\6052(1725) ,
  \4776(2445)  = ~\4772(2105) ,
  \4297(1293)  = \2081(988)  & \4511(1012) ,
  \7412(1039)  = \2308(835) ,
  \7147(3142)  = ~\7145(3080)  | ~\7142(2778) ,
  \2942(859)  = \2886(425)  & \2924(610) ,
  \6297(3436)  = ~\6291(3385) ,
  \6406(1230)  = ~\6402(951) ,
  \617(530)  = \587(402)  & \169(92) ,
  \4048(2594)  = \4047(2302)  | \3971(1124) ,
  \5717(3506)  = ~\5715(3484)  | ~\5712(2077) ,
  \6945(3248)  = ~\6944(3139)  | ~\6943(3194) ,
  \5020(2844)  = ~\5018(2713)  | ~\5011(941) ,
  \4736(2415)  = ~\4732(2051) ,
  \278(536)  = \[55] ,
  \2926(611)  = \2925(514)  | \2899(590) ,
  \5237(720)  = ~\5231(561) ,
  \3175(1558)  = ~\6526(1418)  | ~\6519(928) ,
  \703(542)  = \678(414)  & \156(79) ,
  \538(224)  = \4400(197) ,
  \4847(2932)  = ~\4841(2804) ,
  \398(3713)  = ~\2856(3709)  | ~\2855(3703) ,
  \5281(1058)  = \629(844) ,
  \1989(2654)  = ~\5832(2381)  | ~\5825(2383) ,
  \5956(2316)  = \2354(1983) ,
  \1961(2072)  = \1869(1819)  & (\1914(905)  & \1885(1825) ),
  \3491(3249)  = \3490(3195)  | \3453(2578) ,
  \2054(676)  = \2019(576)  & \100(51) ,
  \1822(1811)  = ~\1821(1518)  | ~\1820(1157) ,
  \5331(1080)  = \731(855) ,
  \3662(601)  = \3642(579)  & \2204(174) ,
  \338(3716)  = \[105] ,
  \6336(3704)  = ~\6332(3697) ,
  \6268(2808)  = ~\6264(2640) ,
  \3233(2119)  = \3186(1845)  & (\3207(936)  & (\3176(1840)  & \3195(1876) )),
  \3792(714)  = \3768(595)  & \47(14) ,
  \4698(766)  = \4677(477)  | \4676(702) ,
  \7156(2774)  = ~\7152(2584) ,
  \7136(2776)  = ~\7132(2589) ,
  \7212(1277)  = ~\7208(978) ,
  \1368(520)  = \1336(405)  & \180(103) ,
  \893(1220)  = ~\4927(508)  | ~\4924(1099) ,
  \3292(1107)  = \3838(1004)  & \4439(209) ,
  \5921(351)  = \3707(243) ,
  \4356(2466)  = \4291(2173)  & (\4300(2153)  & (\4308(2151)  & \4352(2149) )),
  \7372(1263)  = \2077(973) ,
  \391(3094)  = \[62] ,
  \803(1211)  = ~\4895(503)  | ~\4892(1090) ,
  \7232(1033)  = \3804(833) ,
  \3657(504)  = \3622(407)  & \1482(281) ,
  \4601(2406)  = ~\4598(2042) ,
  \3619(3181)  = ~\6851(3120)  | ~\6848(2851) ,
  \4799(3259)  = ~\4793(3203) ,
  \247(3310)  = \3248(3293)  & \3244(1962) ,
  \3670(778)  = \3653(506)  | \3652(668) ,
  \2032(592)  = \1507(418) ,
  \6288(2805)  = ~\6284(2635) ,
  \6506(1272)  = \2163(976) ,
  \3604(2853)  = \3586(2704)  & (\3540(2491)  & \3527(2160) ),
  \1225(1755)  = ~\5262(1452)  | ~\5255(1092) ,
  \381(3092)  = \2558(3017)  & \2564(2929) ,
  \6135(3260)  = ~\6134(3146)  | ~\6133(3204) ,
  \5879(451)  = ~\5873(338) ,
  \4828(2293)  = \3399(1978) ,
  \927(2112)  = \805(1844)  & (\868(934)  & (\792(1841)  & \827(1874) )),
  \6630(1631)  = ~\6626(1297) ,
  \6954(3316)  = ~\6952(2576)  | ~\6945(3248) ,
  \5018(2713)  = ~\5014(2482) ,
  \2732(1496)  = ~\6047(455)  | ~\6044(1251) ,
  \947(2113)  = \868(934)  & \827(1874) ,
  \1458(289)  = ~\1455(166) ,
  \7179(3533)  = ~\7178(3495)  | ~\7177(3516) ,
  \7500(873)  = \4707(763) ,
  \2407(1499)  = ~\5903(457)  | ~\5900(1288) ,
  \1050(930)  = \2946(858)  & \1482(281) ,
  \894(1570)  = ~\4928(1454)  | ~\4921(381) ,
  \5617(3395)  = ~\5611(3348) ,
  \252(3450)  = \[75] ,
  \7611(2193)  = ~\7594(1904)  | ~\7593(1905) ,
  \371(2754)  = ~\4839(316)  | ~\4836(2745) ,
  \3221(557)  = \1210(298)  & \2883(314) ,
  \3787(624)  = \3762(586)  & \190(113) ,
  \4809(3253)  = \3462(3197)  | (\3461(2297)  | (\3460(2284)  | \3393(1121) )),
  \1215(1758)  = ~\5253(1453)  | ~\5250(1101) ,
  \3185(1563)  = ~\6534(1408)  | ~\6527(932) ,
  \524(210)  = \4437(204) ,
  \4046(2303)  = \3979(1126)  & (\3932(1975)  & \3957(1977) ),
  \953(1197)  = \765(774)  & \887(922) ,
  \1524(301)  = \18(5) ,
  \4602(2041)  = \4549(1815) ,
  \1856(2037)  = ~\1850(1812) ,
  \3782(553)  = \3755(412)  & \47(14) ,
  \4286(2693)  = \4270(2459)  & (\4239(2141)  & \4226(1854) ),
  \804(1562)  = ~\4896(1445)  | ~\4889(378) ,
  \5242(917)  = \1007(773) ,
  \2167(990)  = \2148(678)  | \2147(807) ,
  \4335(1653)  = ~\7408(1391)  | ~\7401(1318) ,
  \7485(1166)  = ~\7479(890) ,
  \6087(3435)  = ~\6086(3334)  | ~\6085(3384) ,
  \438(274)  = \1496(173) ,
  \5696(2669)  = ~\5692(2413) ,
  \4386(2698)  = \4369(2486)  & \4356(2466) ,
  \3244(1962)  = ~\3220(1761)  | ~\3227(1925) ,
  \3795(797)  = \3775(740)  & \221(144) ,
  \3152(3305)  = \3150(3241)  & \3146(2871) ,
  \6809(2190)  = ~\6764(1901)  | ~\6763(1918) ,
  \5311(1060)  = ~\5305(845) ,
  \7574(1640)  = ~\7570(1308) ,
  \3344(1970)  = ~\3343(1771)  | ~\3342(1473) ,
  \4640(409)  = \1524(301) ,
  \3596(2450)  = \3571(2096)  & (\3504(1851)  & \3513(1848) ),
  \6375(874)  = \4707(763) ,
  \7108(2592)  = ~\7104(2279) ,
  \6394(1073)  = \711(852) ,
  \4484(754)  = \4464(733)  & \3739(233) ,
  \6261(1944)  = \2724(1722) ,
  \7121(3643)  = ~\7120(3608)  | ~\7119(3631) ,
  \3016(1745)  = ~\6429(1165)  | ~\6426(1070) ,
  \367(3328)  = ~\4832(2597)  | ~\4825(3257) ,
  \4637(2864)  = \4621(2724)  & (\4590(2499)  & \4577(2183) ),
  \5428(963)  = \1418(819) ,
  \1313(2886)  = ~\1312(2542)  & ~\1311(2753) ,
  \5526(2662)  = ~\1715(2391) ,
  \5000(3169)  = ~\4999(3047)  | ~\4998(3111) ,
  \2001(2825)  = ~\2000(2667)  | ~\1999(2400) ,
  \2845(3626)  = \2833(317)  & (\2780(2629)  & \2819(3610) ),
  \4361(2470)  = \4305(1262)  & \4291(2173) ,
  \1373(648)  = \1357(589)  & \141(70) ,
  \7111(3644)  = ~\7110(3609)  | ~\7109(3632) ,
  \5619(3443)  = ~\5617(3395)  | ~\5614(2091) ,
  \1848(1160)  = ~\5775(474)  | ~\5772(1078) ,
  \4470(761)  = \4451(732)  & \3700(247) ,
  \329(3298)  = ~\4776(2445)  | ~\4769(3242) ,
  \2867(3239)  = ~\2866(3115)  | ~\2865(3180) ,
  \5139(3470)  = ~\5138(3413)  | ~\5137(3447) ,
  \7098(2581)  = ~\7094(2263) ,
  \4299(1912)  = ~\7376(1599)  | ~\7369(1344) ,
  \6721(1274)  = \2179(977) ,
  \4888(1460)  = ~\4884(1105) ,
  \1706(2015)  = \1584(877)  & (\1546(1803)  & \1556(1807) ),
  \5912(1717)  = ~\5908(1394) ,
  \1296(2212)  = \1258(1951) ,
  \3544(1922)  = ~\6744(1601)  | ~\6737(1360) ,
  \4402(223)  = ~\4400(197) ,
  \4364(2720)  = \4363(2465)  | (\4362(2468)  | (\4361(2470)  | \4297(1293) )),
  \422(3451)  = \1172(3419) ,
  \5118(3050)  = ~\5116(2840)  | ~\5109(2959) ,
  \4499(1001)  = \4481(696)  | \4480(756) ,
  \4038(2271)  = \3957(1977)  & (\3911(1974)  & (\3932(1975)  & \3997(1980) )),
  \1567(876)  = \751(857)  & \1186(254) ,
  \4521(3186)  = ~\7461(3125)  | ~\7458(2870) ,
  \992(3404)  = \980(3210)  & (\929(2433)  & \967(3355) ),
  \4219(1942)  = ~\7271(1620)  | ~\7268(1046) ,
  \6646(2556)  = ~\6642(2227) ,
  \5841(2392)  = ~\1949(2036)  & ~\1834(878) ,
  \4129(691)  = \4094(584)  & \78(37) ,
  \4924(1099)  = \2933(861) ,
  \692(626)  = \691(523)  | \664(574) ,
  \2965(1805)  = ~\2964(1512)  | ~\2963(1741) ,
  \2556(2801)  = ~\5976(2623)  | ~\5969(1137) ,
  \5532(2946)  = ~\5530(2821)  | ~\5523(1158) ,
  \5157(3565)  = ~\5155(3547)  | ~\5152(2098) ,
  \3127(2725)  = ~\3123(2497) ,
  \5975(1498)  = ~\5969(1137) ,
  \7593(1905)  = ~\7591(1671)  | ~\7588(1336) ,
  \4524(3265)  = \4523(3246)  & (\4520(3243)  & (\4517(3156)  & \3615(3168) )),
  \6701(1281)  = ~\6695(983) ,
  \3027(2040)  = \2965(1805)  & (\2979(886)  & (\2956(1802)  & \2973(1808) )),
  \5355(1438)  = ~\5349(1083) ,
  \5637(3542)  = ~\5631(3525) ,
  \5751(467)  = ~\5745(353) ,
  \4382(2972)  = \4380(2721)  & \4379(2854) ,
  \6781(1286)  = \2085(986) ,
  \254(2888)  = \3249(2223)  & \3046(2813) ,
  \2255(252)  = ~\2253(183) ,
  \5932(1726)  = \4389(1405) ,
  \309(3275)  = ~\4728(2412)  | ~\4721(3217) ,
  \5347(1750)  = ~\5345(1429)  | ~\5342(1079) ,
  \342(3330)  = ~\4799(3259)  | ~\4796(2304) ,
  \6626(1297)  = \2186(989) ,
  \3686(838)  = \3635(408)  | \3666(698) ,
  \4013(2236)  = \3856(1966)  & (\3874(1968)  & \3989(1969) ),
  \5722(2044)  = \1598(1817) ,
  \1628(1176)  = ~\5439(484)  | ~\5436(961) ,
  \967(3355)  = ~\4968(3224)  | ~\4967(3288) ,
  \6795(1591)  = ~\6789(1253) ,
  \5559(3440)  = ~\5553(3391) ,
  \2741(2210)  = ~\6056(1948)  | ~\6049(1049) ,
  \2159(793)  = \2137(738)  & \225(148) ,
  \5393(352)  = \1192(251) ,
  \7507(1002)  = \4473(697)  | \4472(760) ,
  \5808(1237)  = ~\5804(958) ,
  \3956(1778)  = ~\6908(1630)  | ~\6901(332) ,
  \7361(1343)  = \4511(1012) ,
  \3995(1486)  = ~\6923(448)  | ~\6920(1276) ,
  \5357(1753)  = ~\5355(1438)  | ~\5352(1088) ,
  \4928(1454)  = ~\4924(1099) ,
  \6290(3262)  = ~\6288(2805)  | ~\6281(3209) ,
  \6745(1376)  = \3828(1035) ,
  \7165(3427)  = ~\7159(3377) ,
  \7216(1300)  = \2167(990) ,
  \6518(558)  = ~\6514(397) ,
  \6455(1337)  = \4169(1009) ,
  \6122(2923)  = ~\6118(2798) ,
  \5226(1100)  = \2933(861) ,
  \5913(348)  = \3713(241) ,
  \664(574)  = ~\657(404) ,
  \6550(1412)  = ~\6546(1057) ,
  \4251(2476)  = \4198(2157) ,
  \5852(2026)  = \1822(1811) ,
  \3955(1481)  = ~\6907(445)  | ~\6904(1296) ,
  \6599(327)  = \4417(217) ,
  \1553(870)  = \757(856)  & \1192(251) ,
  \6686(2570)  = ~\6682(2244) ,
  \5676(2671)  = ~\5672(2418) ,
  \6332(3697)  = \2849(3692)  | \2848(3693) ,
  \4856(2639)  = ~\4852(2352) ,
  \6493(1647)  = ~\6487(1313) ,
  \6478(1604)  = ~\6474(1269) ,
  \302(3342)  = \2014(3274)  & \2005(2824) ,
  \2(313)  = \1(0) ,
  \1327(3071)  = ~\5376(1961)  | ~\5369(2989) ,
  \5688(3040)  = ~\5686(2830)  | ~\5679(2951) ,
  \4169(1009)  = \4144(706)  | \4143(744) ,
  \1287(2544)  = ~\1284(2220) ,
  \7029(3514)  = ~\7023(3493) ,
  \2505(2336)  = \2391(1134)  & \2372(1986) ,
  \4254(2708)  = ~\4251(2476) ,
  \1280(1751)  = ~\5338(1241)  | ~\5331(1080) ,
  \942(2110)  = \805(1844)  & (\868(934)  & \827(1874) ),
  \574(308)  = ~\5(1) ,
  \3314(1967)  = ~\3313(1766)  | ~\3312(1467) ,
  \2850(3083)  = \2812(2995)  & \2808(2917) ,
  \5572(3501)  = ~\5570(2376)  | ~\5563(3481) ,
  \2241(257)  = ~\2239(181) ,
  \757(856)  = \671(424)  & \710(642) ,
  \3996(1782)  = ~\6924(1613)  | ~\6917(335) ,
  \4282(2983)  = ~\4281(2740)  & ~\4280(2872) ,
  \6355(3119)  = ~\6347(3057) ,
  \5125(3234)  = ~\5119(3175) ,
  \4695(767)  = \4675(482)  | \4674(684) ,
  \352(3318)  = \3486(3004)  & \3491(3249) ,
  \2653(1501)  = ~\6023(459)  | ~\6020(1395) ,
  \3445(2254)  = \3335(1113)  & \3314(1967) ,
  \1883(1177)  = ~\5799(485)  | ~\5796(960) ,
  \6541(1282)  = ~\6535(984) ,
  \7089(3515)  = ~\7087(3497)  | ~\7084(2290) ,
  \5793(365)  = \2226(264) ,
  \1221(2222)  = ~\1217(1960) ,
  \6885(329)  = \4412(219) ,
  \7002(3138)  = ~\7000(2763)  | ~\6993(3076) ,
  \3201(1733)  = ~\6549(1215)  | ~\6546(1057) ,
  \6066(3015)  = ~\6064(2924)  | ~\6057(1136) ,
  \3108(1883)  = ~\6493(1647)  | ~\6490(1299) ,
  \990(3685)  = ~\989(3676) ,
  \1535(302)  = ~\18(5) ,
  \4041(2300)  = \3911(1974)  & (\3979(1126)  & (\3932(1975)  & \3957(1977) )),
  \2295(781)  = \2279(739)  & \239(162) ,
  \5077(3601)  = ~\5071(3585) ,
  \7401(1318)  = \4493(998) ,
  \453(596)  = \572(427) ,
  \805(1844)  = ~\804(1562)  | ~\803(1211) ,
  \7557(1651)  = ~\7551(1316) ,
  \4334(1939)  = ~\7407(1654)  | ~\7404(1042) ,
  \6852(2965)  = ~\6848(2851) ,
  \5764(1075)  = \745(853) ,
  \6341(2538)  = ~\7360(2216)  | ~\7353(1954) ,
  \4561(1897)  = ~\7521(1652)  | ~\7518(1322) ,
  \4571(1898)  = ~\7530(1657)  | ~\7523(1323) ,
  \1775(3666)  = ~\5657(3651)  | ~\5654(2054) ,
  \6365(3129)  = ~\6357(3063) ,
  \4457(583)  = \1530(411) ,
  \2765(2324)  = \2629(1133)  & \2600(1984) ,
  \2755(2325)  = \2629(1133)  & (\2589(1981)  & \2600(1984) ),
  \7353(1954)  = ~\7336(1739)  | ~\7335(1742) ,
  \1541(275)  = ~\1496(173)  | ~\4528(206) ,
  \3713(241)  = ~\3711(188) ,
  \2860(3068)  = ~\6346(2884)  | ~\6337(2961) ,
  \3466(2558)  = \3446(2265)  & \3431(2229) ,
  \5908(1394)  = \2335(1044) ,
  \1711(2012)  = \1556(1807)  & (\1573(1810)  & \1687(1813) ),
  \7238(1708)  = ~\7236(1372)  | ~\7229(1037) ,
  \4077(3659)  = ~\7118(2588)  | ~\7111(3644) ,
  \4180(2159)  = ~\4179(1608)  | ~\4178(1872) ,
  \2352(1489)  = ~\5879(451)  | ~\5876(1259) ,
  \1152(1369)  = ~\5237(720)  | ~\5234(918) ,
  \5246(1194)  = ~\5242(917) ,
  \5657(3651)  = ~\5651(3638) ,
  \5667(3650)  = ~\5661(3637) ,
  \1693(1184)  = ~\5463(489)  | ~\5460(967) ,
  \6996(2561)  = ~\4015(2257)  & (~\4014(2241)  & ~\3868(1110) ),
  \5345(1429)  = ~\5339(1074) ,
  \4609(2729)  = ~\4606(2503) ,
  \5485(3213)  = ~\5484(3103)  | ~\5483(3160) ,
  \6015(458)  = ~\6009(345) ,
  \365(3430)  = \[98] ,
  \6765(1365)  = \2320(1025) ,
  \5504(3438)  = ~\5502(2395)  | ~\5495(3392) ,
  \6495(1311)  = \4166(995) ,
  \4354(1943)  = ~\7432(1724)  | ~\7425(1047) ,
  \7099(3572)  = ~\7097(3552)  | ~\7094(2263) ,
  \1238(1727)  = ~\5287(1413)  | ~\5284(1051) ,
  \496(271)  = \2208(175) ,
  \2838(3672)  = ~\6250(2638)  | ~\6243(3664) ,
  \2799(2531)  = \2724(1722)  & (\2676(1994)  & \2701(1995) ),
  \1312(2542)  = \1288(2219)  & (\1221(2222)  & \1230(2221) ),
  \1653(1179)  = ~\5447(487)  | ~\5444(957) ,
  \2062(657)  = \2032(592)  & \124(63) ,
  \6868(1690)  = ~\6864(1352) ,
  \5142(2123)  = \853(1849) ,
  \389(3021)  = ~\4855(2935)  | ~\4852(2352) ,
  \3478(3001)  = ~\3477(2766)  | ~\3476(2903) ,
  \7327(1064)  = \727(848) ,
  \5415(472)  = ~\5409(356) ,
  \913(1027)  = \784(559)  & \765(774) ,
  \3460(2284)  = \3381(1976)  & \3410(1123) ,
  \5372(1759)  = ~\5280(1457)  | ~\5279(1458) ,
  \1803(1152)  = ~\5759(469)  | ~\5756(1086) ,
  \5888(1593)  = ~\5884(1255) ,
  \5985(336)  = \3751(229) ,
  \579(840)  = \581(421)  & \577(631) ,
  \2162(659)  = \2130(593)  & \121(62) ,
  \4936(1834)  = ~\4932(1547) ,
  \6706(933)  = \3676(777) ,
  \6413(1175)  = ~\6407(903) ,
  \5388(2751)  = ~\5368(2541)  | ~\5367(2540) ,
  \3930(1479)  = ~\6899(443)  | ~\6896(1302) ,
  \3508(2138)  = ~\3504(1851) ,
  \5530(2821)  = ~\5526(2662) ,
  \4816(2586)  = ~\4812(2269) ,
  \3211(827)  = ~\6558(556)  | ~\6551(599) ,
  \4082(3687)  = ~\4081(3679) ,
  \4126(692)  = \4094(584)  & \77(36) ,
  \2675(1798)  = ~\6032(1714)  | ~\6025(349) ,
  \2950(865)  = \2905(426)  & \2928(612) ,
  \546(232)  = \3743(193) ,
  \2500(2322)  = \2384(1132)  & \2354(1983) ,
  \6267(2208)  = ~\6261(1944) ,
  \7537(1684)  = ~\7531(1346) ,
  \332(3304)  = ~\4784(2485)  | ~\4777(3235) ,
  \821(929)  = \2946(858)  & \1482(281) ,
  \322(3302)  = ~\4759(3211)  | ~\4756(2139) ,
  \7317(1068)  = \719(850) ,
  \6298(2880)  = ~\6294(2746) ,
  \1780(3674)  = ~\1779(3648)  | ~\1778(3665) ,
  \4312(1256)  = \2073(971)  & \4505(1014) ,
  \1739(2082)  = \1609(1820)  & (\1677(909)  & (\1630(1824)  & \1655(1827) )),
  \7420(1249)  = \2069(968) ,
  \5132(2135)  = \895(1850) ,
  \7547(1680)  = ~\7541(1342) ,
  \1108(1196)  = \1007(773)  & \1019(923) ,
  \3227(1925)  = ~\3223(1698) ,
  \4938(2202)  = ~\4936(1834)  | ~\4929(564) ,
  \7039(3567)  = ~\7033(3548) ,
  \3450(2274)  = \3393(1121)  & (\3353(1972)  & \3365(1973) ),
  \3531(2480)  = ~\3527(2160) ,
  \3459(3196)  = \3365(1973)  & (\3399(1978)  & (\3381(1976)  & (\3417(1979)  & \2580(3145) ))),
  \4946(1837)  = ~\4942(1551) ,
  \6114(2615)  = ~\6110(2318) ,
  \7595(1801)  = ~\7506(1507)  | ~\7505(1511) ,
  \4316(1899)  = ~\7392(1618)  | ~\7385(1324) ,
  \5457(368)  = \2213(268) ,
  \7139(3006)  = ~\7138(2913)  | ~\7137(2780) ,
  \2929(516)  = \2909(417)  & \212(135) ,
  \1086(935)  = \2938(860)  & \1471(283) ,
  \3415(1484)  = ~\6637(447)  | ~\6634(1275) ,
  \777(370)  = \1198(299)  & \1541(275) ,
  \3816(1021)  = \3792(714)  | \3791(795) ,
  \1383(815)  = \1366(528)  | \1365(644) ,
  \5400(1439)  = ~\5396(1084) ,
  \3931(1776)  = ~\6900(1635)  | ~\6893(330) ,
  \3093(2156)  = ~\3092(1888)  | ~\3091(1870) ,
  \4300(2153)  = ~\4299(1912)  | ~\4298(1867) ,
  \706(640)  = \705(543)  | \685(588) ,
  \7128(2587)  = ~\7124(2270) ,
  \7088(2595)  = ~\7084(2290) ,
  \625(534)  = \606(403)  & \165(88) ,
  \5831(2656)  = ~\5825(2383) ,
  \2059(787)  = \2039(737)  & \233(156) ,
  \2290(569)  = \2259(413)  & \29(8) ,
  \1343(575)  = ~\1336(405) ,
  \7118(2588)  = ~\7114(2272) ,
  \5590(2833)  = ~\5588(2672)  | ~\5581(911) ,
  \1792(3707)  = ~\5744(3698)  | ~\5737(3636) ,
  \3768(595)  = \1507(418) ,
  \2518(2353)  = \2448(1142)  & \2420(1992) ,
  \6717(916)  = ~\6711(772) ,
  \4952(1204)  = \887(922) ,
  \5156(2439)  = ~\5152(2098) ,
  \5174(3700)  = ~\5170(3696) ,
  \1248(1730)  = ~\5296(1411)  | ~\5289(1054) ,
  \5533(3037)  = ~\5532(2946)  | ~\5531(2823) ,
  \5295(1409)  = ~\5289(1054) ,
  \6398(1428)  = ~\6394(1073) ,
  \2779(2527)  = \2655(1991)  & (\2724(1722)  & (\2643(1990)  & (\2676(1994)  & \2701(1995) ))),
  \6703(927)  = \3679(776) ,
  \1914(905)  = \1406(817)  & \2220(266) ,
  \5270(1446)  = ~\5266(1091) ,
  \2548(2922)  = ~\5959(2797)  | ~\5956(2316) ,
  \5383(3066)  = ~\5377(2988) ,
  \1311(2753)  = \1291(2543)  & (\1230(2221)  & \1217(1960) ),
  \6060(2799)  = \2804(2327)  | \2768(2619) ,
  \6908(1630)  = ~\6904(1296) ,
  \4629(2730)  = \4606(2503)  & (\4554(1900)  & \4563(2184) ),
  \2715(1145)  = \2323(1038)  & \3707(243) ,
  \7078(2600)  = ~\7074(2306) ,
  \1357(589)  = ~\1350(415) ,
  \5815(491)  = ~\5809(369) ,
  \2372(1986)  = ~\2371(1788)  | ~\2370(1492) ,
  \6222(3521)  = ~\6220(2646)  | ~\6213(3510) ,
  \4876(401)  = \1198(299) ,
  \6907(445)  = ~\6901(332) ,
  \2920(615)  = \2919(518)  | \2899(590) ,
  \6880(1361)  = \3816(1021) ,
  \1304(2147)  = \1281(1859) ,
  \6226(2347)  = \2643(1990) ,
  \4473(697)  = \4444(582)  & \70(31) ,
  \3416(1781)  = ~\6638(1612)  | ~\6631(334) ,
  \482(253)  = \2253(183) ,
  \4784(2485)  = ~\4780(2168) ,
  \3591(2490)  = \3568(2172) ,
  \3259(2874)  = \3258(2546)  | \3223(1698) ,
  \6743(1693)  = ~\6737(1360) ,
  \2529(2548)  = \2454(1996)  & (\2472(2532)  & \4526(205) ),
  \3350(2261)  = ~\3344(1970) ,
  \3651(509)  = \3622(407)  & \1464(285) ,
  \2862(3185)  = ~\6355(3119)  | ~\6352(2734) ,
  \4535(2093)  = ~\4531(1830) ,
  \6551(599)  = \2872(430) ,
  \7416(1386)  = ~\7412(1039) ,
  \5003(920)  = \765(774) ,
  \3513(1848)  = ~\3512(1616)  | ~\3511(1567) ,
  \4796(2304)  = \3417(1979) ,
  \2806(2755)  = ~\4526(205)  | ~\2771(2634) ,
  \532(218)  = \4415(200) ,
  \384(3016)  = \2406(2344)  & \2564(2929) ,
  \6307(3509)  = ~\6301(3490) ,
  \1686(1522)  = ~\5456(1432)  | ~\5449(359) ,
  \4107(585)  = \1530(411) ,
  \7246(1355)  = ~\7242(1018) ,
  \3117(1930)  = ~\6501(1645)  | ~\6498(1032) ,
  \1134(2131)  = \1038(1843)  & (\1102(940)  & (\1055(1875)  & \1074(1846) )),
  \357(3376)  = ~\4807(3321)  | ~\4804(2266) ,
  \5887(454)  = ~\5881(341) ,
  \5976(2623)  = ~\5972(2331) ,
  \6097(3498)  = ~\6096(3460)  | ~\6095(3478) ,
  \4226(1854)  = ~\4225(1225)  | ~\4224(1574) ,
  \3790(551)  = \3755(412)  & \66(29) ,
  \7522(1660)  = ~\7518(1322) ,
  \4692(768)  = \4673(483)  | \4672(685) ,
  \6264(2640)  = ~\2799(2531)  & (~\2798(2367)  & ~\2693(1143) ),
  \2536(2789)  = \2487(2312)  & \2515(2628) ,
  \6383(880)  = \4704(764) ,
  \7526(1320)  = \4496(999) ,
  \7175(3496)  = ~\7169(3476) ,
  \3438(2239)  = \3327(1111)  & \3295(1965) ,
  \3129(2516)  = \3076(1379)  & (\3052(2192)  & \3062(2194) ),
  \764(603)  = ~\4880(566)  | ~\4873(373) ,
  \6351(2505)  = ~\7344(2203)  | ~\7337(1902) ,
  \4087(3695)  = \4072(3202)  & \4082(3687) ,
  \2843(3689)  = ~\2842(3681) ,
  \4769(3242)  = \1140(3176)  | (\1138(2134)  | (\1137(2117)  | \1068(981) )),
  \4056(3005)  = ~\4053(2910) ,
  \4464(733)  = ~\4457(583) ,
  \3068(1353)  = \3810(823)  & \4172(1008) ,
  \244(3033)  = \1146(2431)  & (\1974(2382)  & (\3466(2558)  & \2537(2915) )),
  \2788(2356)  = \2693(1143)  & \2655(1991) ,
  \4879(495)  = ~\4873(373) ,
  \7497(868)  = \4710(762) ,
  \5359(1957)  = ~\5358(1752)  | ~\5357(1753) ,
  \2757(2602)  = \2756(2339)  | (\2755(2325)  | (\2754(2314)  | \2597(1129) )),
  \3008(1539)  = ~\6422(1226)  | ~\6415(907) ,
  \2635(1135)  = \2091(969)  & \3731(235) ,
  \250(3417)  = \3155(3366)  & \3151(2974) ,
  \1805(1806)  = ~\1804(1513)  | ~\1803(1152) ,
  \4921(381)  = \1464(285) ,
  \2514(2523)  = \2420(1992)  & (\2481(1721)  & (\2409(1989)  & (\2436(1993)  & \2454(1996) ))),
  \2881(3339)  = \2868(3308)  & (\4524(3265)  & \4443(3309) ),
  \3781(621)  = \3762(586)  & \193(116) ,
  \7392(1618)  = ~\7388(1283) ,
  \2524(2525)  = \2481(1721)  & (\2436(1993)  & \2454(1996) ),
  \387(2931)  = ~\4848(2631)  | ~\4841(2804) ,
  \5322(955)  = ~\5318(816) ,
  \3821(1034)  = \3794(724)  | \3793(796) ,
  \2989(889)  = \711(852)  & \4698(766) ,
  \6284(2635)  = ~\2794(2528)  & (~\2793(2364)  & (~\2792(2355)  & ~\2670(1141) )),
  \5436(961)  = \1412(818) ,
  \7592(1674)  = ~\7588(1336) ,
  \2808(2917)  = ~\2753(2603)  | ~\2761(2783) ,
  \307(3389)  = \[90] ,
  \7016(2249)  = \3874(1968) ,
  \7049(2781)  = ~\7047(1485)  | ~\7044(2590) ,
  \264(3121)  = \[59] ,
  \4759(3211)  = ~\4753(3158) ,
  \629(844)  = \581(421)  & \616(729) ,
  \4553(1663)  = ~\7514(1326)  | ~\7507(1002) ,
  \2778(2366)  = \2655(1991)  & (\2715(1145)  & (\2643(1990)  & \2676(1994) )),
  \4729(3218)  = \1968(3163)  | (\1966(2089)  | (\1965(2074)  | \1897(900) )),
  \1376(546)  = \1350(415)  & \151(74) ,
  \4558(2189)  = ~\4554(1900) ,
  \1744(2085)  = \1677(909)  & (\1630(1824)  & \1655(1827) ),
  \7189(3588)  = ~\7188(3550)  | ~\7187(3571) ,
  \5040(3232)  = ~\5038(2686)  | ~\5031(3178) ,
  \2798(2367)  = \2715(1145)  & \2676(1994) ,
  \1795(1804)  = ~\1794(1510)  | ~\1793(1149) ,
  \5108(2843)  = ~\5106(2712)  | ~\5099(1218) ,
  \5929(1048)  = \3682(839) ,
  \3149(3182)  = \3148(3059)  | \3147(3116) ,
  \4225(1225)  = ~\7300(946)  | ~\7293(953) ,
  \5339(1074)  = \745(853) ,
  \7236(1372)  = ~\7232(1033) ,
  \4947(2836)  = ~\4945(2743)  | ~\4942(1551) ,
  \6562(1059)  = \629(844) ,
  \6638(1612)  = ~\6634(1275) ,
  \4679(476)  = \4653(410)  & \2241(257) ,
  \3032(2079)  = \2992(1821)  & (\3013(906)  & (\2982(1816)  & \3001(1823) )),
  \330(3411)  = \[82] ,
  \1055(1875)  = ~\1054(1615)  | ~\1053(1280) ,
  \4306(1864)  = ~\7383(1685)  | ~\7380(1257) ,
  \317(3351)  = ~\4751(3284)  | ~\4748(2075) ,
  \7036(2237)  = \3856(1966) ,
  \2848(3693)  = \2833(317)  & \2843(3689) ,
  \5961(2617)  = ~\2507(2337)  & ~\2384(1132) ,
  \3621(3240)  = ~\3620(3117)  | ~\3619(3181) ,
  \7080(3433)  = ~\7078(2600)  | ~\7071(3378) ,
  \5028(2842)  = ~\5024(2689) ,
  \7026(2225)  = \3845(1963) ,
  \2761(2783)  = ~\2757(2602) ,
  \3141(2492)  = \3093(2156)  & (\3114(1298)  & (\3082(2179)  & \3102(2177) )),
  \4614(2495)  = \4595(2178) ,
  \1235(1958)  = ~\1234(1760)  | ~\1233(1754) ,
  \5627(3485)  = ~\5621(3468) ,
  \341(420)  = \[52] ,
  \6522(1063)  = \645(847) ,
  \697(526)  = \657(404)  & \174(97) ,
  \4678(703)  = \4660(581)  & \63(26) ,
  \5349(1083)  = \757(856) ,
  \2700(1799)  = ~\6040(1710)  | ~\6033(350) ,
  \6337(2961)  = ~\4285(2845)  | ~\4288(2846) ,
  \611(573)  = ~\606(403) ,
  \7551(1316)  = \4151(997) ,
  \1121(1552)  = ~\1117(1193) ,
  \2794(2528)  = \2655(1991)  & (\2724(1722)  & (\2676(1994)  & \2701(1995) )),
  \7162(2305)  = \3997(1980) ,
  \5207(549)  = \1477(394) ,
  \350(3421)  = \[101] ,
  \2813(2930)  = \2775(2803)  & \2784(2802) ,
  \1969(2088)  = \1929(910)  & \1903(1826) ,
  \7247(1691)  = ~\7245(1331)  | ~\7242(1018) ,
  \3957(1977)  = ~\3956(1778)  | ~\3955(1481) ,
  \6653(2761)  = ~\6647(2559) ,
  \6812(2204)  = ~\6754(1933)  | ~\6753(1932) ,
  \2807(2648)  = \2701(1995)  & \2742(2533) ,
  \4128(749)  = \4101(734)  & \4402(223) ,
  \5167(3446)  = \994(3407)  | (\993(3406)  | (\992(3404)  | \991(3405) )),
  \6084(2626)  = ~\6080(2343) ,
  \4740(2066)  = \1885(1825) ,
  \5289(1054)  = \637(842) ,
  \4627(2827)  = ~\4626(2404)  & ~\4625(2678) ,
  \2513(2362)  = \2420(1992)  & (\2465(1144)  & (\2409(1989)  & \2436(1993) )),
  \2523(2363)  = \2436(1993)  & \2465(1144) ,
  \3425(1125)  = \2179(977)  & \4396(225) ,
  \6271(3064)  = ~\6270(2986)  | ~\6269(2878) ,
  \3335(1113)  = \4422(215)  & \3821(1034) ,
  \3136(2475)  = \3082(2179)  & (\3093(2156)  & (\3102(2177)  & (\3110(2175)  & \3122(2158) ))),
  \6212(3473)  = ~\6210(2881)  | ~\6203(3437) ,
  \2435(1797)  = ~\5920(1715)  | ~\5913(348) ,
  \2007(3161)  = \3279(3072)  & \1950(2047) ,
  \7437(2373)  = ~\7602(2021)  | ~\7595(1801) ,
  \1655(1827)  = ~\1654(1538)  | ~\1653(1179) ,
  \2153(791)  = \2137(738)  & \227(150) ,
  \7495(1523)  = ~\7493(1155)  | ~\7490(887) ,
  \2453(1800)  = ~\5928(1709)  | ~\5921(351) ,
  \5824(2380)  = ~\5820(2002) ,
  \6094(2620)  = ~\6090(2328) ,
  \402(395)  = \[41] ,
  \1734(2068)  = \1609(1820)  & (\1669(904)  & \1630(1824) ),
  \5137(3447)  = ~\5135(3409)  | ~\5132(2135) ,
  \1724(2069)  = \1609(1820)  & (\1669(904)  & (\1598(1817)  & \1630(1824) )),
  \1695(1829)  = ~\1694(1542)  | ~\1693(1184) ,
  \4150(704)  = \4107(585)  & \62(25) ,
  \2797(2644)  = \2701(1995)  & (\2676(1994)  & \2742(2533) ),
  \2670(1141)  = \2335(1044)  & \3719(239) ,
  \6104(2605)  = ~\6100(2309) ,
  \5155(3547)  = ~\5149(3528) ,
  \3148(3059)  = \4364(2720)  & \4382(2972) ,
  \6928(2770)  = \4051(2247)  | \4017(2569) ,
  \3183(926)  = \645(847)  & \3679(776) ,
  \4114(735)  = ~\4107(585) ,
  \5473(2826)  = ~\5471(1162)  | ~\5468(2665) ,
  \4670(686)  = \4647(580)  & \83(42) ,
  \2448(1142)  = \2329(1041)  & \3713(241) ,
  \4396(225)  = ~\4394(196) ,
  \5126(2685)  = ~\5122(2443) ,
  \7109(3632)  = ~\7107(3607)  | ~\7104(2279) ,
  \7119(3631)  = ~\7195(3606)  | ~\7192(2278) ,
  \3477(2766)  = ~\6662(2564)  | ~\6655(2568) ,
  \6816(2515)  = ~\6812(2204) ,
  \3200(982)  = \637(842)  & \3673(821) ,
  \1939(2017)  = \1834(878)  & (\1795(1804)  & \1805(1806) ),
  \3997(1980)  = ~\3996(1782)  | ~\3995(1486) ,
  \3775(740)  = ~\3768(595) ,
  \4531(1830)  = ~\4530(1185)  | ~\4529(1545) ,
  \4989(2679)  = ~\4987(1549)  | ~\4980(2511) ,
  \751(857)  = \671(424)  & \708(641) ,
  \5695(3219)  = ~\5689(3164) ,
  \4387(2850)  = \4376(2714)  & \4356(2466) ,
  \6052(1725)  = \4389(1405) ,
  \6032(1714)  = ~\6028(1389) ,
  \4263(2142)  = \4244(1856) ,
  \3467(2760)  = \3431(2229)  & \3453(2578) ,
  \7425(1047)  = \3686(838) ,
  \2300(726)  = \2272(594)  & \29(8) ,
  \6000(1597)  = ~\5996(1260) ,
  \2493(2321)  = \2384(1132)  & (\2343(1982)  & \2354(1983) ),
  \5097(3654)  = ~\5091(3639) ,
  \6179(1946)  = ~\6173(1723) ,
  \1314(2749)  = \1295(2537)  & (\1249(1952)  & \1244(2211) ),
  \5876(1259)  = \2105(972) ,
  \3667(779)  = \3651(509)  | \3650(666) ,
  \5087(3655)  = ~\5081(3640) ,
  \4554(1900)  = ~\4553(1663)  | ~\4552(1664) ,
  \1271(1584)  = ~\5330(1235)  | ~\5323(959) ,
  \4684(669)  = \4660(581)  & \110(55) ,
  \7300(946)  = ~\7296(811) ,
  \5384(1953)  = ~\5380(1736) ,
  \1261(1582)  = ~\5321(1244)  | ~\5318(816) ,
  \6023(459)  = ~\6017(346) ,
  \5471(1162)  = ~\5465(885) ,
  \4369(2486)  = \4317(2170)  & (\4327(2186)  & (\4336(2185)  & (\4344(2188)  & \4355(2207) ))),
  \4277(2876)  = \4258(2716)  & (\4212(1937)  & \4207(2198) ),
  \2550(3013)  = ~\2549(2795)  | ~\2548(2922) ,
  \554(240)  = \3717(189) ,
  \1785(3618)  = \1766(3073)  & (\1754(2950)  & \1757(3594) ),
  \6983(1470)  = \3891(1114) ,
  \2175(975)  = \2152(660)  | \2151(809) ,
  \3176(1840)  = ~\3175(1558)  | ~\3174(1738) ,
  \5726(2408)  = ~\5722(2044) ,
  \1954(2060)  = \1897(900)  & (\1859(1818)  & \1869(1819) ),
  \7614(2181)  = ~\7584(1906)  | ~\7583(1891) ,
  \5380(1736)  = ~\5314(1415)  | ~\5313(1416) ,
  \3070(1675)  = ~\6462(1380)  | ~\6455(1337) ,
  \7541(1342)  = \4511(1012) ,
  \5106(2712)  = ~\5102(2481) ,
  \6107(3555)  = ~\6106(3518)  | ~\6105(3535) ,
  \6186(2811)  = \2807(2648)  | \2801(2645) ,
  \2793(2364)  = \2655(1991)  & (\2715(1145)  & \2676(1994) ),
  \6554(396)  = \1210(298) ,
  \3186(1845)  = ~\3185(1563)  | ~\3184(1729) ,
  \3603(2969)  = ~\3602(2711)  & ~\3601(2856) ,
  \988(3652)  = ~\5098(2446)  | ~\5091(3639) ,
  \4857(2810)  = \2529(2548)  | (\2527(2524)  | \2465(1144) ),
  \6133(3204)  = ~\6131(3149)  | ~\6128(2611) ,
  \7054(2779)  = \4052(2292)  | \4048(2594) ,
  \1240(1950)  = ~\1239(1734)  | ~\1238(1727) ,
  \1793(1149)  = ~\5751(467)  | ~\5748(1085) ,
  \4606(2503)  = \4572(2187) ,
  \6442(1006)  = \3813(822) ,
  \4563(2184)  = ~\4562(1895)  | ~\4561(1897) ,
  \4887(500)  = ~\4881(375) ,
  \6828(2701)  = ~\6826(2467)  | ~\6819(2152) ,
  \2213(268)  = ~\2211(176) ,
  \2809(2893)  = \2806(2755)  & \2784(2802) ,
  \4630(2977)  = ~\4629(2730)  & ~\4628(2865) ,
  \4121(228)  = ~\4393(195) ,
  \1885(1825)  = ~\1884(1536)  | ~\1883(1177) ,
  \5404(1087)  = \751(857) ,
  \7265(1285)  = \2065(985) ,
  \4525(862)  = \2886(425)  & \2918(736) ,
  \5993(339)  = \3745(231) ,
  \5737(3636)  = \1785(3618)  | (\1784(3617)  | (\1783(3615)  | \1782(3616) )),
  \6453(1673)  = ~\6447(1335) ,
  \7531(1346)  = \4505(1014) ,
  \4259(2487)  = \4221(2171) ,
  \1821(1518)  = ~\5768(1430)  | ~\5761(357) ,
  \412(3369)  = \[69] ,
  \3582(2705)  = ~\3579(2473) ,
  \1949(2036)  = \1841(883)  & \1822(1811) ,
  \5935(1402)  = ~\5929(1048) ,
  \6755(1328)  = \3838(1004) ,
  \6932(2905)  = ~\6928(2770) ,
  \1153(1700)  = ~\5238(1195)  | ~\5231(561) ,
  \6118(2798)  = ~\2768(2619) ,
  \6799(1289)  = \2111(987) ,
  \5423(478)  = ~\5417(360) ,
  \6629(446)  = ~\6623(333) ,
  \4489(709)  = \4457(583)  & \56(19) ,
  \4990(2953)  = ~\4989(2679)  | ~\4988(2834) ,
  \7205(1273)  = \2163(976) ,
  \6714(775)  = \3661(496)  | \3660(608) ,
  \1897(900)  = \1412(818)  & \2226(264) ,
  \2980(1748)  = ~\6397(1167)  | ~\6394(1073) ,
  \1488(279)  = ~\1486(171) ,
  \628(637)  = \627(535)  | \611(573) ,
  \2047(802)  = \2026(730)  & \203(126) ,
  \5284(1051)  = ~\579(840) ,
  \7478(1181)  = ~\7474(908) ,
  \7369(1344)  = \4508(1013) ,
  \7367(1681)  = ~\7361(1343) ,
  \7006(2259)  = \3989(1969) ,
  \7409(1321)  = \4490(1000) ,
  \3932(1975)  = ~\3931(1776)  | ~\3930(1479) ,
  \5047(3410)  = ~\5041(3360) ,
  \5863(1520)  = ~\5857(1159) ,
  \3536(2174)  = ~\3535(1885)  | ~\3534(1882) ,
  \1207(307)  = ~\9(2)  | ~\12(3) ,
  \2147(807)  = \2124(731)  & \196(119) ,
  \6893(330)  = \4407(221) ,
  \394(3095)  = \[63] ,
  \4807(3321)  = ~\4801(3250) ,
  \3410(1123)  = \2186(989)  & \4402(223) ,
  \1391(813)  = \1370(521)  | \1369(646) ,
  \6642(2227)  = \3283(1964) ,
  \490(263)  = \2230(179) ,
  \6752(1702)  = ~\6748(1373) ,
  \5321(1244)  = ~\5315(965) ,
  \410(387)  = \[45] ,
  \3602(2711)  = \3579(2473)  & (\3527(2160)  & \3536(2174) ),
  \1210(298)  = \38(11) ,
  \5162(2166)  = \827(1874) ,
  \2048(653)  = \2019(576)  & \130(65) ,
  \5146(2452)  = ~\5142(2123) ,
  \5136(2453)  = ~\5132(2135) ,
  \1630(1824)  = ~\1629(1535)  | ~\1628(1176) ,
  \5735(3596)  = ~\5729(3582) ,
  \4057(3586)  = ~\6981(3568)  | ~\6978(2235) ,
  \6236(2360)  = \2676(1994) ,
  \4719(3192)  = ~\4713(3136) ,
  \5996(1260)  = \2105(972) ,
  \540(227)  = \4393(195) ,
  \6202(3336)  = ~\6200(2933)  | ~\6193(3263) ,
  \5669(1182)  = \1677(909) ,
  \3629(578)  = ~\3622(407) ,
  \6789(1253)  = \2099(970) ,
  \5057(3489)  = ~\5051(3471) ,
  \6965(3492)  = ~\6964(3454)  | ~\6963(3474) ,
  \4211(1716)  = ~\7264(1387)  | ~\7257(1043) ,
  \5229(510)  = ~\5223(382) ,
  \6317(3558)  = ~\6311(3537) ,
  \1158(1927)  = ~\1157(1699)  | ~\1156(1368) ,
  \886(604)  = ~\4920(565)  | ~\4913(497) ,
  \715(851)  = \650(423)  & \694(627) ,
  \4959(3170)  = ~\4958(3048)  | ~\4957(3112) ,
  \6216(2369)  = \2701(1995) ,
  \6639(2560)  = \3440(2234)  | (\3439(2252)  | (\3438(2239)  | \3308(1109) )),
  \5895(456)  = ~\5889(343) ,
  \2923(513)  = \2892(416)  & \215(138) ,
  \1316(2882)  = ~\1315(2534)  & ~\1314(2749) ,
  \4481(696)  = \4457(583)  & \73(32) ,
  \1023(1205)  = ~\1019(923) ,
  \1647(899)  = \1412(818)  & \2226(264) ,
  \868(934)  = \2938(860)  & \1471(283) ,
  \7407(1654)  = ~\7401(1318) ,
  \6246(2351)  = \2655(1991) ,
  \7601(1997)  = ~\7595(1801) ,
  \5230(1455)  = ~\5226(1100) ,
  \6570(1329)  = \3838(1004) ,
  \5280(1457)  = ~\5278(1103)  | ~\5271(863) ,
  \1381(651)  = \1357(589)  & \135(68) ,
  \6915(437)  = ~\6909(324) ,
  \6256(2350)  = \2655(1991) ,
  \257(2860)  = \3249(2223)  & (\3035(2374)  & (\3156(2706)  & (\4386(2698)  & \89(48) ))),
  \2470(1945)  = ~\5935(1402)  | ~\5932(1726) ,
  \6145(3434)  = ~\6144(3333)  | ~\6143(3383) ,
  \5760(1441)  = ~\5756(1086) ,
  \6682(2244)  = \3314(1967) ,
  \1370(521)  = \1336(405)  & \179(102) ,
  \3607(2875)  = \3590(2717)  & (\3559(2205)  & \3554(2510) ),
  \5610(3216)  = ~\5608(2670)  | ~\5601(3166) ,
  \7177(3516)  = ~\7175(3496)  | ~\7172(2291) ,
  \3458(2294)  = \3365(1973)  & (\3425(1125)  & (\3381(1976)  & \3399(1978) )),
  \700(630)  = \699(527)  | \664(574) ,
  \3800(700)  = \3768(595)  & \66(29) ,
  \6124(3014)  = ~\6122(2923)  | ~\6115(1494) ,
  \2186(989)  = \2158(677)  | \2157(792) ,
  \2655(1991)  = ~\2654(1795)  | ~\2653(1501) ,
  \1440(3030)  = \1788(2375)  & (\4089(2553)  & \2854(2916) ),
  \4284(2456)  = \4263(2142)  & (\4226(1854)  & \4235(1855) ),
  \7380(1257)  = \2073(971) ,
  \4198(2157)  = ~\4197(1921)  | ~\4196(1605) ,
  \2039(737)  = ~\2032(592) ,
  \4157(1010)  = \4132(707)  | \4131(748) ,
  \5864(2397)  = ~\5860(2025) ,
  \5070(3545)  = ~\5068(2440)  | ~\5061(3527) ,
  \1709(2016)  = \1584(877)  & \1556(1807) ,
  \5444(957)  = \1406(817) ,
  \6904(1296)  = \2186(989) ,
  \5951(2790)  = ~\5945(2609) ,
  \5820(2002)  = \1795(1804) ,
  \3648(665)  = \3629(578)  & \114(59) ,
  \2148(678)  = \2117(577)  & \97(50) ,
  \5839(2664)  = ~\5833(2393) ,
  \3147(3116)  = \4385(3060)  & \4381(2964) ,
  \4727(3278)  = ~\4721(3217) ,
  \4929(564)  = ~\1198(299)  & ~\1519(374) ,
  \2238(259)  = ~\2236(180) ,
  \5589(2677)  = ~\5587(1183)  | ~\5584(2419) ,
  \4996(3045)  = ~\4990(2953) ,
  \5385(2962)  = ~\1322(2847)  | ~\1325(2848) ,
  \5660(3598)  = ~\5736(2421)  | ~\5729(3582) ,
  \5650(3599)  = ~\5648(2422)  | ~\5641(3583) ,
  \3184(1729)  = ~\6533(1212)  | ~\6530(1053) ,
  \3417(1979)  = ~\3416(1781)  | ~\3415(1484) ,
  \6748(1373)  = \3821(1034) ,
  \3843(1463)  = ~\6859(431)  | ~\6856(1327) ,
  \2111(987)  = \2064(675)  | \2063(789) ,
  \6818(2732)  = ~\6816(2515)  | ~\6809(2190) ,
  \3025(2005)  = \2970(872)  & \2956(1802) ,
  \1749(2022)  = \1573(1810)  & \1687(1813) ,
  \637(842)  = \581(421)  & \620(633) ,
  \4184(2479)  = ~\4180(2159) ,
  \1499(273)  = ~\1496(173) ,
  \7431(1401)  = ~\7425(1047) ,
  \5401(355)  = \1186(254) ,
  \5011(941)  = ~\2933(861)  & ~\1464(285) ,
  \7067(3256)  = ~\7061(3199) ,
  \2600(1984)  = ~\2599(1786)  | ~\2598(1490) ,
  \5736(2421)  = ~\5732(2063) ,
  \5408(1442)  = ~\5404(1087) ,
  \6020(1395)  = \2335(1044) ,
  \3464(3200)  = \3399(1978)  & (\3417(1979)  & \2580(3145) ),
  \6578(1350)  = \3833(1016) ,
  \6470(1357)  = ~\6466(1019) ,
  \723(849)  = \650(423)  & \698(629) ,
  \2522(2550)  = \2420(1992)  & (\2454(1996)  & (\2436(1993)  & (\2472(2532)  & \4526(205) ))),
  \2578(3082)  = \2571(3018)  & \2495(2601) ,
  \962(2839)  = \924(2441)  & \933(2683) ,
  \5706(2428)  = ~\5702(2090) ,
  \3762(586)  = ~\3755(412) ,
  \3579(2473)  = \3545(2155) ,
  \7260(1040)  = \2308(835) ,
  \5166(2483)  = ~\5162(2166) ,
  \7090(3494)  = ~\7088(2595)  | ~\7081(3477) ,
  \5716(2427)  = ~\5712(2077) ,
  \594(572)  = ~\587(402) ,
  \372(2890)  = ~\4840(2879)  | ~\4833(207) ,
  \3174(1738)  = ~\6525(1207)  | ~\6522(1063) ,
  \1880(895)  = \1418(819)  & \2232(262) ,
  \1850(1812)  = ~\1849(1521)  | ~\1848(1160) ,
  \4581(2500)  = ~\4577(2183) ,
  \3557(1935)  = ~\6779(1713)  | ~\6776(1384) ,
  \2818(3575)  = ~\6114(2615)  | ~\6107(3555) ,
  \4308(2151)  = ~\4307(1915)  | ~\4306(1864) ,
  \4855(2935)  = ~\4849(2807) ,
  \4788(2118)  = \1074(1846) ,
  \3844(1762)  = ~\6860(1665)  | ~\6853(318) ,
  \440(277)  = \1492(172) ,
  \6607(328)  = \4412(219) ,
  \3021(1831)  = ~\3020(1543)  | ~\3019(1581) ,
  \4744(2423)  = ~\4740(2066) ,
  \851(1217)  = ~\4911(507)  | ~\4908(1096) ,
  \4516(3024)  = ~\7442(2814)  | ~\7433(2949) ,
  \1233(1754)  = ~\5269(1459)  | ~\5266(1091) ,
  \305(3343)  = \2014(3274)  & \1850(1812) ,
  \4216(2206)  = ~\4212(1937) ,
  \5801(366)  = \2220(266) ,
  \5896(1588)  = ~\5892(1250) ,
  \5964(2315)  = \2354(1983) ,
  \4673(483)  = \4640(409)  & \2226(264) ,
  \4272(2710)  = \4247(2477)  & (\4180(2159)  & \4189(2176) ),
  \4062(3587)  = ~\7039(3567)  | ~\7036(2237) ,
  \6176(2809)  = \2797(2644)  | (\2796(2529)  | (\2795(2368)  | \2693(1143) )),
  \1714(2031)  = \1590(882)  & \1573(1810) ,
  \7336(1739)  = ~\7334(1422)  | ~\7327(1064) ,
  \6193(3263)  = ~\6192(3154)  | ~\6191(3208) ,
  \6196(2806)  = \2791(2637)  | (\2790(2526)  | (\2789(2365)  | (\2788(2356)  | \2670(1141) ))),
  \6414(1229)  = ~\6410(950) ,
  \6711(772)  = \3663(493)  | \3662(601) ,
  \2308(835)  = \2290(569)  | \2289(617) ,
  \2303(784)  = \2279(739)  & \236(159) ,
  \2472(2532)  = ~\2471(2209)  | ~\2470(1945) ,
  \4262(2715)  = ~\4259(2487) ,
  \4817(3254)  = \3464(3200)  | (\3463(2296)  | \3410(1123) ),
  \5215(379)  = \1471(283) ,
  \5598(2831)  = ~\5594(2675) ,
  \7326(1743)  = ~\7324(1426)  | ~\7317(1068) ,
  \6634(1275)  = \2179(977) ,
  \6391(891)  = \4698(766) ,
  \355(3317)  = \3350(2261)  & \3491(3249) ,
  \2259(413)  = \1535(302) ,
  \6486(1637)  = ~\6482(1304) ,
  \5759(469)  = ~\5753(354) ,
  \852(1568)  = ~\4912(1451)  | ~\4905(380) ,
  \3001(1823)  = ~\3000(1534)  | ~\2999(1578) ,
  \6048(1589)  = ~\6044(1251) ,
  \5128(3231)  = ~\5126(2685)  | ~\5119(3175) ,
  \3034(2403)  = \3033(2092)  | (\3032(2079)  | (\3031(2061)  | (\3030(2055)  | \2989(889) ))),
  \7438(2650)  = ~\7437(2373)  | ~\7436(2394) ,
  \7505(1511)  = ~\7503(1146)  | ~\7500(873) ,
  \1596(1168)  = ~\5423(478)  | ~\5420(1082) ,
  \7583(1891)  = ~\7581(1677)  | ~\7578(1312) ,
  \7582(1646)  = ~\7578(1312) ,
  \2784(2802)  = ~\2780(2629) ,
  \3463(2296)  = \3425(1125)  & \3399(1978) ,
  \6758(1351)  = \3833(1016) ,
  \5707(3442)  = ~\5705(3394)  | ~\5702(2090) ,
  \7168(3432)  = ~\7166(2599)  | ~\7159(3377) ,
  \1284(2220)  = \1235(1958) ,
  \7176(2596)  = ~\7172(2291) ,
  \7166(2599)  = ~\7162(2305) ,
  \2161(794)  = \2137(738)  & \224(147) ,
  \4085(3629)  = \4067(3144)  & (\4053(2910)  & \4064(3605) ),
  \4478(757)  = \4451(732)  & \3719(239) ,
  \5483(3160)  = ~\5481(3105)  | ~\5478(2388) ,
  \5920(1715)  = ~\5916(1390) ,
  \5678(2832)  = ~\5676(2671)  | ~\5669(1182) ,
  \7208(978)  = \2144(663)  | \2143(806) ,
  \6232(3578)  = ~\6230(2633)  | ~\6223(3557) ,
  \5181(494)  = ~\5175(372) ,
  \3118(1644)  = ~\6502(1371)  | ~\6495(1311) ,
  \5705(3394)  = ~\5699(3347) ,
  \4748(2075)  = \1903(1826) ,
  \4011(2243)  = \3885(1112)  & \3856(1966) ,
  \4051(2247)  = \3874(1968)  & \3989(1969) ,
  \4343(1658)  = ~\7416(1386)  | ~\7409(1321) ,
  \7356(1955)  = ~\7326(1743)  | ~\7325(1746) ,
  \6654(2557)  = ~\6650(2228) ,
  \1315(2534)  = \1292(2213)  & (\1240(1950)  & \1249(1952) ),
  \2973(1808)  = ~\2972(1515)  | ~\2971(1744) ,
  \3155(3366)  = ~\3152(3305) ,
  \5725(3543)  = ~\5719(3526) ,
  \4026(2287)  = \3911(1974)  & (\3971(1124)  & (\3899(1971)  & \3932(1975) )),
  \945(2128)  = \877(939)  & (\827(1874)  & \853(1849) ),
  \1471(283)  = ~\1469(169) ,
  \1244(2211)  = ~\1240(1950) ,
  \262(2993)  = \3249(2223)  & (\3035(2374)  & (\3156(2706)  & \4388(2971) )),
  \691(523)  = \657(404)  & \177(100) ,
  \4036(2286)  = \3911(1974)  & (\3971(1124)  & \3932(1975) ),
  \6822(2150)  = ~\6798(1863)  | ~\6797(1862) ,
  \7308(1227)  = ~\7304(948) ,
  \6719(1202)  = ~\6717(916)  | ~\6714(775) ,
  \7196(2591)  = ~\7192(2278) ,
  \2249(255)  = ~\2247(182) ,
  \2210(270)  = ~\2208(175) ,
  \5816(1245)  = ~\5812(966) ,
  \1778(3665)  = ~\5667(3650)  | ~\5664(2052) ,
  \2763(2338)  = \2600(1984)  & (\2635(1135)  & \2618(1985) ),
  \368(3431)  = \[99] ,
  \6031(462)  = ~\6025(349) ,
  \2588(1783)  = ~\5992(1625)  | ~\5985(336) ,
  \4594(1890)  = ~\7574(1640)  | ~\7567(1310) ,
  \4584(1893)  = ~\7565(1679)  | ~\7562(1314) ,
  \2933(861)  = \2886(425)  & \2920(615) ,
  \4197(1921)  = ~\7228(1606)  | ~\7221(1020) ,
  \7493(1155)  = ~\7487(881) ,
  \7503(1146)  = ~\7497(868) ,
  \418(3449)  = \[85] ,
  \3121(1894)  = ~\6510(1607)  | ~\6503(1315) ,
  \1038(1843)  = ~\1037(1561)  | ~\1036(1210) ,
  \4072(3202)  = ~\4067(3144) ,
  \4865(2877)  = \2531(2547)  | \2481(1721) ,
  \6063(1495)  = ~\6057(1136) ,
  \374(3152)  = \2571(3018)  & \2547(3084) ,
  \6709(1206)  = ~\6703(927) ,
  \4307(1915)  = ~\7384(1594)  | ~\7377(1347) ,
  \6943(3194)  = ~\6941(3141)  | ~\6938(2562) ,
  \321(3715)  = \[104] ,
  \912(1550)  = ~\908(1192) ,
  \4519(3124)  = ~\7452(2975)  | ~\7443(3061) ,
  \6573(432)  = ~\6567(319) ,
  \5969(1137)  = ~\3731(235)  & ~\2091(969) ,
  \1751(2828)  = \1721(2410)  & \1730(2668) ,
  \2892(416)  = \1503(303) ,
  \297(3266)  = \1987(2942)  & \2008(3214) ,
  \3575(2095)  = \3522(1839) ,
  \5594(2675)  = \1750(2078)  | \1746(2424) ,
  \4767(3297)  = ~\4761(3233) ,
  \2503(2323)  = \2384(1132)  & \2354(1983) ,
  \7598(1809)  = ~\7496(1516)  | ~\7495(1523) ,
  \916(1030)  = \784(559)  & \765(774) ,
  \6155(3499)  = ~\6154(3461)  | ~\6153(3479) ,
  \2981(1526)  = ~\6398(1428)  | ~\6391(891) ,
  \1944(2009)  = \1805(1806)  & (\1822(1811)  & \1850(1812) ),
  \1145(3179)  = \1093(1853)  & \3271(3101) ,
  \3554(2510)  = ~\3550(2199) ,
  \4864(2641)  = ~\4860(2358) ,
  \3277(2891)  = \3466(2558)  & (\2532(2788)  & \4526(205) ),
  \335(3300)  = ~\4792(2449)  | ~\4785(3237) ,
  \6335(3656)  = ~\6329(3641) ,
  \267(3027)  = \997(2432)  & (\1788(2375)  & \4091(2899) ),
  \5515(3539)  = ~\5514(3502)  | ~\5513(3524) ,
  \6773(1388)  = \2329(1041) ,
  \2305(826)  = \2288(555)  | \2287(620) ,
  \6764(1901)  = ~\6762(1689)  | ~\6755(1328) ,
  \4689(769)  = \4671(488)  | \4670(686) ,
  \1571(1156)  = ~\5415(472)  | ~\5412(1076) ,
  \2370(1492)  = ~\5887(454)  | ~\5884(1255) ,
  \3091(1870)  = ~\6477(1639)  | ~\6474(1269) ,
  \1006(602)  = ~\5182(563)  | ~\5175(372) ,
  \1941(2379)  = \1940(2032)  | (\1939(2017)  | (\1938(2006)  | \1802(871) )),
  \4483(712)  = \4457(583)  & \53(16) ,
  \4305(1262)  = \2077(973)  & \4508(1013) ,
  \3231(2109)  = \3192(931)  & \3176(1840) ,
  \4895(503)  = ~\4889(378) ,
  \2156(662)  = \2130(593)  & \118(61) ,
  \4285(2845)  = ~\4284(2456)  & ~\4283(2694) ,
  \6065(2927)  = ~\6063(1495)  | ~\6060(2799) ,
  \4967(3288)  = ~\4965(3227)  | ~\4962(919) ,
  \1127(2116)  = \1038(1843)  & (\1086(935)  & (\1026(1842)  & \1055(1875) )),
  \6637(447)  = ~\6631(334) ,
  \5288(1406)  = ~\5284(1051) ,
  \2823(3576)  = ~\6172(2616)  | ~\6165(3554) ,
  \6095(3478)  = ~\6093(3463)  | ~\6090(2328) ,
  \2641(1500)  = ~\6015(458)  | ~\6012(1287) ,
  \1137(2117)  = \1055(1875)  & \1086(935) ,
  \5194(1106)  = \2950(865) ,
  \7447(2735)  = ~\7618(2498)  | ~\7611(2193) ,
  \7457(2736)  = ~\7610(2508)  | ~\7603(2196) ,
  \3885(1112)  = \3828(1035)  & \4429(213) ,
  \2155(800)  = \2137(738)  & \217(140) ,
  \3022(1998)  = \2956(1802)  & (\2965(1805)  & (\2973(1808)  & \3018(1814) )),
  \6685(1768)  = ~\6679(1469) ,
  \6606(1692)  = ~\6602(1359) ,
  \5860(2025)  = \1822(1811) ,
  \4016(2258)  = \3891(1114)  & \3874(1968) ,
  \5772(1078)  = \737(854) ,
  \1295(2537)  = ~\1292(2213) ,
  \4348(1385)  = \2308(835)  & \4490(1000) ,
  \1053(1280)  = ~\5213(672)  | ~\5210(1094) ,
  \4549(1815)  = ~\4548(1525)  | ~\4547(1532) ,
  \6549(1215)  = ~\6543(937) ,
  \5431(481)  = ~\5425(363) ,
  \6955(3423)  = ~\6954(3316)  | ~\6953(3374) ,
  \6180(2936)  = ~\6176(2809) ,
  \3443(2253)  = \3335(1113)  & \3314(1967) ,
  \242(2955)  = \1146(2431)  & \1982(2816) ,
  \1116(1031)  = \1014(560)  & \1007(773) ,
  \2991(1531)  = ~\6406(1230)  | ~\6399(897) ,
  \6183(3131)  = ~\6182(3065)  | ~\6181(2987) ,
  \2909(417)  = \1503(303) ,
  \6190(2939)  = ~\6186(2811) ,
  \853(1849)  = ~\852(1568)  | ~\851(1217) ,
  \3707(243)  = ~\3705(187) ,
  \5367(2540)  = ~\5365(2218)  | ~\5362(1956) ,
  \1303(2462)  = ~\1300(2146) ,
  \5303(1417)  = ~\5297(1062) ,
  \2003(2399)  = ~\5863(1520)  | ~\5860(2025) ,
  \6016(1622)  = ~\6012(1287) ,
  \2865(3180)  = ~\6365(3129)  | ~\6362(2849) ,
  \737(854)  = \671(424)  & \704(639) ,
  \7359(2215)  = ~\7353(1954) ,
  \5313(1416)  = ~\5311(1060)  | ~\5308(846) ,
  \4407(221)  = ~\4405(198) ,
  \5488(2039)  = \1687(1813) ,
  \[100]  = \346(3311)  | \345(3370) ,
  \4342(1936)  = ~\7415(1659)  | ~\7412(1039) ,
  \[101]  = \349(3314)  | \348(3371) ,
  \[102]  = \352(3318)  | \351(3372) ,
  \1256(1728)  = ~\5303(1417)  | ~\5300(1052) ,
  \6923(448)  = ~\6917(335) ,
  \[103]  = \355(3317)  | \354(3375) ,
  \[104]  = ~\320(3711) ,
  \4617(2722)  = ~\4614(2495) ,
  \6346(2884)  = ~\6342(2750) ,
  \[105]  = ~\337(3712) ,
  \[106]  = ~\369(3714) ,
  \6200(2933)  = ~\6196(2806) ,
  \5562(3439)  = ~\5560(2396)  | ~\5553(3391) ,
  \5916(1390)  = \2329(1041) ,
  \2931(517)  = \2909(417)  & \211(134) ,
  \[107]  = ~\398(3713) ,
  \5231(561)  = ~\1519(374)  & ~\1198(299) ,
  \1019(923)  = ~\1018(606)  | ~\1017(831) ,
  \4576(1650)  = ~\7558(1341)  | ~\7551(1316) ,
  \1754(2950)  = ~\1751(2828) ,
  \1482(281)  = ~\1480(170) ,
  \2495(2601)  = \2494(2333)  | (\2493(2321)  | (\2492(2313)  | \2351(1128) )),
  \2549(2795)  = ~\5960(2614)  | ~\5953(2618) ,
  \2061(788)  = \2039(737)  & \232(155) ,
  \1267(2144)  = ~\1263(1857) ,
  \5495(3392)  = ~\5494(3273)  | ~\5493(3345) ,
  \6421(1180)  = ~\6415(907) ,
  \5008(3289)  = ~\5006(3226)  | ~\5003(920) ,
  \6463(1309)  = \4163(994) ,
  \622(634)  = \621(532)  | \594(572) ,
  \6761(1666)  = ~\6755(1328) ,
  \1002(2682)  = \929(2433)  & \902(1199) ,
  \7565(1679)  = ~\7559(1340) ,
  \925(2103)  = \821(929)  & \792(1841) ,
  \6754(1933)  = ~\6752(1702)  | ~\6745(1376) ,
  \6105(3535)  = ~\6103(3519)  | ~\6100(2309) ,
  \7178(3495)  = ~\7176(2596)  | ~\7169(3476) ,
  \5239(719)  = \1014(560) ,
  \2329(1041)  = \2302(727)  | \2301(783) ,
  \2558(3017)  = ~\2557(2928) ,
  \6028(1389)  = \2329(1041) ,
  \1849(1521)  = ~\5776(1433)  | ~\5769(358) ,
  \5865(337)  = \3751(229) ,
  \2928(612)  = \2927(515)  | \2914(591) ,
  \2527(2524)  = \2481(1721)  & \2454(1996) ,
  \5498(2023)  = \1573(1810) ,
  \4333(1397)  = \2316(837)  & \4496(999) ,
  \3656(667)  = \3629(578)  & \112(57) ,
  \6008(1592)  = ~\6004(1254) ,
  \619(531)  = \587(402)  & \168(91) ,
  \6671(1116)  = ~\4422(215)  & ~\3821(1034) ,
  \7280(1586)  = ~\7276(1247) ,
  \3486(3004)  = ~\3485(2909) ,
  \5640(3541)  = ~\5638(2409)  | ~\5631(3525) ,
  \7510(1003)  = \4471(699)  | \4470(761) ,
  \2420(1992)  = ~\2419(1796)  | ~\2418(1502) ,
  \4289(1880)  = ~\7367(1681)  | ~\7364(1292) ,
  \2289(617)  = \2266(587)  & \207(130) ,
  \6694(945)  = ~\6690(780) ,
  \2056(674)  = \2032(592)  & \103(52) ,
  \2232(262)  = ~\2230(179) ,
  \4032(2773)  = ~\4028(2579) ,
  \4840(2879)  = ~\4836(2745) ,
  \1279(1585)  = ~\5337(1435)  | ~\5334(962) ,
  \705(543)  = \678(414)  & \155(78) ,
  \645(847)  = \601(422)  & \624(635) ,
  \7462(2981)  = ~\7458(2870) ,
  \1160(3173)  = \3271(3101)  & \1122(2101) ,
  \1629(1535)  = ~\5440(1240)  | ~\5433(364) ,
  \1140(3176)  = \1074(1846)  & (\1055(1875)  & (\1093(1853)  & \3271(3101) )),
  \279(304)  = \[37] ,
  \6172(2616)  = ~\6168(2320) ,
  \6356(2869)  = ~\6352(2734) ,
  \312(3279)  = ~\4736(2415)  | ~\4729(3218) ,
  \3363(1477)  = ~\6613(441)  | ~\6610(1266) ,
  \6618(1303)  = \2192(991) ,
  \1669(904)  = \1406(817)  & \2220(266) ,
  \3076(1379)  = \3807(834)  & \4169(1009) ,
  \4147(705)  = \4107(585)  & \61(24) ,
  \7559(1340)  = \4157(1010) ,
  \7186(2580)  = ~\7182(2262) ,
  \6044(1251)  = \2091(969) ,
  \6004(1254)  = \2099(970) ,
  \4172(1008)  = \4147(705)  | \4146(743) ,
  \7013(3422)  = ~\7012(3315)  | ~\7011(3373) ,
  \6314(2346)  = \2643(1990) ,
  \4212(1937)  = ~\4211(1716)  | ~\4210(1712) ,
  \7097(3552)  = ~\7091(3532) ,
  \6381(1151)  = ~\6375(874) ,
  \333(3416)  = \[83] ,
  \1258(1951)  = ~\1257(1737)  | ~\1256(1728) ,
  \7320(1071)  = \715(851) ,
  \2857(293)  = \240(163)  & (\228(151)  & (\184(107)  & \150(73) )),
  \5391(3055)  = ~\5385(2962) ,
  \4374(2518)  = \4327(2186)  & (\4348(1385)  & (\4317(2170)  & \4336(2185) )),
  \7032(3511)  = ~\7030(2554)  | ~\7023(3493) ,
  \2400(1988)  = ~\2399(1792)  | ~\2398(1497) ,
  \3293(1465)  = ~\6581(433)  | ~\6578(1350) ,
  \2733(1791)  = ~\6048(1589)  | ~\6041(342) ,
  \1367(650)  = \1343(575)  & \138(69) ,
  \6142(2625)  = ~\6138(2342) ,
  \4686(770)  = \4669(490)  | \4668(701) ,
  \7057(3081)  = ~\7051(3007) ,
  \7452(2975)  = ~\7448(2862) ,
  \3794(724)  = \3768(595)  & \35(10) ,
  \2406(2344)  = ~\2400(1988) ,
  \2297(790)  = \2279(739)  & \229(152) ,
  \6808(1879)  = ~\6806(1598)  | ~\6799(1289) ,
  \5024(2689)  = \956(2124)  | \950(2448) ,
  \272(3287)  = \1161(3229)  & \1176(1838) ,
  \1756(3561)  = ~\5522(2389)  | ~\5515(3539) ,
  \4892(1090)  = \2946(858) ,
  \671(424)  = \1207(307) ,
  \446(393)  = \1475(295) ,
  \3659(499)  = \3635(408)  & \1488(279) ,
  \3789(625)  = \3762(586)  & \189(112) ,
  \5348(1749)  = ~\5346(1434)  | ~\5339(1074) ,
  \5090(3602)  = ~\5166(2483)  | ~\5159(3584) ,
  \2408(1793)  = ~\5904(1623)  | ~\5897(344) ,
  \1737(2056)  = \1647(899)  & \1609(1820) ,
  \526(212)  = \4432(203) ,
  \6152(2621)  = ~\6148(2329) ,
  \353(3425)  = \[102] ,
  \5329(1238)  = ~\5323(959) ,
  \3797(798)  = \3775(740)  & \220(143) ,
  \3617(3126)  = ~\6844(2979)  | ~\6837(3056) ,
  \3294(1764)  = ~\6582(1688)  | ~\6575(320) ,
  \3597(2841)  = ~\3596(2450)  & ~\3595(2688) ,
  \6771(1697)  = ~\6765(1365) ,
  \4777(3235)  = \1143(3177)  | (\1141(2133)  | \1086(935) ),
  \5080(3603)  = ~\5078(2484)  | ~\5071(3585) ,
  \3784(567)  = \3755(412)  & \35(10) ,
  \1375(643)  = \1357(589)  & \147(72) ,
  \3139(2474)  = \3099(1268)  & \3082(2179) ,
  \3845(1963)  = ~\3844(1762)  | ~\3843(1463) ,
  \7530(1657)  = ~\7526(1320) ,
  \5817(2384)  = \1944(2009)  | (\1943(2034)  | (\1942(2018)  | \1816(875) )),
  \5247(1098)  = \2933(861) ,
  \4937(1929)  = ~\4935(722)  | ~\4932(1547) ,
  \2740(1947)  = ~\6055(1403)  | ~\6052(1725) ,
  \3364(1774)  = ~\6614(1602)  | ~\6607(328) ,
  \3599(2436)  = \3575(2095)  & (\3508(2138)  & \3517(2120) ),
  \1901(1178)  = ~\5807(486)  | ~\5804(958) ,
  \5984(2622)  = ~\5980(2330) ,
  \4486(753)  = \4464(733)  & \3745(231) ,
  \1884(1536)  = ~\5800(1239)  | ~\5793(365) ,
  \4093(3710)  = ~\7204(3706)  | ~\7197(3642) ,
  \2742(2533)  = ~\2741(2210)  | ~\2740(1947) ,
  \1598(1817)  = ~\1597(1527)  | ~\1596(1168) ,
  \4080(3658)  = ~\7128(2587)  | ~\7121(3643) ,
  \4939(2512)  = ~\4938(2202)  | ~\4937(1929) ,
  \5223(382)  = \1464(285) ,
  \345(3370)  = \3497(3319)  & \3475(3074) ,
  \4125(750)  = \4101(734)  & \4396(225) ,
  \1512(300)  = \18(5) ,
  \4472(760)  = \4451(732)  & \3703(245) ,
  \2091(969)  = \2058(654)  | \2057(786) ,
  \2693(1143)  = \2329(1041)  & \3713(241) ,
  \4681(471)  = \4653(410)  & \2249(255) ,
  \5601(3166)  = ~\5600(3041)  | ~\5599(3107) ,
  \5034(2444)  = \940(2107)  | (\939(2125)  | (\938(2111)  | (\937(2162)  | \821(929) ))),
  \5541(3159)  = ~\5539(3104)  | ~\5536(2387) ,
  \5768(1430)  = ~\5764(1075) ,
  \3521(1557)  = ~\6710(1213)  | ~\6703(927) ,
  \7514(1326)  = ~\7510(1003) ,
  \2543(3009)  = ~\2542(2786)  | ~\2541(2918) ,
  \1146(2431)  = \1122(2101)  & \1108(1196) ,
  \2316(837)  = \2294(571)  | \2293(619) ,
  \4244(1856)  = ~\4243(1747)  | ~\4242(1580) ,
  \4548(1525)  = ~\7486(1173)  | ~\7479(890) ,
  \7264(1387)  = ~\7260(1040) ,
  \6474(1269)  = \2175(975) ,
  \6798(1863)  = ~\6796(1590)  | ~\6789(1253) ,
  \694(627)  = \693(524)  | \664(574) ,
  \5019(2691)  = ~\5017(1219)  | ~\5014(2482) ,
  \392(3022)  = ~\4863(2938)  | ~\4860(2358) ,
  \2876(389)  = \4514(292)  & \2857(293) ,
  \3481(3000)  = ~\3480(2765)  | ~\3479(2902) ,
  \6206(2747)  = \2742(2533) ,
  \7187(3571)  = ~\7185(3553)  | ~\7182(2262) ,
  \5158(3544)  = ~\5156(2439)  | ~\5149(3528) ,
  \1866(893)  = \731(855)  & \1178(261) ,
  \920(2100)  = \792(1841)  & (\805(1844)  & (\827(1874)  & (\853(1849)  & \895(1850) ))),
  \265(2835)  = \1002(2682)  | \908(1192) ,
  \1694(1542)  = ~\5464(1246)  | ~\5457(368) ,
  \295(3352)  = \[73] ,
  \1115(371)  = \1198(299)  & \1541(275) ,
  \1317(2748)  = \1299(2536)  & (\1253(2214)  & \1240(1950) ),
  \3605(2703)  = \3583(2472)  & (\3531(2480)  & \3540(2491) ),
  \5698(3215)  = ~\5696(2669)  | ~\5689(3164) ,
  \3511(1567)  = ~\6701(1281)  | ~\6698(938) ,
  \7344(2203)  = ~\7340(1931) ,
  \4896(1445)  = ~\4892(1090) ,
  \5959(2797)  = ~\5953(2618) ,
  \7388(1283)  = \2065(985) ,
  \7220(1633)  = ~\7216(1300) ,
  \887(922)  = ~\886(604)  | ~\885(832) ,
  \2553(3012)  = ~\2552(2794)  | ~\2551(2921) ,
  \1794(1510)  = ~\5752(1440)  | ~\5745(353) ,
  \5198(1461)  = ~\5194(1106) ,
  \940(2107)  = \853(1849)  & (\805(1844)  & (\827(1874)  & \895(1850) )),
  \4530(1185)  = ~\7470(915)  | ~\7463(913) ,
  \5715(3484)  = ~\5709(3467) ,
  \1330(3067)  = ~\5384(1953)  | ~\5377(2988) ,
  \382(3148)  = \[67] ,
  \7330(1067)  = \723(849) ,
  \7544(1345)  = \4508(1013) ,
  \5116(2840)  = ~\5112(2687) ,
  \2841(3662)  = ~\6260(2636)  | ~\6253(3645) ,
  \1903(1826)  = ~\1902(1537)  | ~\1901(1178) ,
  \5165(3600)  = ~\5159(3584) ,
  \4737(3220)  = \1971(3165)  | (\1969(2088)  | \1914(905) ),
  \1654(1538)  = ~\5448(1236)  | ~\5441(367) ,
  \6934(3003)  = ~\6932(2905)  | ~\6925(1115) ,
  \4844(2345)  = \2409(1989) ,
  \5767(473)  = ~\5761(357) ,
  \7283(1294)  = \2081(988) ,
  \6530(1053)  = \641(841) ,
  \3462(3197)  = \3399(1978)  & (\3381(1976)  & (\3417(1979)  & \2580(3145) )),
  \6001(340)  = \3739(233) ,
  \3223(1698)  = \3222(1366)  | \3221(557) ,
  \5828(2003)  = \1795(1804) ,
  \1804(1513)  = ~\5760(1441)  | ~\5753(354) ,
  \2598(1490)  = ~\5999(452)  | ~\5996(1260) ,
  \273(3402)  = \[86] ,
  \310(3393)  = \[77] ,
  \4633(2978)  = ~\4632(2731)  & ~\4631(2866) ,
  \3606(2966)  = ~\3605(2703)  & ~\3604(2853) ,
  \6402(951)  = \1395(814) ,
  \4586(2182)  = ~\4585(1908)  | ~\4584(1893) ,
  \5297(1062)  = \645(847) ,
  \6581(433)  = ~\6575(320) ,
  \2069(968)  = \2048(653)  | \2047(802) ,
  \7534(1348)  = \4502(1015) ,
  \6615(331)  = \4407(221) ,
  \5308(846)  = \601(422)  & \626(636) ,
  \7268(1046)  = \2316(837) ,
  \3050(1903)  = ~\6445(1670)  | ~\6442(1006) ,
  \3751(229)  = ~\3749(194) ,
  \3071(2195)  = ~\3070(1675)  | ~\3069(1934) ,
  \2618(1985)  = ~\2617(1787)  | ~\2616(1491) ,
  \325(3358)  = ~\4767(3297)  | ~\4764(2102) ,
  \3504(1851)  = ~\3503(1221)  | ~\3502(1573) ,
  \3308(1109)  = \3833(1016)  & \4434(211) ,
  \5464(1246)  = ~\5460(967) ,
  \2541(2918)  = ~\5943(2791)  | ~\5940(2310) ,
  \6233(3613)  = ~\6232(3578)  | ~\6231(3593) ,
  \4196(1605)  = ~\7227(1358)  | ~\7224(1270) ,
  \4538(1540)  = ~\7477(1174)  | ~\7474(908) ,
  \1968(3163)  = \1903(1826)  & (\1885(1825)  & (\1921(1832)  & \3279(3072) )),
  \6661(2768)  = ~\6655(2568) ,
  \4973(1548)  = ~\917(1190) ,
  \3441(2240)  = \3327(1111)  & \3295(1965) ,
  \4632(2731)  = \4610(2502)  & (\4558(2189)  & \4567(2501) ),
  \3030(2055)  = \2998(896)  & \2982(1816) ,
  \4502(1015)  = \4483(712)  | \4482(755) ,
  \4824(2593)  = ~\4820(2281) ,
  \397(3097)  = \[64] ,
  \6300(3453)  = ~\6298(2880)  | ~\6291(3385) ,
  \4517(3156)  = ~\4516(3024)  | ~\4515(3099) ,
  \6986(2769)  = ~\4017(2569) ,
  \1761(3562)  = ~\5580(2390)  | ~\5573(3538) ,
  \6901(332)  = \4402(223) ,
  \[37]  = ~\15(4) ,
  \6073(3150)  = ~\6067(3088) ,
  \5505(3480)  = ~\5504(3438)  | ~\5503(3465) ,
  \5274(864)  = \2905(426)  & \2930(613) ,
  \1742(2065)  = \1655(1827)  & (\1630(1824)  & \1695(1829) ),
  \1093(1853)  = ~\1092(1572)  | ~\1091(1224) ,
  \2551(2921)  = ~\5967(2796)  | ~\5964(2315) ,
  \7352(2464)  = ~\7348(2148) ,
  \2963(1741)  = ~\6381(1151)  | ~\6378(1066) ,
  \4653(410)  = \1524(301) ,
  \4089(2553)  = \4020(2264)  & \4004(2224) ,
  \2561(2925)  = ~\2560(2800)  | ~\2559(2624) ,
  \3574(2438)  = ~\3571(2096) ,
  \6310(3500)  = ~\6308(2647)  | ~\6301(3490) ,
  \2555(2627)  = ~\5975(1498)  | ~\5972(2331) ,
  \4144(706)  = \4107(585)  & \60(23) ,
  \4775(3303)  = ~\4769(3242) ,
  \5832(2381)  = ~\5828(2003) ,
  \[41]  = ~\401(310)  | ~\400(297) ,
  \[42]  = ~\2857(293) ,
  \5543(3212)  = ~\5542(3102)  | ~\5541(3159) ,
  \[43]  = ~\4514(292) ,
  \360(3379)  = ~\4815(3325)  | ~\4812(2269) ,
  \5014(2482)  = \946(2122)  | (\945(2128)  | (\944(2114)  | \845(980) )),
  \5481(3105)  = ~\5475(3038) ,
  \6503(1315)  = \4151(997) ,
  \[44]  = ~\4442(290) ,
  \6859(431)  = ~\6853(318) ,
  \2499(2782)  = ~\2495(2601) ,
  \[45]  = ~\1501(291) ,
  \1102(940)  = \2933(861)  & \1464(285) ,
  \4920(565)  = ~\4916(400) ,
  \2008(3214)  = \2007(3161)  | \1957(2411) ,
  \6253(3645)  = ~\6252(3614)  | ~\6251(3634) ,
  \1573(1810)  = ~\1572(1517)  | ~\1571(1156) ,
  \[48]  = ~\574(308)  | ~\1197(165) ,
  \6736(1629)  = ~\6732(1295) ,
  \5740(3694)  = \1787(3678)  | \1786(3686) ,
  \[49]  = ~\1205(305) ,
  \2999(1578)  = ~\6413(1175)  | ~\6410(950) ,
  \965(2958)  = ~\962(2839) ,
  \1841(883)  = \2241(257)  & \737(854) ,
  \1994(2945)  = ~\1993(2659)  | ~\1992(2820) ,
  \5903(457)  = ~\5897(344) ,
  \1122(2101)  = \1074(1846)  & (\1026(1842)  & (\1055(1875)  & (\1093(1853)  & \1038(1843) ))),
  \2515(2628)  = \2514(2523)  | (\2513(2362)  | (\2512(2354)  | (\2511(2348)  | \2417(1138) ))),
  \6450(1017)  = \3810(823) ,
  \3009(1828)  = ~\3008(1539)  | ~\3007(1575) ,
  \4429(213)  = ~\4427(202) ,
  \1319(2883)  = ~\1318(2535)  & ~\1317(2748) ,
  \5508(2001)  = \1546(1803) ,
  \929(2433)  = \928(2126)  | (\927(2112)  | (\926(2163)  | (\925(2103)  | \802(924) ))),
  \1263(1857)  = ~\1262(1234)  | ~\1261(1582) ,
  \7273(1258)  = \2073(971) ,
  \[50]  = ~\574(308)  | ~\1197(165) ,
  \745(853)  = \671(424)  & \706(640) ,
  \5362(1956)  = ~\5348(1749)  | ~\5347(1750) ,
  \[51]  = ~\575(309)  | ~\1184(294) ,
  \6975(3549)  = ~\6974(3512)  | ~\6973(3531) ,
  \[52]  = ~\1205(305) ,
  \657(404)  = \1512(300) ,
  \[53]  = ~\280(391) ,
  \6162(2604)  = ~\6158(2308) ,
  \[55]  = \572(427)  & \163(86) ,
  \7290(1600)  = ~\7286(1264) ,
  \[56]  = ~\372(2890)  | ~\371(2754) ,
  \2366(1130)  = \2105(972)  & \3745(231) ,
  \[57]  = \245(2897)  | (\244(3033)  | (\243(3032)  | (\242(2955)  | \241(2837) ))),
  \390(2934)  = ~\4856(2639)  | ~\4849(2807) ,
  \6281(3209)  = ~\6280(3096)  | ~\6279(3155) ,
  \[58]  = \257(2860)  | (\256(2991)  | (\255(2990)  | (\254(2888)  | \3259(2874) ))),
  \3431(2229)  = \3283(1964)  & (\3314(1967)  & (\3344(1970)  & \3295(1965) )),
  \3393(1121)  = \2192(991)  & \4407(221) ,
  \4903(671)  = ~\4897(548) ,
  \[59]  = \263(2858)  | (\262(2993)  | (\261(2992)  | (\260(2889)  | \3259(2874) ))),
  \5099(1218)  = \877(939) ,
  \1350(415)  = \1503(303) ,
  \4122(751)  = \4101(734)  & \4121(228) ,
  \3908(1118)  = \3816(1021)  & \4417(217) ,
  \5944(2606)  = ~\5940(2310) ,
  \7334(1422)  = ~\7330(1067) ,
  \3534(1882)  = ~\6735(1634)  | ~\6732(1295) ,
  \6040(1710)  = ~\6036(1383) ,
  \5253(1453)  = ~\5247(1098) ,
  \6931(1471)  = ~\6925(1115) ,
  \2000(2667)  = ~\5856(2398)  | ~\5849(884) ,
  \2353(1785)  = ~\5880(1596)  | ~\5873(338) ,
  \731(855)  = \671(424)  & \702(638) ,
  \7197(3642)  = \4086(3630)  | (\4085(3629)  | (\4084(3627)  | \4083(3628) )),
  \[60]  = \269(2896)  | (\268(3028)  | (\267(3027)  | (\266(2956)  | \265(2835) ))),
  \4053(2910)  = \4023(2582)  & \4032(2773) ,
  \4287(2457)  = \4267(2143)  & (\4230(2140)  & \4239(2141) ),
  \[61]  = ~\387(2931)  | ~\386(3020) ,
  \1947(2035)  = \1841(883)  & \1822(1811) ,
  \[62]  = ~\390(2934)  | ~\389(3021) ,
  \548(234)  = \3737(192) ,
  \5788(964)  = \1418(819) ,
  \3813(822)  = \3790(551)  | \3789(625) ,
  \6461(1676)  = ~\6455(1337) ,
  \[63]  = ~\393(2937)  | ~\392(3022) ,
  \6270(2986)  = ~\6268(2808)  | ~\6261(1944) ,
  \4598(2042)  = \4549(1815) ,
  \[64]  = ~\396(2941)  | ~\395(3023) ,
  \4999(3047)  = ~\4997(1555)  | ~\4990(2953) ,
  \[65]  = \375(3090)  | \374(3152) ,
  \4873(373)  = \1541(275) ,
  \6519(928)  = \3679(776) ,
  \[66]  = \378(3091)  | \377(3153) ,
  \5884(1255)  = \2099(970) ,
  \5518(2011)  = \1556(1807) ,
  \7041(1127)  = ~\2179(977)  & ~\4396(225) ,
  \3476(2903)  = ~\6661(2768)  | ~\6658(2233) ,
  \[67]  = \381(3092)  | \380(3086) ,
  \7324(1426)  = ~\7320(1071) ,
  \4388(2971)  = \4387(2850)  | \4364(2720) ,
  \2050(656)  = \2019(576)  & \127(64) ,
  \[68]  = \384(3016)  | \383(3089) ,
  \5873(338)  = \3745(231) ,
  \5512(2377)  = ~\5508(2001) ,
  \[69]  = ~\4443(3309) ,
  \5170(3696)  = \996(3683)  | \995(3691) ,
  \4166(995)  = \4141(690)  | \4140(745) ,
  \3109(1892)  = ~\6494(1632)  | ~\6487(1313) ,
  \7417(1349)  = \4502(1015) ,
  \1783(3615)  = \1771(3137)  & (\1726(2407)  & \1757(3594) ),
  \1973(3167)  = \1921(1832)  & \3279(3072) ,
  \4622(2673)  = \4601(2406)  & (\4540(1822)  & \4535(2093) ),
  \7094(2263)  = \3899(1971) ,
  \5745(353)  = \1192(251) ,
  \2434(1503)  = ~\5919(461)  | ~\5916(1390) ,
  \6191(3208)  = ~\6189(3187)  | ~\6186(2811) ,
  \5189(607)  = ~\5183(498) ,
  \399(3717)  = \[107] ,
  \5342(1079)  = \737(854) ,
  \7377(1347)  = \4505(1014) ,
  \2064(675)  = \2032(592)  & \100(51) ,
  \1399(820)  = \1376(546)  | \1375(643) ,
  \6165(3554)  = ~\6164(3517)  | ~\6163(3534) ,
  \7023(3493)  = ~\7022(3455)  | ~\7021(3475) ,
  \1172(3419)  = \1171(3307)  | \1170(3367) ,
  \5630(3482)  = ~\5628(2426)  | ~\5621(3468) ,
  \[70]  = ~\4524(3265) ,
  \627(535)  = \606(403)  & \164(87) ,
  \1677(909)  = \1399(820)  & \2213(268) ,
  \[71]  = ~\2868(3308) ,
  \708(641)  = \707(544)  | \685(588) ,
  \245(2897)  = \1146(2431)  & (\1974(2382)  & (\3466(2558)  & (\2532(2788)  & \4526(205) ))),
  \[72]  = \248(3306)  | \247(3310) ,
  \7549(1913)  = ~\7547(1680)  | ~\7544(1345) ,
  \2150(680)  = \2117(577)  & \94(49) ,
  \4475(695)  = \4444(582)  & \74(33) ,
  \[73]  = ~\294(3223)  | ~\293(3285) ,
  \5305(845)  = \601(422)  & \628(637) ,
  \5452(1077)  = \737(854) ,
  \[74]  = ~\323(3238)  | ~\322(3302) ,
  \5352(1088)  = \751(857) ,
  \[75]  = \251(3365)  | \250(3417) ,
  \[76]  = \275(3286)  | \274(3353) ,
  \6650(2228)  = \3283(1964) ,
  \5292(1056)  = \633(843) ,
  \4067(3144)  = \2851(3008)  | \2850(3083) ,
  \[77]  = ~\309(3275)  | ~\308(3346) ,
  \2398(1497)  = ~\5895(456)  | ~\5892(1250) ,
  \[78]  = ~\312(3279)  | ~\311(3349) ,
  \1328(3191)  = ~\1327(3071)  | ~\1326(3135) ,
  \369(3714)  = ~\4093(3710)  | ~\4092(3705) ,
  \[79]  = ~\315(3281)  | ~\314(3350) ,
  \3590(2717)  = ~\3587(2489) ,
  \1962(2086)  = \1869(1819)  & (\1929(910)  & (\1885(1825)  & \1903(1826) )),
  \986(3677)  = ~\985(3653)  | ~\984(3668) ,
  \5522(2389)  = ~\5518(2011) ,
  \432(428)  = \573(311) ,
  \6274(2812)  = ~\2801(2645) ,
  \6990(2904)  = ~\6986(2769) ,
  \2207(272)  = ~\2204(174) ,
  \6843(3118)  = ~\6837(3056) ,
  \3650(666)  = \3629(578)  & \113(58) ,
  \4233(1576)  = ~\7307(1228)  | ~\7304(948) ,
  \7539(1916)  = ~\7537(1684)  | ~\7534(1348) ,
  \5412(1076)  = \745(853) ,
  \7375(1682)  = ~\7369(1344) ,
  \534(220)  = \4410(199) ,
  \5502(2395)  = ~\5498(2023) ,
  \[80]  = ~\318(3283)  | ~\317(3351) ,
  \1726(2407)  = \1725(2081)  | (\1724(2069)  | (\1723(2058)  | (\1722(2049)  | \1606(892) ))),
  \6526(1418)  = ~\6522(1063) ,
  \6566(1414)  = ~\6562(1059) ,
  \[81]  = ~\326(3294)  | ~\325(3358) ,
  \1454(2894)  = \4089(2553)  & (\2852(2785)  & \4526(205) ),
  \[82]  = ~\329(3298)  | ~\328(3361) ,
  \7137(2780)  = ~\7135(1780)  | ~\7132(2589) ,
  \[83]  = ~\332(3304)  | ~\331(3364) ,
  \4815(3325)  = ~\4809(3253) ,
  \5584(2419)  = \1742(2065)  | (\1741(2083)  | (\1740(2071)  | \1647(899) )),
  \3653(506)  = \3622(407)  & \1471(283) ,
  \3080(1920)  = ~\6469(1642)  | ~\6466(1019) ,
  \5135(3409)  = ~\5129(3359) ,
  \[84]  = ~\335(3300)  | ~\334(3362) ,
  \6304(2370)  = \2701(1995) ,
  \[85]  = ~\417(3415) ,
  \448(284)  = \1469(169) ,
  \914(1200)  = \765(774)  & \887(922) ,
  \6501(1645)  = ~\6495(1311) ,
  \[86]  = \272(3287)  | \271(3354) ,
  \1003(3702)  = ~\5173(3469)  | ~\5170(3696) ,
  \7252(825)  = \2286(554)  | \2285(616) ,
  \308(3346)  = ~\4727(3278)  | ~\4724(2048) ,
  \[87]  = \297(3266)  | \296(3340) ,
  \7466(771)  = \4667(492)  | \4666(687) ,
  \7071(3378)  = ~\7070(3252)  | ~\7069(3323) ,
  \4804(2266)  = \3353(1972) ,
  \1364(519)  = \1336(405)  & \181(104) ,
  \5460(967)  = \1399(820) ,
  \[88]  = \300(3267)  | \299(3341) ,
  \6361(2702)  = ~\7352(2464)  | ~\7345(2154) ,
  \7011(3373)  = ~\7009(3312)  | ~\7006(2259) ,
  \[89]  = \303(3271)  | \302(3342) ,
  \5983(1789)  = ~\5977(1493) ,
  \6469(1642)  = ~\6463(1309) ,
  \938(2111)  = \805(1844)  & (\868(934)  & \827(1874) ),
  \5493(3345)  = ~\5491(3269)  | ~\5488(2039) ,
  \5202(1089)  = \2946(858) ,
  \4201(1695)  = ~\7255(1364)  | ~\7252(825) ,
  \4247(2477)  = \4198(2157) ,
  \3060(1919)  = ~\6453(1673)  | ~\6450(1017) ,
  \484(256)  = \2247(182) ,
  \2699(1505)  = ~\6039(463)  | ~\6036(1383) ,
  \1216(1757)  = ~\5254(1456)  | ~\5247(1098) ,
  \5271(863)  = \2905(426)  & \2932(614) ,
  \5857(1159)  = \1841(883) ,
  \7486(1173)  = ~\7482(898) ,
  \[90]  = \306(3270)  | \305(3343) ,
  \5365(2218)  = ~\5359(1957) ,
  \996(3683)  = \986(3677)  & \975(3157) ,
  \[91]  = ~\343(3258)  | ~\342(3330) ,
  \4047(2302)  = \3979(1126)  & \3957(1977) ,
  \1005(721)  = ~\5181(494)  | ~\5178(399) ,
  \2846(3623)  = \2828(208)  & (\2813(2930)  & \2824(3611) ),
  \4326(1655)  = ~\7400(1398)  | ~\7393(1319) ,
  \5031(3178)  = ~\5030(3051)  | ~\5029(3114) ,
  \2855(3703)  = ~\6335(3656)  | ~\6332(3697) ,
  \6085(3384)  = ~\6083(3332)  | ~\6080(2343) ,
  \6278(2940)  = ~\6274(2812) ,
  \1378(538)  = \1350(415)  & \160(83) ,
  \1942(2018)  = \1834(878)  & \1805(1806) ,
  \2431(1140)  = \2335(1044)  & \3719(239) ,
  \[96]  = ~\358(3320)  | ~\357(3376) ,
  \[97]  = ~\361(3324)  | ~\360(3379) ,
  \[98]  = ~\364(3326)  | ~\363(3380) ,
  \5604(2414)  = \1736(2053)  | (\1735(2080)  | (\1734(2068)  | (\1733(2057)  | \1624(894) ))),
  \[99]  = ~\367(3328)  | ~\366(3381) ,
  \6837(3056)  = ~\3603(2969)  | ~\3606(2966) ,
  \5312(1061)  = ~\5308(846) ,
  \5587(1183)  = ~\5581(911) ,
  \2292(570)  = \2259(413)  & \26(7) ,
  \3853(1108)  = \3838(1004)  & \4439(209) ,
  \2391(1134)  = \3731(235)  & \2091(969) ,
  \3234(2137)  = \3186(1845)  & (\3209(942)  & (\3176(1840)  & (\3195(1876)  & \3203(1847) ))),
  \6590(1707)  = ~\6586(1378) ,
  \3295(1965)  = ~\3294(1764)  | ~\3293(1465) ,
  \7415(1659)  = ~\7409(1321) ,
  \3365(1973)  = ~\3364(1774)  | ~\3363(1477) ,
  \3480(2765)  = ~\6670(2563)  | ~\6663(2567) ,
  \5708(3399)  = ~\5706(2428)  | ~\5699(3347) ,
  \255(2990)  = \3249(2223)  & (\3035(2374)  & \3164(2980) ),
  \4628(2865)  = \4609(2729)  & (\4563(2184)  & \4558(2189) ),
  \2643(1990)  = ~\2642(1794)  | ~\2641(1500) ,
  \5409(356)  = \2249(255) ,
  \7107(3607)  = ~\7101(3589) ,
  \1318(2535)  = \1296(2212)  & (\1244(2211)  & \1253(2214) ),
  \928(2126)  = \805(1844)  & (\877(939)  & (\792(1841)  & (\827(1874)  & \853(1849) ))),
  \3783(622)  = \3762(586)  & \192(115) ,
  \5809(369)  = \2213(268) ,
  \7114(2272)  = \3911(1974) ,
  \4014(2241)  = \3885(1112)  & \3856(1966) ,
  \2780(2629)  = \2779(2527)  | (\2778(2366)  | (\2777(2357)  | (\2776(2349)  | \2652(1139) ))),
  \3470(2758)  = ~\6646(2556)  | ~\6639(2560) ,
  \1132(2164)  = \1068(981)  & \1038(1843) ,
  \2105(972)  = \2062(657)  | \2061(788) ,
  \358(3320)  = ~\4808(2583)  | ~\4801(3250) ,
  \4273(2968)  = ~\4272(2710)  & ~\4271(2857) ,
  \993(3406)  = \975(3157)  & (\962(2839)  & \971(3356) ),
  \4039(2275)  = \3949(1122)  & \3911(1974) ,
  \4756(2139)  = \1093(1853) ,
  \2756(2339)  = \2600(1984)  & (\2635(1135)  & (\2589(1981)  & \2618(1985) )),
  \5728(3540)  = ~\5726(2408)  | ~\5719(3526) ,
  \1054(1615)  = ~\5214(1449)  | ~\5207(549) ,
  \1998(3036)  = ~\1997(2944) ,
  \7584(1906)  = ~\7582(1646)  | ~\7575(1338) ,
  \948(2130)  = \877(939)  & (\827(1874)  & \853(1849) ),
  \7124(2270)  = \3911(1974) ,
  \6647(2559)  = ~\3442(2251)  & (~\3441(2240)  & ~\3308(1109) ),
  \4667(492)  = \4640(409)  & \2210(270) ,
  \7104(2279)  = \3932(1975) ,
  \924(2441)  = ~\920(2100) ,
  \4792(2449)  = ~\4788(2118) ,
  \3642(579)  = ~\3635(408) ,
  \2956(1802)  = ~\2955(1508)  | ~\2954(1740) ,
  \3615(3168)  = ~\3614(3044)  | ~\3613(3108) ,
  \3239(3025)  = \3035(2374)  & \3164(2980) ,
  \5847(2663)  = ~\5841(2392) ,
  \7594(1904)  = ~\7592(1674)  | ~\7585(1334) ,
  \377(3153)  = \2571(3018)  & \2554(3085) ,
  \6324(2359)  = \2676(1994) ,
  \3013(906)  = \1387(812)  & \4689(769) ,
  \5346(1434)  = ~\5342(1079) ,
  \401(310)  = ~\5(1) ,
  \3791(795)  = \3775(740)  & \223(146) ,
  \4280(2872)  = \4262(2715)  & (\4216(2206)  & \4203(1923) ),
  \4957(3112)  = ~\4955(3046)  | ~\4952(1204) ,
  \4735(3280)  = ~\4729(3218) ,
  \1518(278)  = \1492(172)  & \4528(206) ,
  \4336(2185)  = ~\4335(1653)  | ~\4334(1939) ,
  \2776(2349)  = \2670(1141)  & \2643(1990) ,
  \1816(875)  = \751(857)  & \1186(254) ,
  \2964(1512)  = ~\6382(1421)  | ~\6375(874) ,
  \7316(1231)  = ~\7312(952) ,
  \4863(2938)  = ~\4857(2810) ,
  \6796(1590)  = ~\6792(1252) ,
  \6203(3437)  = ~\6202(3336)  | ~\6201(3386) ,
  \4088(3688)  = \4078(3680)  & \4067(3144) ,
  \1707(2029)  = \1556(1807)  & (\1590(882)  & (\1546(1803)  & \1573(1810) )),
  \6517(598)  = ~\6511(429) ,
  \6399(897)  = \4695(767) ,
  \699(527)  = \657(404)  & \173(96) ,
  \3810(823)  = \3788(552)  | \3787(624) ,
  \5775(474)  = ~\5769(358) ,
  \7084(2290)  = \3957(1977) ,
  \4480(756)  = \4464(733)  & \3725(237) ,
  \3587(2489)  = \3568(2172) ,
  \5358(1752)  = ~\5356(1443)  | ~\5349(1083) ,
  \1036(1210)  = ~\5205(502)  | ~\5202(1089) ,
  \2766(2340)  = \2600(1984)  & (\2635(1135)  & \2618(1985) ),
  \7609(2507)  = ~\7603(2196) ,
  \5677(2676)  = ~\5675(1541)  | ~\5672(2418) ,
  \4078(3680)  = ~\4077(3659)  | ~\4076(3670) ,
  \3456(2273)  = \3393(1121)  & \3365(1973) ,
  \4412(219)  = ~\4410(199) ,
  \4004(2224)  = \3845(1963)  & (\3856(1966)  & (\3874(1968)  & \3989(1969) )),
  \7142(2778)  = ~\4048(2594) ,
  \4163(994)  = \4138(689)  | \4137(746) ,
  \2977(879)  = \719(850)  & \4704(764) ,
  \4288(2846)  = ~\4287(2457)  & ~\4286(2693) ,
  \6802(1261)  = \2105(972) ,
  \1802(871)  = \757(856)  & \1192(251) ,
  \2351(1128)  = \2111(987)  & \3751(229) ,
  \6806(1598)  = ~\6802(1261) ,
  \1786(3686)  = \1771(3137)  & \1781(3684) ,
  \3446(2265)  = \3399(1978)  & (\3353(1972)  & (\3381(1976)  & (\3417(1979)  & \3365(1973) ))),
  \6446(1332)  = ~\6442(1006) ,
  \6429(1165)  = ~\6423(888) ,
  \6410(950)  = \1391(813) ,
  \4362(2468)  = \4312(1256)  & (\4291(2173)  & \4300(2153) ),
  \5416(1431)  = ~\5412(1076) ,
  \3682(839)  = \3635(408)  | \3665(600) ,
  \1501(291)  = \199(122)  & (\188(111)  & (\172(95)  & \162(85) )),
  \5277(1102)  = ~\5271(863) ,
  \6623(333)  = \4402(223) ,
  \2922(609)  = \2921(512)  | \2899(590) ,
  \5553(3391)  = ~\5552(3272)  | ~\5551(3344) ,
  \6792(1252)  = \2091(969) ,
  \6039(463)  = ~\6033(350) ,
  \2506(2332)  = \2372(1986)  & \2400(1988) ,
  \5050(3414)  = ~\5048(2454)  | ~\5041(3360) ,
  \3868(1110)  = \3833(1016)  & \4434(211) ,
  \5456(1432)  = ~\5452(1077) ,
  \6776(1384)  = \2323(1038) ,
  \5356(1443)  = ~\5352(1088) ,
  \5060(3486)  = ~\5058(2451)  | ~\5051(3471) ,
  \6422(1226)  = ~\6418(947) ,
  \6780(1711)  = ~\6776(1384) ,
  \6123(2926)  = ~\6121(1790)  | ~\6118(2798) ,
  \6724(979)  = \2154(664)  | \2153(791) ,
  \6389(1154)  = ~\6383(880) ,
  \1554(1153)  = ~\5407(470)  | ~\5404(1087) ,
  \4275(2707)  = \4251(2476)  & (\4184(2479)  & \4193(2493) ),
  \5928(1709)  = ~\5924(1382) ,
  \5296(1411)  = ~\5292(1056) ,
  \4009(2256)  = \3856(1966)  & (\3891(1114)  & (\3845(1963)  & \3874(1968) )),
  \1176(1838)  = ~\1112(1553)  | ~\1121(1552) ,
  \4349(1400)  = \3695(1050)  & \3686(838) ,
  \3487(2574)  = ~\6685(1768)  | ~\6682(2244) ,
  \6586(1378)  = \3828(1035) ,
  \7129(1483)  = \3979(1126) ,
  \6320(3556)  = ~\6318(2632)  | ~\6311(3537) ,
  \4752(2425)  = ~\4748(2075) ,
  \7276(1247)  = \2069(968) ,
  \1746(2424)  = \1745(2084)  | \1669(904) ,
  \7155(3255)  = ~\7149(3198) ,
  \2674(1504)  = ~\6031(462)  | ~\6028(1389) ,
  \6574(1667)  = ~\6570(1329) ,
  \5206(1444)  = ~\5202(1089) ,
  \3059(1330)  = \3813(822)  & \4175(1007) ,
  \3436(2250)  = \3295(1965)  & (\3335(1113)  & (\3283(1964)  & \3314(1967) )),
  \4389(1405)  = \1535(302)  & \2320(1025) ,
  \404(390)  = \[42] ,
  \6243(3664)  = ~\6242(3635)  | ~\6241(3646) ,
  \1974(2382)  = \1950(2047)  & \1935(2004) ,
  \248(3306)  = \3223(1698)  & \3245(3230) ,
  \3461(2297)  = \3425(1125)  & (\3381(1976)  & \3399(1978) ),
  \6494(1632)  = ~\6490(1299) ,
  \4825(3257)  = \3465(3201)  | \3425(1125) ,
  \5686(2830)  = ~\5682(2674) ,
  \6067(3088)  = ~\6066(3015)  | ~\6065(2927) ,
  \5849(884)  = ~\2241(257)  & ~\737(854) ,
  \4083(3628)  = \4072(3202)  & (\4032(2773)  & \4064(3605) ),
  \4044(2280)  = \3957(1977)  & (\3932(1975)  & \3997(1980) ),
  \2580(3145)  = \2579(3011)  | \2578(3082) ,
  \2886(425)  = \1207(307) ,
  \6662(2564)  = ~\6658(2233) ,
  \6679(1469)  = \3335(1113) ,
  \5972(2331)  = \2372(1986) ,
  \3610(2873)  = \3594(2719)  & (\3563(2517)  & \3550(2199) ),
  \1722(2049)  = \1624(894)  & \1598(1817) ,
  \943(2127)  = \805(1844)  & (\877(939)  & (\827(1874)  & \853(1849) )),
  \3437(2551)  = \3436(2250)  | (\3435(2238)  | (\3434(2230)  | \3292(1107) )),
  \4325(1941)  = ~\7399(1656)  | ~\7396(1045) ,
  \4672(685)  = \4647(580)  & \84(43) ,
  \1712(2014)  = \1584(877)  & \1556(1807) ,
  \2302(727)  = \2272(594)  & \26(7) ,
  \5513(3524)  = ~\5511(3503)  | ~\5508(2001) ,
  \7064(2585)  = \4038(2271)  | (\4037(2298)  | (\4036(2286)  | (\4035(2276)  | \3926(1120) ))),
  \6867(434)  = ~\6861(321) ,
  \4380(2721)  = ~\89(48)  | ~\4369(2486) ,
  \4900(1093)  = \2942(859) ,
  \1292(2213)  = \1258(1951) ,
  \6963(3474)  = ~\6961(3457)  | ~\6958(2248) ,
  \5689(3164)  = ~\5688(3040)  | ~\5687(3106) ,
  \685(588)  = ~\678(414) ,
  \1730(2668)  = ~\1726(2407) ,
  \4562(1895)  = ~\7522(1660)  | ~\7515(1317) ,
  \4956(1556)  = ~\4952(1204) ,
  \556(242)  = \3711(188) ,
  \7463(913)  = \4686(770) ,
  \1026(1842)  = ~\1025(1560)  | ~\1024(1209) ,
  \6076(3147)  = ~\6074(2793)  | ~\6067(3088) ,
  \6948(2260)  = \3989(1969) ,
  \2077(973)  = \2052(658)  | \2051(804) ,
  \5620(3400)  = ~\5618(2429)  | ~\5611(3348) ,
  \7474(908)  = \4689(769) ,
  \5439(484)  = ~\5433(364) ,
  \542(246)  = \3701(186) ,
  \3451(2283)  = \3365(1973)  & (\3410(1123)  & (\3353(1972)  & \3381(1976) )),
  \5573(3538)  = ~\5572(3501)  | ~\5571(3523) ,
  \1624(894)  = \1418(819)  & \2232(262) ,
  \1919(1188)  = ~\5815(491)  | ~\5812(966) ,
  \1035(925)  = \2950(865)  & \1488(279) ,
  \1091(1224)  = ~\5229(510)  | ~\5226(1100) ;
endmodule

