// IWLS benchmark module "C5315.iscas" printed on Wed May 29 16:29:45 2002
module C5315 (\1(0) , \4(1) , \11(2) , \14(3) , \17(4) , \20(5) , \23(6) , \24(7) , \25(8) , \26(9) , \27(10) , \31(11) , \34(12) , \37(13) , \40(14) , \43(15) , \46(16) , \49(17) , \52(18) , \53(19) , \54(20) , \61(21) , \64(22) , \67(23) , \70(24) , \73(25) , \76(26) , \79(27) , \80(28) , \81(29) , \82(30) , \83(31) , \86(32) , \87(33) , \88(34) , \91(35) , \94(36) , \97(37) , \100(38) , \103(39) , \106(40) , \109(41) , \112(42) , \113(43) , \114(44) , \115(45) , \116(46) , \117(47) , \118(48) , \119(49) , \120(50) , \121(51) , \122(52) , \123(53) , \126(54) , \127(55) , \128(56) , \129(57) , \130(58) , \131(59) , \132(60) , \135(61) , \136(62) , \137(63) , \140(64) , \141(65) , \145(66) , \146(67) , \149(68) , \152(69) , \155(70) , \158(71) , \161(72) , \164(73) , \167(74) , \170(75) , \173(76) , \176(77) , \179(78) , \182(79) , \185(80) , \188(81) , \191(82) , \194(83) , \197(84) , \200(85) , \203(86) , \206(87) , \209(88) , \210(89) , \217(90) , \218(91) , \225(92) , \226(93) , \233(94) , \234(95) , \241(96) , \242(97) , \245(98) , \248(99) , \251(100) , \254(101) , \257(102) , \264(103) , \265(104) , \272(105) , \273(106) , \280(107) , \281(108) , \288(109) , \289(110) , \292(111) , \293(112) , \299(113) , \302(114) , \307(115) , \308(116) , \315(117) , \316(118) , \323(119) , \324(120) , \331(121) , \332(122) , \335(123) , \338(124) , \341(125) , \348(126) , \351(127) , \358(128) , \361(129) , \366(130) , \369(131) , \372(132) , \373(133) , \374(134) , \386(135) , \389(136) , \400(137) , \411(138) , \422(139) , \435(140) , \446(141) , \457(142) , \468(143) , \479(144) , \490(145) , \503(146) , \514(147) , \523(148) , \534(149) , \545(150) , \549(151) , \552(152) , \556(153) , \559(154) , \562(155) , \1497(156) , \1689(157) , \1690(158) , \1691(159) , \1694(160) , \2174(161) , \2358(162) , \2824(163) , \3173(164) , \3546(165) , \3548(166) , \3550(167) , \3552(168) , \3717(169) , \3724(170) , \4087(171) , \4088(172) , \4089(173) , \4090(174) , \4091(175) , \4092(176) , \4115(177) , \144(354) , \298(299) , \973(202) , \594(224) , \599(269) , \600(259) , \601(220) , \602(222) , \603(225) , \604(223) , \611(275) , \612(263) , \810(356) , \848(330) , \849(219) , \850(217) , \851(218) , \634(665) , \815(627) , \845(845) , \847(465) , \926(624) , \923(619) , \921(664) , \892(408) , \887(528) , \606(407) , \656(621) , \809(655) , \993(850) , \978(851) , \949(852) , \939(853) , \889(734) , \593(733) , \636(1280) , \704(1281) , \717(1282) , \820(1283) , \639(1275) , \673(1276) , \707(1277) , \715(1278) , \598(1623) , \610(1519) , \588(1696) , \615(1750) , \626(1752) , \632(1692) , \1002(1920) , \1004(1977) , \591(1894) , \618(1925) , \621(1893) , \629(1926) , \822(1933) , \838(2064) , \861(2070) , \623(2152) , \722(2131) , \832(2133) , \834(2123) , \836(2128) , \859(2132) , \871(2127) , \873(2124) , \875(2125) , \877(2126) , \998(2163) , \1000(2168) , \575(2240) , \585(2236) , \661(2178) , \693(2179) , \747(2187) , \752(2189) , \757(2190) , \762(2184) , \787(2186) , \792(2188) , \797(2191) , \802(2183) , \642(2222) , \664(2223) , \667(2224) , \670(2225) , \676(2229) , \696(2226) , \699(2227) , \702(2228) , \818(2273) , \813(2260) , \824(2274) , \826(2275) , \828(2233) , \830(2182) , \854(2268) , \863(2276) , \865(2277) , \867(2237) , \869(2181) , \712(2297) , \727(2298) , \732(2300) , \737(2279) , \742(2238) , \772(2299) , \777(2278) , \782(2239) , \645(2271) , \648(2295) , \651(2314) , \654(2315) , \679(2272) , \682(2296) , \685(2316) , \688(2317) , \843(2455) , \882(2456) , \767(2479) , \807(2480) , \658(2483) , \690(2484) );
input
  \131(59) ,
  \126(54) ,
  \4092(176) ,
  \386(135) ,
  \372(132) ,
  \64(22) ,
  \366(130) ,
  \446(141) ,
  \292(111) ,
  \226(93) ,
  \145(66) ,
  \3552(168) ,
  \210(89) ,
  \43(15) ,
  \185(80) ,
  \3546(165) ,
  \119(49) ,
  \332(122) ,
  \422(139) ,
  \245(98) ,
  \103(39) ,
  \83(31) ,
  \164(73) ,
  \25(8) ,
  \316(118) ,
  \302(114) ,
  \562(155) ,
  \556(153) ,
  \552(152) ,
  \97(37) ,
  \203(86) ,
  \122(52) ,
  \4(1) ,
  \117(47) ,
  \81(29) ,
  \76(26) ,
  \273(106) ,
  \257(102) ,
  \17(4) ,
  \1497(156) ,
  \4087(171) ,
  \141(65) ,
  \197(84) ,
  \217(90) ,
  \136(62) ,
  \120(50) ,
  \115(45) ,
  \34(12) ,
  \176(77) ,
  \373(133) ,
  \457(142) ,
  \3173(164) ,
  \241(96) ,
  \293(112) ,
  \155(70) ,
  \523(148) ,
  \53(19) ,
  \503(146) ,
  \1(0) ,
  \3717(169) ,
  \129(57) ,
  \113(43) ,
  \88(34) ,
  \323(119) ,
  \27(10) ,
  \14(3) ,
  \307(115) ,
  \234(95) ,
  \67(23) ,
  \26(9) ,
  \46(16) ,
  \188(81) ,
  \132(60) ,
  \288(109) ,
  \127(55) ,
  \280(107) ,
  \91(35) ,
  \264(103) ,
  \248(99) ,
  \86(32) ,
  \1690(158) ,
  \254(101) ,
  \106(40) ,
  \167(74) ,
  \70(24) ,
  \4090(174) ,
  \490(145) ,
  \1694(160) ,
  \2174(161) ,
  \4088(172) ,
  \2358(162) ,
  \146(67) ,
  \468(143) ,
  \191(82) ,
  \130(58) ,
  \374(134) ,
  \206(87) ,
  \3724(170) ,
  \11(2) ,
  \170(75) ,
  \2824(163) ,
  \534(149) ,
  \79(27) ,
  \3550(167) ,
  \23(6) ,
  \3548(166) ,
  \358(128) ,
  \514(147) ,
  \338(124) ,
  \348(126) ,
  \225(92) ,
  \324(120) ,
  \400(137) ,
  \123(53) ,
  \118(48) ,
  \37(13) ,
  \179(78) ,
  \82(30) ,
  \308(116) ,
  \158(71) ,
  \61(21) ,
  \281(108) ,
  \218(91) ,
  \265(104) ,
  \137(63) ,
  \182(79) ,
  \40(14) ,
  \1691(159) ,
  \1689(157) ,
  \121(51) ,
  \251(100) ,
  \20(5) ,
  \116(46) ,
  \80(28) ,
  \4091(175) ,
  \242(97) ,
  \4089(173) ,
  \100(38) ,
  \479(144) ,
  \161(72) ,
  \389(136) ,
  \299(113) ,
  \54(20) ,
  \140(64) ,
  \369(131) ,
  \49(17) ,
  \135(61) ,
  \289(110) ,
  \435(140) ,
  \94(36) ,
  \200(85) ,
  \114(44) ,
  \361(129) ,
  \109(41) ,
  \341(125) ,
  \4115(177) ,
  \351(127) ,
  \73(25) ,
  \335(123) ,
  \24(7) ,
  \331(121) ,
  \411(138) ,
  \149(68) ,
  \52(18) ,
  \194(83) ,
  \315(117) ,
  \209(88) ,
  \128(56) ,
  \112(42) ,
  \31(11) ,
  \559(154) ,
  \87(33) ,
  \173(76) ,
  \549(151) ,
  \545(150) ,
  \233(94) ,
  \272(105) ,
  \152(69) ;
output
  \861(2070) ,
  \615(1750) ,
  \298(299) ,
  \807(2480) ,
  \767(2479) ,
  \600(259) ,
  \658(2483) ,
  \859(2132) ,
  \877(2126) ,
  \634(665) ,
  \843(2455) ,
  \836(2128) ,
  \722(2131) ,
  \882(2456) ,
  \707(1277) ,
  \875(2125) ,
  \834(2123) ,
  \832(2133) ,
  \717(1282) ,
  \690(2484) ,
  \639(1275) ,
  \873(2124) ,
  \851(218) ,
  \599(269) ,
  \849(219) ,
  \715(1278) ,
  \848(330) ,
  \871(2127) ,
  \636(1280) ,
  \704(1281) ,
  \1002(1920) ,
  \820(1283) ,
  \601(220) ,
  \673(1276) ,
  \1004(1977) ,
  \611(275) ,
  \144(354) ,
  \847(465) ,
  \815(627) ,
  \588(1696) ,
  \810(356) ,
  \993(850) ,
  \921(664) ,
  \632(1692) ,
  \809(655) ,
  \887(528) ,
  \602(222) ,
  \598(1623) ,
  \889(734) ,
  \656(621) ,
  \612(263) ,
  \732(2300) ,
  \688(2317) ,
  \973(202) ,
  \926(624) ,
  \685(2316) ,
  \654(2315) ,
  \777(2278) ,
  \818(2273) ,
  \737(2279) ,
  \651(2314) ,
  \826(2275) ,
  \865(2277) ,
  \1000(2168) ,
  \679(2272) ,
  \824(2274) ,
  \978(851) ,
  \863(2276) ,
  \854(2268) ,
  \648(2295) ,
  \645(2271) ,
  \813(2260) ,
  \727(2298) ,
  \603(225) ,
  \682(2296) ,
  \772(2299) ,
  \712(2297) ,
  \699(2227) ,
  \828(2233) ,
  \845(845) ,
  \892(408) ,
  \676(2229) ,
  \696(2226) ,
  \667(2224) ,
  \867(2237) ,
  \923(619) ,
  \591(1894) ,
  \629(1926) ,
  \618(1925) ,
  \664(2223) ,
  \621(1893) ,
  \610(1519) ,
  \782(2239) ,
  \869(2181) ,
  \642(2222) ,
  \585(2236) ,
  \742(2238) ,
  \594(224) ,
  \575(2240) ,
  \787(2186) ,
  \670(2225) ,
  \747(2187) ,
  \606(407) ,
  \702(2228) ,
  \850(217) ,
  \949(852) ,
  \822(1933) ,
  \802(2183) ,
  \623(2152) ,
  \939(853) ,
  \838(2064) ,
  \752(2189) ,
  \792(2188) ,
  \830(2182) ,
  \998(2163) ,
  \762(2184) ,
  \604(223) ,
  \693(2179) ,
  \757(2190) ,
  \797(2191) ,
  \661(2178) ,
  \593(733) ,
  \626(1752) ;
wire
  \2646(548) ,
  \4938(1989) ,
  \1837(1038) ,
  \4961(1474) ,
  \3998(367) ,
  \2752(544) ,
  \2959(489) ,
  \3249(486) ,
  \2675(896) ,
  \3570(382) ,
  \3449(1624) ,
  \4981(1488) ,
  \4582(2265) ,
  \1207(1811) ,
  \3467(1396) ,
  \4027(2235) ,
  \5251(1922) ,
  \576(1776) ,
  \2335(1869) ,
  \2581(894) ,
  \774(2195) ,
  \2442(195) ,
  \2879(960) ,
  \734(2196) ,
  \5362(586) ,
  \3119(470) ,
  \5121(1048) ,
  \2922(518) ,
  \3132(513) ,
  \4786(421) ,
  \3540(2164) ,
  \1849(1148) ,
  \4068(1980) ,
  \5034(2203) ,
  \3125(485) ,
  \4956(2267) ,
  \3476(1399) ,
  \2811(1298) ,
  \1224(1777) ,
  \773(2194) ,
  \5340(318) ,
  \2906(525) ,
  \1237(1818) ,
  \5331(1387) ,
  \733(2197) ,
  \2875(956) ,
  \3965(2153) ,
  \5366(598) ,
  \633(365) ,
  \2809(1234) ,
  \4507(1571) ,
  \2871(957) ,
  \4503(2288) ,
  \4086(2231) ,
  \2361(325) ,
  \5285(1424) ,
  \4481(1904) ,
  \2454(385) ,
  \3475(1398) ,
  \3358(350) ,
  \5096(491) ,
  \4207(1545) ,
  \3497(1626) ,
  \1889(1850) ,
  \1660(799) ,
  \4199(1544) ,
  \4432(2210) ,
  \4991(1414) ,
  \1948(1993) ,
  \3466(1395) ,
  \3891(1305) ,
  \1729(1146) ,
  \1287(1160) ,
  \3305(476) ,
  \5108(300) ,
  \4840(2262) ,
  \2337(2033) ,
  \5196(1092) ,
  \4660(1050) ,
  \4284(240) ,
  \5348(335) ,
  \2572(436) ,
  \1151(1195) ,
  \3542(2023) ,
  \5165(1097) ,
  \5151(1375) ,
  \3215(487) ,
  \2566(440) ,
  \4492(2215) ,
  \1388(1181) ,
  \3219(488) ,
  \1033(1161) ,
  \4899(2207) ,
  \3136(529) ,
  \4591(2287) ,
  \4527(1582) ,
  \4085(2232) ,
  \779(2139) ,
  \1225(1819) ,
  \1776(1131) ,
  \5399(946) ,
  \3837(1653) ,
  \3555(332) ,
  \3289(871) ,
  \5150(1373) ,
  \1204(1813) ,
  \3485(1388) ,
  \2081(970) ,
  \1022(1164) ,
  \1276(1165) ,
  \3458(1607) ,
  \1766(1135) ,
  \1846(1147) ,
  \689(2482) ,
  \1222(1820) ,
  \1757(1141) ,
  \4183(257) ,
  \4935(1917) ,
  \2430(383) ,
  \5161(1385) ,
  \4215(1541) ,
  \4615(1581) ,
  \778(2138) ,
  \3472(1641) ,
  \659(2121) ,
  \3887(1654) ,
  \4822(1995) ,
  \3972(184) ,
  \3285(876) ,
  \4780(230) ,
  \2991(857) ,
  \4595(1574) ,
  \4957(2216) ,
  \1242(1829) ,
  \3962(2154) ,
  \5090(274) ,
  \4500(2286) ,
  \1252(1824) ,
  \4569(1905) ,
  \4537(1592) ,
  \4788(229) ,
  \5286(1431) ,
  \4231(1521) ,
  \5160(1380) ,
  \4937(1938) ,
  \4547(1591) ,
  \1935(1994) ,
  \739(2140) ,
  \1885(1858) ,
  \2344(795) ,
  \764(2471) ,
  \2985(858) ,
  \4167(251) ,
  \879(2452) ,
  \657(2481) ,
  \4148(1098) ,
  \2639(316) ,
  \2631(323) ,
  \1775(983) ,
  \4764(237) ,
  \3481(1643) ,
  \1789(865) ,
  \5429(1642) ,
  \2635(317) ,
  \1051(1156) ,
  \3231(981) ,
  \804(2470) ,
  \1919(1874) ,
  \5015(1915) ,
  \4306(447) ,
  \4879(1944) ,
  \1954(1997) ,
  \2561(336) ,
  \4223(1540) ,
  \738(2141) ,
  \5284(1437) ,
  \3387(699) ,
  \2059(975) ,
  \4391(1547) ,
  \4880(1996) ,
  \3232(418) ,
  \763(2472) ,
  \2541(346) ,
  \4104(1462) ,
  \1852(1149) ,
  \1886(1975) ,
  \1909(1876) ,
  \4401(1537) ,
  \5098(290) ,
  \1749(988) ,
  \4558(1359) ,
  \4859(1384) ,
  \3651(2193) ,
  \5328(1077) ,
  \1664(1870) ,
  \4319(1091) ,
  \2549(341) ,
  \2338(796) ,
  \2597(667) ,
  \2600(388) ,
  \2066(1299) ,
  \1943(1992) ,
  \1305(1157) ,
  \4869(1378) ,
  \568(2008) ,
  \4156(1094) ,
  \2193(2403) ,
  \2709(1183) ,
  \2545(345) ,
  \4585(1594) ,
  \2776(939) ,
  \3346(943) ,
  \5209(925) ,
  \1462(1817) ,
  \3342(942) ,
  \1882(1857) ,
  \3926(1667) ,
  \2575(881) ,
  \4010(1981) ,
  \2772(937) ,
  \844(657) ,
  \1115(1185) ,
  \2405(329) ,
  \719(2030) ,
  \2341(2032) ,
  \1363(1184) ,
  \567(2009) ,
  \3895(738) ,
  \5025(1987) ,
  \1489(2393) ,
  \4743(1415) ,
  \3282(928) ,
  \3845(963) ,
  \4707(1377) ,
  \3790(2025) ,
  \3090(753) ,
  \4114(359) ,
  \3444(1368) ,
  \5069(1487) ,
  \2192(2404) ,
  \5409(1998) ,
  \3241(968) ,
  \582(2106) ,
  \4381(1529) ,
  \1528(215) ,
  \2139(1792) ,
  \4324(249) ,
  \569(2012) ,
  \3080(751) ,
  \1342(1189) ,
  \803(2469) ,
  \1893(1972) ,
  \2569(884) ,
  \4164(1090) ,
  \2766(593) ,
  \1215(1948) ,
  \4699(1382) ,
  \3255(854) ,
  \4652(920) ,
  \3453(1361) ,
  \5325(1070) ,
  \5321(1421) ,
  \2191(2402) ,
  \2171(2400) ,
  \3443(1369) ,
  \2328(2473) ,
  \1883(1974) ,
  \4900(2281) ,
  \758(2031) ,
  \5134(1054) ,
  \5320(1418) ,
  \3461(1370) ,
  \4300(244) ,
  \4357(1957) ,
  \1420(1175) ,
  \5145(1058) ,
  \5199(1089) ,
  \4802(411) ,
  \3616(182) ,
  \5049(1475) ,
  \1133(1180) ,
  \3961(2116) ,
  \1793(1128) ,
  \3906(938) ,
  \5155(1069) ,
  \2019(978) ,
  \5016(1968) ,
  \1811(1125) ,
  \1924(1872) ,
  \4715(1376) ,
  \2001(987) ,
  \1219(1900) ,
  \1914(1875) ,
  \2619(1171) ,
  \5189(1082) ,
  \4072(821) ,
  \3538(2117) ,
  \1875(1279) ,
  \2190(2401) ,
  \1214(1801) ,
  \2615(1155) ,
  \671(966) ,
  \5213(1061) ,
  \572(2113) ,
  \3411(878) ,
  \3251(861) ,
  \2655(306) ,
  \1598(610) ,
  \4841(2208) ,
  \3301(870) ,
  \2651(307) ,
  \3076(907) ,
  \5299(1122) ,
  \691(2122) ,
  \1487(2384) ,
  \5389(1499) ,
  \4436(2283) ,
  \2692(902) ,
  \2536(591) ,
  \2148(1615) ,
  \3192(829) ,
  \3062(901) ,
  \4799(1045) ,
  \3421(888) ,
  \2705(1186) ,
  \4378(2284) ,
  \1890(1973) ,
  \1212(1949) ,
  \4804(234) ,
  \1488(2372) ,
  \2702(910) ,
  \4412(1343) ,
  \2623(1167) ,
  \4821(1943) ,
  \4878(1880) ,
  \2713(1178) ,
  \5223(1629) ,
  \4835(1502) ,
  \4683(1362) ,
  \1494(2394) ,
  \5141(1053) ,
  \5045(2289) ,
  \3245(869) ,
  \2699(393) ,
  \4303(1099) ,
  \3254(759) ,
  \589(1711) ,
  \3857(1450) ,
  \840(2451) ,
  \2873(680) ,
  \3959(1466) ,
  \2128(1619) ,
  \1680(615) ,
  \5392(1635) ,
  \5142(1062) ,
  \5186(1085) ,
  \2877(679) ,
  \2159(1621) ,
  \1211(1803) ,
  \4561(1911) ,
  \3529(1767) ,
  \5242(1628) ,
  \2847(656) ,
  \1439(1539) ,
  \2689(391) ,
  \1206(1892) ,
  \798(2028) ,
  \4819(1878) ,
  \1169(1525) ,
  \3914(771) ,
  \4474(1964) ,
  \2897(520) ,
  \856(2029) ,
  \1330(1168) ,
  \3244(758) ,
  \4877(1884) ,
  \1953(1881) ,
  \3250(760) ,
  \4327(1086) ,
  \2278(612) ,
  \3735(2142) ,
  \1674(614) ,
  \3930(1666) ,
  \4311(1093) ,
  \3883(1473) ,
  \3786(808) ,
  \4756(1363) ,
  \5365(775) ,
  \619(1710) ,
  \5296(1127) ,
  \1236(1896) ,
  \3508(1766) ,
  \1246(1906) ,
  \3069(713) ,
  \5375(776) ,
  \2925(875) ,
  \4415(1958) ,
  \3009(856) ,
  \1437(1530) ,
  \4668(1044) ,
  \2893(519) ,
  \1200(1934) ,
  \4698(1851) ,
  \3131(730) ,
  \2756(558) ,
  \3322(597) ,
  \4266(1823) ,
  \3015(863) ,
  \5042(2280) ,
  \5184(1080) ,
  \3334(765) ,
  \4838(2218) ,
  \3135(736) ,
  \3306(594) ,
  \5422(1638) ,
  \2915(873) ,
  \2755(746) ,
  \4903(1517) ,
  \5001(1413) ,
  \2333(2478) ,
  \1177(1524) ,
  \2007(1134) ,
  \1901(1882) ,
  \5244(1966) ,
  \2349(2092) ,
  \2097(1138) ,
  \4829(1855) ,
  \2911(874) ,
  \3410(755) ,
  \570(2001) ,
  \2894(294) ,
  \4242(1341) ,
  \5232(1640) ,
  \2134(1614) ,
  \4893(1500) ,
  \3399(703) ,
  \3640(637) ,
  \5229(1467) ,
  \2154(1617) ,
  \3233(689) ,
  \3395(705) ,
  \2607(669) ,
  \5315(1136) ,
  \2144(1613) ,
  \1203(1891) ,
  \3420(757) ,
  \2890(293) ,
  \5152(1075) ,
  \3083(545) ,
  \4497(1595) ,
  \2751(741) ,
  \3504(1754) ,
  \2611(1159) ,
  \3003(675) ,
  \3543(2120) ,
  \5304(1133) ,
  \1492(2385) ,
  \4896(2217) ,
  \1445(1533) ,
  \5036(2259) ,
  \2762(581) ,
  \771(649) ,
  \1166(1522) ,
  \4434(2263) ,
  \1493(2373) ,
  \4494(2266) ,
  \2145(1620) ,
  \4343(1084) ,
  \2828(206) ,
  \5212(1071) ,
  \3526(1773) ,
  \2153(1618) ,
  \1272(1898) ,
  \4955(1366) ,
  \4376(2264) ,
  \4477(1825) ,
  \5233(1639) ,
  \5222(1634) ,
  \2330(2474) ,
  \2717(1191) ,
  \1199(1865) ,
  \1223(1899) ,
  \2556(580) ,
  \4258(1830) ,
  \2642(555) ,
  \2749(739) ,
  \3956(1465) ,
  \5219(1458) ,
  \1174(1527) ,
  \1444(1531) ,
  \1168(1542) ,
  \3938(1096) ,
  \3126(492) ,
  \4691(1381) ,
  \4578(2160) ,
  \3286(991) ,
  \4927(1379) ,
  \4409(1807) ,
  \4719(1515) ,
  \3348(1043) ,
  \2576(995) ,
  \5396(1110) ,
  \5216(1460) ,
  \4917(1383) ,
  \5347(550) ,
  \2201(2453) ,
  \4247(1553) ,
  \3300(762) ,
  \4429(1560) ,
  \2552(579) ,
  \2929(749) ,
  \4580(2214) ,
  \4887(1854) ,
  \3509(1637) ,
  \2666(458) ,
  \3437(1047) ,
  \3268(292) ,
  \2672(453) ,
  \3283(432) ,
  \761(643) ,
  \705(964) ,
  \4365(1810) ,
  \3963(2107) ,
  \2356(803) ,
  \1216(1999) ,
  \5226(1468) ,
  \1659(2476) ,
  \1251(1903) ,
  \3428(1036) ,
  \3979(374) ,
  \1442(1535) ,
  \1241(1907) ,
  \4954(2204) ,
  \3112(495) ,
  \5059(1496) ,
  \3431(720) ,
  \4791(1049) ,
  \1231(1897) ,
  \3260(295) ,
  \3905(744) ,
  \4472(1836) ,
  \5181(1111) ,
  \1210(1890) ,
  \5312(1145) ,
  \3264(291) ,
  \3065(708) ,
  \2150(1616) ,
  \2595(387) ,
  \1173(1523) ,
  \4202(1814) ,
  \3061(709) ,
  \1524(2454) ,
  \1742(992) ,
  \2113(1632) ,
  \2304(208) ,
  \2065(1124) ,
  \4727(1514) ,
  \3500(1755) ,
  \1947(1941) ,
  \3531(1757) ,
  \[10] ,
  \1483(1895) ,
  \3267(516) ,
  \[11] ,
  \1926(1937) ,
  \2992(969) ,
  \2355(2091) ,
  \3765(371) ,
  \4274(1838) ,
  \[12] ,
  \3047(547) ,
  \3934(1095) ,
  \1171(1526) ,
  \1604(611) ,
  \[13] ,
  \[14] ,
  \5363(576) ,
  \3129(727) ,
  \3512(1768) ,
  \5236(1457) ,
  \2973(423) ,
  \1898(1946) ,
  \[15] ,
  \3967(1769) ,
  \3043(546) ,
  \5252(1976) ,
  \[16] ,
  \3263(523) ,
  \5425(1470) ,
  \[17] ,
  \3326(475) ,
  \5373(588) ,
  \[18] ,
  \1931(1914) ,
  \4172(1087) ,
  \[19] ,
  \3396(892) ,
  \3493(503) ,
  \4491(1833) ,
  \581(2045) ,
  \5335(303) ,
  \3397(1012) ,
  \4210(1812) ,
  \4218(1804) ,
  \5009(1664) ,
  \1916(1940) ,
  \3734(629) ,
  \1440(1534) ,
  \2151(1622) ,
  \2343(2093) ,
  \721(646) ,
  \3514(1057) ,
  \4366(2110) ,
  \3382(333) ,
  \3745(376) ,
  \[20] ,
  \4471(1828) ,
  \2121(1633) ,
  \1481(1528) ,
  \1208(1950) ,
  \5351(319) ,
  \4255(1589) ,
  \4690(1852) ,
  \2898(288) ,
  \2252(2094) ,
  \1238(1953) ,
  \3960(2108) ,
  \1892(1848) ,
  \2968(266) ,
  \5029(1668) ,
  \2939(1144) ,
  \[26] ,
  \1930(1840) ,
  \[27] ,
  \4605(1549) ,
  \[28] ,
  \2964(267) ,
  \1657(2475) ,
  \4820(1879) ,
  \2020(1130) ,
  \3329(702) ,
  \5097(484) ,
  \3086(899) ,
  \3553(198) ,
  \2927(510) ,
  \3505(1636) ,
  \2382(327) ,
  \3929(1786) ,
  \1248(1959) ,
  \3001(395) ,
  \5386(1461) ,
  \857(849) ,
  \2260(603) ,
  \1521(2450) ,
  \4226(1802) ,
  \4346(468) ,
  \2347(2088) ,
  \3056(462) ,
  \5005(1491) ,
  \5243(1459) ,
  \4936(1873) ,
  \5403(1103) ,
  \4019(2137) ,
  \2250(2090) ,
  \[34] ,
  \[35] ,
  \4263(1586) ,
  \2130(1753) ,
  \3869(1447) ,
  \[36] ,
  \2119(1153) ,
  \[37] ,
  \2866(958) ,
  \[38] ,
  \4180(1083) ,
  \1580(605) ,
  \[39] ,
  \3897(935) ,
  \4423(1809) ,
  \2912(990) ,
  \3287(427) ,
  \3338(1003) ,
  \3892(1490) ,
  \3918(1715) ,
  \5359(338) ,
  \3501(1625) ,
  \5085(258) ,
  \3532(1627) ,
  \1888(1924) ,
  \2040(1129) ,
  \711(630) ,
  \4845(1516) ,
  \3066(898) ,
  \3059(1027) ,
  \4581(2161) ,
  \1205(1951) ,
  \4123(443) ,
  \801(642) ,
  \[40] ,
  \2271(790) ,
  \5294(1699) ,
  \3362(344) ,
  \3366(343) ,
  \[41] ,
  \3352(1042) ,
  \[42] ,
  \5369(348) ,
  \2254(606) ,
  \[43] ,
  \1213(1889) ,
  \[44] ,
  \1266(1954) ,
  \791(658) ,
  \[45] ,
  \4643(430) ,
  \4484(2114) ,
  \3347(1002) ,
  \4250(1831) ,
  \[46] ,
  \1921(1939) ,
  \4077(2135) ,
  \3392(879) ,
  \[47] ,
  \1243(1961) ,
  \[48] ,
  \3882(1405) ,
  \2986(972) ,
  \4832(2166) ,
  \3440(284) ,
  \4175(248) ,
  \1662(2477) ,
  \1952(1945) ,
  \5063(1671) ,
  \2281(210) ,
  \1253(1960) ,
  \2353(2089) ,
  \2913(428) ,
  \1847(1509) ,
  \5126(912) ,
  \2976(866) ,
  \[51] ,
  \4667(415) ,
  \[52] ,
  \3167(931) ,
  \[53] ,
  \2574(698) ,
  \3247(417) ,
  \[54] ,
  \3288(693) ,
  \2116(1152) ,
  \[55] ,
  \1701(355) ,
  \[56] ,
  \4322(459) ,
  \4424(2109) ,
  \3881(1402) ,
  \[57] ,
  \4110(298) ,
  \2980(690) ,
  \[58] ,
  \4151(245) ,
  \1855(1507) ,
  \[59] ,
  \1884(1928) ,
  \4716(989) ,
  \4890(2165) ,
  \781(652) ,
  \3933(1785) ,
  \2293(401) ,
  \2948(282) ,
  \3757(181) ,
  \2960(273) ,
  \4812(986) ,
  \4351(1805) ,
  \[60] ,
  \597(1202) ,
  \4271(1570) ,
  \4671(227) ,
  \[61] ,
  \5073(1662) ,
  \4371(1561) ,
  \[62] ,
  \3468(1469) ,
  \4783(921) ,
  \[63] ,
  \5053(1656) ,
  \3477(1471) ,
  \3284(696) ,
  \[64] ,
  \1486(1952) ,
  \3067(1019) ,
  \[65] ,
  \[66] ,
  \[67] ,
  \5173(1104) ,
  \2605(389) ,
  \3416(893) ,
  \2942(1137) ,
  \4083(2130) ,
  \3737(186) ,
  \4025(2129) ,
  \3343(1004) ,
  \4655(231) ,
  \5394(1676) ,
  \2331(798) ,
  \751(659) ,
  \[70] ,
  \[71] ,
  \5162(1100) ,
  \3036(314) ,
  \[72] ,
  \[73] ,
  \3032(315) ,
  \[74] ,
  \5322(932) ,
  \2734(276) ,
  \1467(1596) ,
  \1457(1597) ,
  \3208(281) ,
  \1764(1508) ,
  \[75] ,
  \1271(1955) ,
  \3175(221) ,
  \2166(2399) ,
  \4026(2185) ,
  \[76] ,
  \3556(324) ,
  \[77] ,
  \3204(280) ,
  \[78] ,
  \4340(256) ,
  \5393(1677) ,
  \[79] ,
  \3401(1008) ,
  \3922(1714) ,
  \4119(242) ,
  \5268(1166) ,
  \1178(1559) ,
  \2036(864) ,
  \4022(2136) ,
  \1881(1927) ,
  \1469(1583) ,
  \3777(2209) ,
  \4631(236) ,
  \1179(1552) ,
  \5170(1107) ,
  \2767(936) ,
  \1256(2049) ,
  \3224(264) ,
  \2802(950) ,
  \4559(1827) ,
  \5289(1158) ,
  \1220(1956) ,
  \[80] ,
  \1189(1567) ,
  \3220(265) ,
  \741(651) ,
  \[81] ,
  \3331(1005) ,
  \1288(1328) ,
  \1891(1923) ,
  \3486(1464) ,
  \5206(929) ,
  \[82] ,
  \4639(235) ,
  \[83] ,
  \3085(752) ,
  \5383(1689) ,
  \2122(1151) ,
  \[84] ,
  \2916(985) ,
  \[85] ,
  \4135(238) ,
  \[86] ,
  \[87] ,
  \3075(750) ,
  \1591(789) ,
  \1389(1347) ,
  \[88] ,
  \3071(1030) ,
  \3063(1022) ,
  \[89] ,
  \1181(1590) ,
  \3181(205) ,
  \731(650) ,
  \1086(1554) ,
  \3314(260) ,
  \2882(302) ,
  \3835(2206) ,
  \3137(914) ,
  \5046(2325) ,
  \4194(662) ,
  \1176(1558) ,
  \1845(1226) ,
  \3256(301) ,
  \4080(2134) ,
  \3445(1455) ,
  \3052(304) ,
  \[90] ,
  \3896(740) ,
  \1688(663) ,
  \1806(974) ,
  \[91] ,
  \4308(253) ,
  \4084(2180) ,
  \4876(1315) ,
  \3143(919) ,
  \[92] ,
  \1609(214) ,
  \[93] ,
  \5054(2338) ,
  \1258(2112) ,
  \2990(686) ,
  \[94] ,
  \1579(787) ,
  \[95] ,
  \1468(1572) ,
  \[96] ,
  \2067(1403) ,
  \3861(1444) ,
  \[97] ,
  \5055(2327) ,
  \[98] ,
  \2155(1657) ,
  \1678(2099) ,
  \2914(694) ,
  \4096(2167) ,
  \[99] ,
  \1175(1556) ,
  \3433(918) ,
  \3281(767) ,
  \1585(785) ,
  \2259(784) ,
  \4948(2149) ,
  \2984(687) ,
  \3860(1441) ,
  \2910(695) ,
  \4579(1832) ,
  \1473(1599) ,
  \1466(1577) ,
  \1209(2000) ,
  \3199(639) ,
  \1454(1593) ,
  \1576(2097) ,
  \1456(1578) ,
  \2765(783) ,
  \2265(788) ,
  \3901(1081) ,
  \1447(1565) ,
  \2160(1916) ,
  \3463(1456) ,
  \2687(905) ,
  \3377(578) ,
  \5052(2336) ,
  \3406(883) ,
  \2279(625) ,
  \2933(933) ,
  \3454(1453) ,
  \1465(1584) ,
  \1455(1585) ,
  \2880(684) ,
  \5279(1170) ,
  \3496(725) ,
  \4355(1886) ,
  \4565(1826) ,
  \1475(1579) ,
  \2179(207) ,
  \5276(1154) ,
  \4347(1246) ,
  \1188(1587) ,
  \3373(577) ,
  \5039(1199) ,
  \3236(860) ,
  \3870(1434) ,
  \1446(1564) ,
  \3866(1726) ,
  \4103(1386) ,
  \3325(781) ,
  \2761(774) ,
  \5329(1232) ,
  \3321(780) ,
  \1471(1598) ,
  \2868(681) ,
  \1516(2407) ,
  \4178(1249) ,
  \4931(1842) ,
  \2857(844) ,
  \2662(711) ,
  \2963(490) ,
  \5044(2312) ,
  \3549(200) ,
  \1509(2431) ,
  \2759(773) ,
  \3309(778) ,
  \3910(1088) ,
  \5066(2383) ,
  \3492(726) ,
  \4413(1887) ,
  \1676(2095) ,
  \1172(1557) ,
  \3783(809) ,
  \2135(1673) ,
  \4113(1859) ,
  \5258(2022) ,
  \1515(2408) ,
  \3088(539) ,
  \5149(1217) ,
  \1899(1680) ,
  \1183(1568) ,
  \2663(904) ,
  \1267(2003) ,
  \1472(1580) ,
  \1257(2004) ,
  \5372(782) ,
  \4368(2156) ,
  \1474(1573) ,
  \4730(1317) ,
  \1684(2098) ,
  \3345(769) ,
  \2142(1410) ,
  \1507(2428) ,
  \1508(2435) ,
  \3341(768) ,
  \4099(1240) ,
  \1514(2406) ,
  \1263(2111) ,
  \1513(2405) ,
  \5006(1198) ,
  \2169(2389) ,
  \5101(289) ,
  \1078(1340) ,
  \1519(2445) ,
  \1306(1325) ,
  \1421(1342) ,
  \1277(1333) ,
  \4017(836) ,
  \1856(1513) ,
  \5111(296) ,
  \2042(1408) ,
  \3357(589) ,
  \5307(862) ,
  \1518(2436) ,
  \5148(1221) ,
  \3073(560) ,
  \1192(1569) ,
  \3528(1861) ,
  \1443(1562) ,
  \3405(754) ,
  \3393(994) ,
  \881(370) ,
  \4888(2118) ,
  \4186(1245) ,
  \4487(1743) ,
  \3890(1411) ,
  \3008(676) ,
  \3696(378) ,
  \1482(1575) ,
  \3415(756) ,
  \1331(1336) ,
  \2125(1688) ,
  \4094(527) ,
  \4275(1728) ,
  \1170(1555) ,
  \1682(2096) ,
  \2345(613) ,
  \5159(1230) ,
  \4268(1747) ,
  \3243(498) ,
  \3848(1864) ,
  \1506(2432) ,
  \2351(616) ,
  \5158(1239) ,
  \5064(2370) ,
  \1087(1337) ,
  \1470(1576) ,
  \1854(1512) ,
  \5263(1179) ,
  \2825(204) ,
  \1517(2440) ,
  \3390(435) ,
  \4023(818) ,
  \4746(1782) ,
  \4259(1738) ,
  \4467(1735) ,
  \2165(2378) ,
  \766(644) ,
  \1441(1563) ,
  \5271(1187) ,
  \4331(1248) ,
  \4290(441) ,
  \4426(2155) ,
  \4946(2103) ,
  \1853(1510) ,
  \1895(1681) ,
  \5056(2350) ,
  \1182(1588) ,
  \3525(1863) ,
  \5214(1220) ,
  \1273(2005) ,
  \5065(2359) ,
  \776(632) ,
  \4572(2115) ,
  \3523(1749) ,
  \3432(722) ,
  \3280(522) ,
  \4560(1837) ,
  \3398(445) ,
  \3847(805) ,
  \3018(1126) ,
  \2697(897) ,
  \2099(1419) ,
  \4187(469) ,
  \4419(1702) ,
  \5413(2046) ,
  \2586(704) ,
  \3122(719) ,
  \3422(716) ,
  \2009(1416) ,
  \4684(1759) ,
  \1262(2002) ,
  \1949(2040) ,
  \4267(1736) ,
  \852(255) ,
  \4163(463) ,
  \3253(480) ,
  \3333(473) ,
  \5354(572) ,
  \5260(1182) ,
  \4298(438) ,
  \3394(449) ,
  \2650(549) ,
  \5406(2013) ,
  \4493(2162) ,
  \4998(2416) ,
  \2164(2388) ,
  \1451(1551) ,
  \1132(1346) ,
  \2967(483) ,
  \3027(561) ,
  \4367(2048) ,
  \4754(1781) ,
  \2658(541) ,
  \4825(1761) ,
  \2316(399) ,
  \4889(2060) ,
  \3207(499) ,
  \846(254) ,
  \4009(1287) ,
  \4395(1713) ,
  \3672(380) ,
  \2587(891) ,
  \2988(410) ,
  \2654(542) ,
  \2393(328) ,
  \1850(1511) ,
  \3317(474) ,
  \2584(446) ,
  \790(830) ,
  \5062(2358) ,
  \5215(1233) ,
  \1511(2434) ,
  \3520(1748) ,
  \3336(701) ,
  \1863(1675) ,
  \3227(479) ,
  \4425(2047) ,
  \4251(1720) ,
  \4260(1727) ,
  \1512(2438) ,
  \1477(1600) ,
  \5332(308) ,
  \2750(537) ,
  \4195(1746) ,
  \4433(1724) ,
  \4692(1758) ,
  \3123(478) ,
  \3012(1132) ,
  \5088(477) ,
  \3197(953) ,
  \4794(416) ,
  \1510(2427) ,
  \4676(360) ,
  \5140(1211) ,
  \3632(377) ,
  \4770(434) ,
  \5330(1231) ,
  \2146(1409) ,
  \3660(190) ,
  \4219(1705) ,
  \5250(2016) ,
  \2170(2379) ,
  \1778(1307) ,
  \3403(565) ,
  \3176(362) ,
  \770(838) ,
  \736(633) ,
  \4375(1725) ,
  \3223(481) ,
  \5019(1779) ,
  \4883(1760) ,
  \1476(1601) ,
  \3006(396) ,
  \5414(2018) ,
  \3558(192) ,
  \3413(567) ,
  \726(631) ,
  \4405(1700) ,
  \1021(1332) ,
  \4067(1284) ,
  \2748(535) ,
  \2867(962) ,
  \4778(425) ,
  \780(826) ,
  \3170(1076) ,
  \1934(2039) ,
  \4244(1739) ,
  \4738(1791) ,
  \4147(451) ,
  \806(645) ,
  \796(661) ,
  \3134(521) ,
  \2822(361) ,
  \2997(867) ,
  \3684(188) ,
  \1777(979) ,
  \1268(2050) ,
  \4056(366) ,
  \4276(243) ,
  \2826(364) ,
  \2418(193) ,
  \5193(1244) ,
  \4227(1704) ,
  \3622(372) ,
  \4252(1737) ,
  \3021(1123) ,
  \3733(1868) ,
  \4453(1712) ,
  \4490(2159) ,
  \3297(877) ,
  \3966(1862) ,
  \816(628) ,
  \3237(973) ,
  \1032(1329) ,
  \760(835) ,
  \5192(1247) ,
  \3728(196) ,
  \1661(601) ,
  \2106(1040) ,
  \4015(1289) ,
  \2089(1039) ,
  \4994(2410) ,
  \4830(2119) ,
  \4358(2006) ,
  \2977(980) ,
  \4292(239) ,
  \1578(2101) ,
  \1520(2448) ,
  \2339(600) ,
  \4796(226) ,
  \750(831) ,
  \2798(948) ,
  \5082(262) ,
  \4570(2056) ,
  \2158(1501) ,
  \5013(1783) ,
  \4795(1208) ,
  \2117(1504) ,
  \2918(533) ,
  \4073(1286) ,
  \880(815) ,
  \5024(2036) ,
  \4463(1701) ,
  \4706(1798) ,
  \4666(1209) ,
  \720(848) ,
  \5356(347) ,
  \4803(1205) ,
  \1191(1649) ,
  \3852(1190) ,
  \2794(947) ,
  \1942(2041) ,
  \1887(2021) ,
  \1098(1354) ,
  \5137(922) ,
  \1868(1609) ,
  \4299(1267) ,
  \3234(414) ,
  \730(839) ,
  \2816(353) ,
  \3130(505) ,
  \1050(1324) ,
  \4159(252) ,
  \786(653) ,
  \4416(2007) ,
  \4196(1707) ,
  \5033(1787) ,
  \3391(697) ,
  \4772(232) ,
  \2643(311) ,
  \2647(312) ,
  \1857(1608) ,
  \740(827) ,
  \2975(691) ,
  \1552(213) ,
  \756(660) ,
  \2627(322) ,
  \4815(1794) ,
  \2788(945) ,
  \2780(940) ,
  \4030(183) ,
  \1668(599) ,
  \2131(1493) ,
  \2784(944) ,
  \1983(1321) ,
  \4012(1288) ,
  \4483(2010) ,
  \2553(342) ,
  \4831(2061) ,
  \4204(1706) ,
  \2593(885) ,
  \2557(337) ,
  \4714(1797) ,
  \4810(429) ,
  \2268(2251) ,
  \4934(1784) ,
  \4626(2421) ,
  \4923(1228) ,
  \1195(1605) ,
  \3198(843) ,
  \5072(2392) ,
  \5125(1207) ,
  \3105(278) ,
  \3228(424) ,
  \4945(1788) ,
  \4203(1708) ,
  \4674(1204) ,
  \2163(1969) ,
  \2512(379) ,
  \1792(1303) ,
  \5428(1770) ,
  \1810(1300) ,
  \2810(1078) ,
  \2603(895) ,
  \3925(1815) ,
  \3628(187) ,
  \1666(2035) ,
  \4361(1703) ,
  \1672(2100) ,
  \4873(1799) ,
  \2123(1505) ,
  \4332(247) ,
  \4138(1266) ,
  \1894(2020) ,
  \5124(1206) ,
  \2124(1506) ,
  \1184(1604) ,
  \2936(1072) ,
  \4070(1285) ,
  \646(2269) ,
  \1823(971) ,
  \5225(1762) ,
  \1193(1606) ,
  \4913(1237) ,
  \3949(1843) ,
  \5133(1201) ,
  \4779(1213) ,
  \728(2250) ,
  \746(654) ,
  \4146(1263) ,
  \2721(277) ,
  \3296(763) ,
  \3339(1162) ,
  \4339(1262) ,
  \3846(1982) ,
  \800(834) ,
  \5022(2017) ,
  \1261(2051) ,
  \2276(2253) ,
  \2149(1480) ,
  \4634(1222) ,
  \5077(2441) ,
  \4154(1259) ,
  \4534(2419) ,
  \4544(2418) ,
  \3946(1835) ,
  \595(1463) ,
  \3788(1984) ,
  \3452(1196) ,
  \1502(216) ,
  \4480(2014) ,
  \4627(2446) ,
  \710(822) ,
  \4211(1709) ,
  \3639(2463) ,
  \1114(1351) ,
  \4855(1238) ,
  \5169(1258) ,
  \3203(951) ,
  \2945(1079) ,
  \3780(816) ,
  \2813(977) ,
  \1756(1316) ,
  \1429(1358) ,
  \3238(409) ,
  \1448(1698) ,
  \4018(1290) ,
  \1289(1428) ,
  \1728(1320) ,
  \4532(2413) ,
  \4542(2412) ,
  \3337(886) ,
  \3229(692) ,
  \3836(1120) ,
  \1564(404) ,
  \2147(1476) ,
  \2120(1503) ,
  \4307(1260) ,
  \1878(1647) ,
  \1869(1645) ,
  \1936(2105) ,
  \2238(400) ,
  \2274(2252) ,
  \2540(592) ,
  \3424(913) ,
  \4865(1227) ,
  \4988(2391) ,
  \4013(2027) ,
  \4388(2330) ,
  \4315(1254) ,
  \3658(2460) ,
  \4868(2381) ,
  \1540(406) ,
  \4608(2366) ,
  \4996(2409) ,
  \1190(1603) ,
  \3070(909) ,
  \1686(618) ,
  \4016(2073) ,
  \3843(1983) ,
  \5224(1756) ,
  \[3] ,
  \2500(189) ,
  \4687(1235) ,
  \4682(648) ,
  \[4] ,
  \649(2292) ,
  \3328(916) ,
  \[5] ,
  \1765(1311) ,
  \4071(2026) ,
  \[6] ,
  \4609(1716) ,
  \3649(2458) ,
  \[7] ,
  \[8] ,
  \3785(1985) ,
  \4623(2442) ,
  \577(1967) ,
  \4162(1255) ,
  \[9] ,
  \635(1114) ,
  \3656(2467) ,
  \3943(1834) ,
  \3196(640) ,
  \4078(812) ,
  \3921(1816) ,
  \2691(671) ,
  \4291(1269) ,
  \4997(2390) ,
  \2881(678) ,
  \819(1117) ,
  \3636(2461) ,
  \5235(1772) ,
  \1197(1650) ,
  \1944(2104) ,
  \1596(2258) ,
  \5168(1261) ,
  \4695(1236) ,
  \1584(2146) ,
  \1343(1355) ,
  \2758(569) ,
  \1364(1350) ,
  \4323(1252) ,
  \1867(1481) ,
  \3657(2459) ,
  \4116(1112) ,
  \4279(1113) ,
  \1670(2034) ,
  \5303(1297) ,
  \3058(906) ,
  \4947(2038) ,
  \3645(2464) ,
  \2588(1009) ,
  \4642(1219) ,
  \4170(1251) ,
  \4620(2415) ,
  \1196(1651) ,
  \4397(2345) ,
  \4599(1730) ,
  \3133(732) ,
  \2889(526) ,
  \5176(1268) ,
  \3519(1839) ,
  \4122(1273) ,
  \5234(1771) ,
  \578(1988) ,
  \716(1116) ,
  \4619(1732) ,
  \3239(685) ,
  \2133(1478) ,
  \4828(2043) ,
  \4446(2331) ,
  \5177(1265) ,
  \2869(677) ,
  \2152(1479) ,
  \3782(1986) ,
  \2143(1477) ,
  \3310(595) ,
  \3654(2468) ,
  \4514(2354) ,
  \1874(1646) ,
  \4455(2344) ,
  \3078(553) ,
  \3844(814) ,
  \566(1979) ,
  \3655(2465) ,
  \2270(2254) ,
  \2258(2144) ,
  \4074(2072) ,
  \2708(1352) ,
  \4703(1225) ,
  \5004(2422) ,
  \4540(2426) ,
  \4550(2425) ,
  \1877(1472) ,
  \1194(1652) ,
  \3318(596) ,
  \3653(2466) ,
  \1594(2255) ,
  \2886(297) ,
  \4589(1744) ,
  \3646(636) ,
  \3187(397) ,
  \579(1990) ,
  \1150(1360) ,
  \2908(930) ,
  \3057(712) ,
  \5081(2444) ,
  \3947(1963) ,
  \4568(2015) ,
  \628(1853) ,
  \4650(1212) ,
  \2678(467) ,
  \2764(587) ,
  \3235(688) ,
  \4739(1674) ,
  \2754(551) ,
  \686(2294) ,
  \5116(731) ,
  \637(965) ,
  \4283(1274) ,
  \3332(1163) ,
  \1582(2145) ,
  \3484(1241) ,
  \5106(728) ,
  \3295(515) ,
  \3952(1844) ,
  \1697(357) ,
  \4082(2071) ,
  \703(1115) ,
  \4130(1270) ,
  \1872(1648) ,
  \4944(2037) ,
  \2753(743) ,
  \4024(2068) ,
  \4014(820) ,
  \3642(2462) ,
  \4394(2342) ,
  \5247(1847) ,
  \2638(556) ,
  \2630(563) ,
  \2256(2143) ,
  \2634(564) ,
  \3259(532) ,
  \4711(1224) ,
  \2132(1489) ,
  \713(967) ,
  \5405(1264) ,
  \3731(1121) ,
  \1365(1445) ,
  \5203(1250) ,
  \5074(2414) ,
  \2728(494) ,
  \4523(2364) ,
  \4849(1686) ,
  \1064(996) ,
  \1332(1435) ,
  \2570(999) ,
  \1278(1433) ,
  \4611(2363) ,
  \3147(723) ,
  \4886(2044) ,
  \1843(1630) ,
  \4452(2343) ,
  \4951(1200) ,
  \2747(737) ,
  \4444(2322) ,
  \4918(2356) ,
  \4386(2321) ,
  \3055(538) ,
  \1217(1723) ,
  \1307(1427) ,
  \2226(209) ,
  \1344(1449) ,
  \5026(2102) ,
  \4555(1734) ,
  \3652(2457) ,
  \4811(1218) ,
  \5402(1271) ,
  \5185(1272) ,
  \4020(819) ,
  \4771(1223) ,
  \2660(461) ,
  \5355(559) ,
  \2578(450) ,
  \2564(573) ,
  \4602(2355) ,
  \2041(1304) ,
  \4679(1197) ,
  \1089(1436) ,
  \680(2270) ,
  \683(2291) ,
  \4618(2395) ,
  \5104(514) ,
  \2760(575) ,
  \2548(584) ,
  \4839(1679) ,
  \2560(574) ,
  \3913(745) ,
  \5202(1253) ,
  \4521(1717) ,
  \3944(1962) ,
  \2676(1018) ,
  \4708(1684) ,
  \3128(497) ,
  \5319(1312) ,
  \3051(540) ,
  \1602(2257) ,
  \2544(585) ,
  \4978(2360) ,
  \1116(1446) ,
  \4987(2369) ,
  \1478(1731) ,
  \2664(1026) ,
  \5080(2420) ,
  \1860(1486) ,
  \4111(1765) ,
  \3423(718) ,
  \2350(800) ,
  \4387(2306) ,
  \4976(2351) ,
  \2021(1306) ,
  \1861(1482) ,
  \3271(517) ,
  \4575(1742) ,
  \2999(419) ,
  \3127(724) ,
  \4862(2368) ,
  \4112(1774) ,
  \3937(1256) ,
  \4897(1678) ,
  \652(2293) ,
  \2885(534) ,
  \3092(279) ,
  \5338(543) ,
  \718(1867) ,
  \1526(622) ,
  \1134(1442) ,
  \4520(2365) ,
  \1851(1631) ,
  \1422(1439) ,
  \4524(2387) ,
  \3838(804) ,
  \3948(1919) ,
  \855(1866) ,
  \1915(1790) ,
  \4511(1729) ,
  \3064(454) ,
  \4612(2386) ,
  \4522(2377) ,
  \1870(1483) ,
  \2979(420) ,
  \2202(626) ,
  \4531(1733) ,
  \4445(2307) ,
  \1600(2256) ,
  \785(840) ,
  \5114(530) ,
  \5376(1808) ,
  \1873(1611) ,
  \3202(638) ,
  \4748(1658) ,
  \842(368) ,
  \4079(1119) ,
  \3060(457) ,
  \1597(791) ,
  \5318(1319) ,
  \3522(1845) ,
  \5089(471) ,
  \3533(1846) ,
  \5412(2057) ,
  \3290(984) ,
  \3489(504) ,
  \1592(607) ,
  \3839(1291) ,
  \1390(1443) ,
  \4287(1108) ,
  \3299(507) ,
  \1458(1719) ,
  \5343(313) ,
  \3787(1296) ,
  \3378(334) ,
  \3953(1971) ,
  \2878(961) ,
  \3778(1293) ,
  \1185(1721) ,
  \1606(623) ,
  \2701(673) ,
  \5293(1326) ,
  \4571(2011) ,
  \5014(1841) ,
  \4384(2309) ,
  \5266(1348) ,
  \5267(1345) ,
  \795(833) ,
  \2008(1310) ,
  \1862(1610) ,
  \[100] ,
  \1903(1793) ,
  \[101] ,
  \1318(997) ,
  \3991(179) ,
  \3068(466) ,
  \[102] ,
  \765(847) ,
  \2582(1013) ,
  \4335(1101) ,
  \4364(2053) ,
  \4541(1741) ,
  \4501(1745) ,
  \1929(1751) ,
  \[103] ,
  \1859(1495) ,
  \3276(285) ,
  \[104] ,
  \4533(2398) ,
  \[105] ,
  \3194(954) ,
  \[106] ,
  \4107(1644) ,
  \3551(199) ,
  \4543(2397) ,
  \4155(448) ,
  \[107] ,
  \3462(1210) ,
  \3418(568) ,
  \4860(2357) ,
  \4848(2303) ,
  \2874(959) ,
  \839(2241) ,
  \[108] ,
  \2098(1314) ,
  \4732(1670) ,
  \1128(1025) ,
  \4551(1740) ,
  \[109] ,
  \1667(797) ,
  \3968(1930) ,
  \4723(1683) ,
  \2272(609) ,
  \853(2202) ,
  \2720(1357) ,
  \1871(1612) ,
  \812(2205) ,
  \1586(604) ,
  \3370(339) ,
  \5420(2058) ,
  \1046(1001) ,
  \3536(2059) ,
  \3279(506) ,
  \2370(326) ,
  \1221(1722) ,
  \[110] ,
  \4131(442) ,
  \4442(2308) ,
  \2277(792) ,
  \3970(1978) ,
  \[111] ,
  \1673(794) ,
  \4926(2380) ,
  \4295(1106) ,
  \3272(286) ,
  \[112] ,
  \607(1425) ,
  \1023(1432) ,
  \[113] ,
  \4076(1118) ,
  \3374(340) ,
  \2266(608) ,
  \4610(2376) ,
  \5282(1322) ,
  \3408(566) ,
  \769(2246) ,
  \3275(508) ,
  \[114] ,
  \[115] ,
  \3795(185) ,
  \[116] ,
  \4037(373) ,
  \2870(955) ,
  \4984(2371) ,
  \4968(2326) ,
  \4908(2320) ,
  \580(1991) ,
  \3779(1936) ,
  \709(2245) ,
  \[117] ,
  \5178(934) ,
  \4338(452) ,
  \2670(1023) ,
  \[118] ,
  \[119] ,
  \4986(2382) ,
  \4928(1665) ,
  \1100(1448) ,
  \4552(1194) ,
  \3950(1970) ,
  \878(2242) ,
  \2537(352) ,
  \4763(1659) ,
  \4651(426) ,
  \745(841) ,
  \4314(464) ,
  \1900(1795) ,
  \4966(2318) ,
  \2533(351) ,
  \2901(511) ,
  \4422(2054) ,
  \5093(268) ,
  \3554(331) ,
  \677(2220) ,
  \1359(1029) ,
  \4755(1660) ,
  \[120] ,
  \596(1412) ,
  \4731(1682) ,
  \775(824) ,
  \[121] ,
  \4675(412) ,
  \729(2248) ,
  \[122] ,
  \1866(1407) ,
  \708(2243) ,
  \4659(422) ,
  \3784(1295) ,
  \3941(1257) ,
  \1034(1429) ,
  \608(1440) ,
  \3721(197) ,
  \4530(2396) ,
  \3862(1566) ,
  \1704(1073) ,
  \4482(2055) ,
  \755(832) ,
  \2332(602) ,
  \4139(437) ,
  \3951(1918) ,
  \4330(456) ,
  \5035(2148) ,
  \4635(433) ,
  \1145(1020) ,
  \609(1430) ,
  \1876(1400) ,
  \5283(1338) ,
  \1052(1426) ,
  \768(2244) ,
  \5274(1334) ,
  \2682(1031) ,
  \1453(1718) ,
  \3388(882) ,
  \4700(1685) ,
  \817(2230) ,
  \3803(375) ,
  \2681(911) ,
  \3354(349) ,
  \4977(2339) ,
  \2955(502) ,
  \1080(1438) ,
  \2952(283) ,
  \4920(2367) ,
  \4965(1655) ,
  \5374(949) ,
  \3216(271) ,
  \4124(1109) ,
  \3212(270) ,
  \4919(2348) ,
  \4759(1484) ,
  \2598(880) ,
  \4964(2313) ,
  \2951(501) ,
  \5379(1518) ,
  \4132(1105) ,
  \3823(369) ,
  \2956(272) ,
  \1588(2200) ,
  \3044(310) ,
  \3842(1292) ,
  \805(846) ,
  \1404(1021) ,
  \2264(2199) ,
  \4049(178) ,
  \3781(1294) ,
  \4985(1663) ,
  \643(2221) ,
  \4143(246) ,
  \1412(1033) ,
  \2814(1308) ,
  \3874(1203) ,
  \1978(1068) ,
  \4663(228) ,
  \2608(890) ,
  \3524(1913) ,
  \2592(666) ,
  \3541(2062) ,
  \3878(1367) ,
  \3527(1932) ,
  \814(203) ,
  \5032(2147) ,
  \735(825) ,
  \4907(1687) ,
  \1794(1406) ,
  \3958(1243) ,
  \1324(1017) ,
  \3211(500) ,
  \1031(1006) ,
  \4740(1661) ,
  \4995(1492) ,
  \3518(1371) ,
  \1812(1404) ,
  \2618(1323) ,
  \1896(1796) ,
  \4858(2340) ,
  \1633(212) ,
  \4916(2341) ,
  \4127(241) ,
  \4974(2337) ,
  \724(2247) ,
  \4647(233) ,
  \3535(1921) ,
  \2812(1301) ,
  \4140(1102) ,
  \4975(1672) ,
  \841(813) ,
  \1984(1423) ,
  \1603(793) ,
  \2262(2198) ,
  \725(823) ,
  \5023(1871) ,
  \2018(982) ,
  \3517(1214) ,
  \1966(1067) ,
  \4851(2304) ,
  \3954(1392) ,
  \5302(1302) ,
  \3793(2065) ,
  \1111(1028) ,
  \1724(1066) ,
  \1925(1780) ,
  \723(2249) ,
  \3792(2066) ,
  \3028(321) ,
  \2902(287) ,
  \3851(2063) ,
  \3850(2069) ,
  \3200(952) ,
  \3815(180) ,
  \3024(320) ,
  \1341(1010) ,
  \4316(250) ,
  \3155(924) ,
  \3293(761) ,
  \2905(509) ,
  \3353(1330) ,
  \2115(1229) ,
  \3091(908) ,
  \3165(927) ,
  \1958(1074) ,
  \3515(1372) ,
  \3151(923) ,
  \3361(590) ,
  \3161(926) ,
  \3516(1215) ,
  \3081(900) ,
  \3335(915) ,
  \1712(1065) ,
  \3521(1912) ,
  \1902(1775) ,
  \2909(431) ,
  \3955(1242) ,
  \3791(2067) ,
  \3240(855) ,
  \4941(1669) ,
  \1286(1007) ,
  \4818(1139) ,
  \4069(837) ,
  \3385(570) ,
  \3048(305) ,
  \4909(2305) ,
  \4598(2334) ,
  \3139(917) ,
  \4971(1497) ,
  \1382(1024) ,
  \3302(261) ,
  \3330(887) ,
  \3381(571) ,
  \789(2078) ,
  \4021(1401) ,
  \5195(1391) ,
  \2716(1344) ,
  \5417(1877) ,
  \4081(810) ,
  \574(2158) ,
  \3195(828) ,
  \4910(2329) ,
  \5255(1860) ,
  \4354(1176) ,
  \2203(211) ,
  \1160(1034) ,
  \5310(1309) ,
  \3099(496) ,
  \3040(309) ,
  \1767(1417) ,
  \5295(1536) ,
  \3915(941) ,
  \3945(1908) ,
  \5205(1394) ,
  \4235(1691) ,
  \4406(1177) ,
  \668(2177) ,
  \4398(2362) ,
  \584(2151) ,
  \5194(1390) ,
  \2680(714) ,
  \1645(403) ,
  \2763(777) ,
  \2996(674) ,
  \1097(1011) ,
  \3840(1935) ,
  \4404(2375) ,
  \2696(672) ,
  \2215(402) ,
  \4502(2311) ,
  \4396(2353) ,
  \573(2157) ,
  \3350(1331) ,
  \2253(786) ,
  \4504(2324) ,
  \749(2083) ,
  \2614(1327) ,
  \3193(641) ,
  \2994(394) ,
  \4456(2361) ,
  \5204(1393) ,
  \4075(817) ,
  \4191(1602) ,
  \2808(1318) ,
  \2694(392) ,
  \2876(683) ,
  \4724(1142) ,
  \1758(1420) ,
  \788(2075) ,
  \583(2150) ,
  \5385(1885) ,
  \3853(1356) ,
  \4967(2301) ,
  \2668(710) ,
  \5129(1041) ,
  \2930(872) ,
  \2686(670) ,
  \5311(976) ,
  \2872(682) ,
  \2757(770) ,
  \3313(779) ,
  \5292(1543) ,
  \4751(1485) ,
  \3400(889) ,
  \3513(1216) ,
  \3530(1929) ,
  \3292(531) ,
  \3369(582) ,
  \4628(1063) ,
  \2807(1313) ,
  \4861(2349) ,
  \4243(1690) ,
  \1301(1000) ,
  \4958(2290) ,
  \2684(390) ,
  \799(2080) ,
  \2669(903) ,
  \3547(201) ,
  \4906(2302) ,
  \2907(764) ,
  \5395(1856) ,
  \759(2085) ,
  \1995(993) ,
  \4747(1494) ,
  \4385(1695) ,
  \3230(868) ,
  \3365(583) ,
  \697(2175) ,
  \4762(1454) ,
  \3789(807) ,
  \5364(772) ,
  \811(2219) ,
  \2626(1335) ,
  \4236(1173) ,
  \1590(2201) ,
  \4212(1694) ,
  \1920(1789) ,
  \3004(859) ,
  \1152(1452) ,
  \1621(405) ,
  \3942(1909) ,
  \4513(2332) ,
  \5043(1365) ,
  \5118(1046) ,
  \748(2086) ,
  \4722(1143) ,
  \4592(2323) ,
  \5382(1888) ,
  \2189(2437) ,
  \4470(1193) ,
  \5117(735) ,
  \4228(1015) ,
  \4462(2374) ,
  \1099(1188) ,
  \3957(1389) ,
  \2741(493) ,
  \4852(2328) ,
  \620(1800) ,
  \617(1849) ,
  \4590(2310) ,
  \5107(729) ,
  \5012(1364) ,
  \4636(1060) ,
  \2602(668) ,
  \4234(1174) ,
  \784(2077) ,
  \3201(842) ,
  \4870(1140) ,
  \4220(1693) ,
  \4658(1051) ,
  \700(2176) ,
  \5404(1397) ,
  \4454(2352) ,
  \665(2174) ,
  \2712(1349) ,
  \1698(358) ,
  \794(2079) ,
  \1982(1150) ,
  \5239(1374) ,
  \1198(1778) ,
  \2187(2423) ,
  \694(2172) ,
  \674(2171) ,
  \3643(634) ,
  \3327(766) ,
  \4735(1498) ,
  \590(1806) ,
  \2357(617) ,
  \2188(2433) ,
  \793(2076) ,
  \4898(2261) ,
  \3637(635) ,
  \2838(398) ,
  \2184(2411) ,
  \4443(1697) ,
  \627(1764) ,
  \744(2081) ,
  \1079(1172) ,
  \4562(1965) ,
  \1071(1014) ,
  \4510(2335) ,
  \2183(2417) ,
  \858(647) ,
  \2195(2429) ,
  \2827(620) ,
  \3389(998) ,
  \5105(512) ,
  \2198(2449) ,
  \4011(811) ,
  \783(2074) ,
  \5132(1035) ,
  \4348(1016) ,
  \4377(2213) ,
  \4512(2346) ,
  \5259(1931) ,
  \1685(802) ,
  \2580(706) ,
  \3545(2169) ,
  \2924(748) ,
  \4239(1520) ,
  \753(2087) ,
  \3841(806) ,
  \2185(2424) ,
  \4600(2347) ,
  \4588(2285) ,
  \616(1763) ,
  \2920(747) ,
  \3039(552) ,
  \3035(554) ,
  \743(2082) ,
  \2186(2430) ,
  \4601(2333) ,
  \754(2084) ,
  \1679(801) ,
  \5115(524) ,
  \3849(2024) ,
  \5275(1353) ,
  \2197(2447) ,
  \3537(2019) ,
  \4282(444) ,
  \3118(715) ,
  \2476(191) ,
  \4842(2282) ,
  \1088(1169) ,
  \662(2173) ,
  \3904(742) ,
  \2674(707) ,
  \4644(1055) ,
  \4787(1052) ,
  \4414(1902) ,
  \5346(557) ,
  \1829(1037) ,
  \3594(384) ,
  \5339(536) ,
  \5384(1947) ,
  \2622(1339) ,
  \3120(717) ,
  \4473(1910) ,
  \4850(2319) ,
  \4449(1546) ,
  \3386(439) ,
  \4171(460) ,
  \2590(386) ,
  \1218(1821) ,
  \4356(1901) ,
  \3871(1548) ,
  \4439(1532) ,
  \4459(1538) ,
  \2971(482) ,
  \4775(1056) ,
  \4807(1059) ,
  \3124(721) ,
  \571(2052) ,
  \1730(1422) ,
  \2196(2443) ,
  \4188(363) ,
  \3964(2042) ,
  \640(2170) ,
  \1247(1822) ,
  \4464(1032) ,
  \4179(455) ,
  \1430(1451) ,
  \2194(2439) ,
  \4435(2212) ,
  \2488(381) ,
  \5421(1942) ,
  \4517(1550) ,
  \1428(1192) ,
  \3031(562) ,
  \4374(2211) ,
  \4767(1064) ,
  \3582(194) ,
  \4028(2234) ,
  \3648(2192) ,
  \2568(700) ,
  \3121(472) ,
  \1897(1883) ,
  \2982(413) ;
assign
  \2646(548)  = ~\2643(311) ,
  \4938(1989)  = ~\4937(1938)  | ~\4936(1873) ,
  \1837(1038)  = \3137(914) ,
  \4961(1474)  = \2067(1403) ,
  \3998(367)  = ~\3991(179) ,
  \2752(544)  = \2721(277)  & \280(107) ,
  \2959(489)  = ~\2956(272) ,
  \3249(486)  = \3212(270)  & \3555(332) ,
  \2675(896)  = \2674(707)  | \2672(453) ,
  \3570(382)  = ~\3558(192) ,
  \3449(1624)  = ~\3445(1455) ,
  \4981(1488)  = \2042(1408) ,
  \4582(2265)  = ~\4581(2161)  | ~\4580(2214) ,
  \861(2070)  = \[57] ,
  \615(1750)  = \[46] ,
  \1207(1811)  = ~\4211(1709)  | ~\4204(1706) ,
  \3467(1396)  = ~\5169(1258)  | ~\5162(1100) ,
  \4027(2235)  = \4020(819)  | (\4019(2137)  | \4018(1290) ),
  \5251(1922)  = ~\5247(1847) ,
  \576(1776)  = ~\1878(1647) ,
  \2335(1869)  = \2316(399)  & (\2293(401)  & \3848(1864) ),
  \2581(894)  = \2580(706)  | \2578(450) ,
  \774(2195)  = \3696(378)  & (\3660(190)  & \4026(2185) ),
  \2442(195)  = \4087(171) ,
  \2879(960)  = \2857(844)  & (\2828(206)  & \25(8) ),
  \734(2196)  = \3594(384)  & (\3558(192)  & \4026(2185) ),
  \5362(586)  = ~\5356(347) ,
  \3119(470)  = \3092(279)  & \372(132) ,
  \5121(1048)  = \3143(919) ,
  \2922(518)  = \2890(293)  & \3554(331) ,
  \298(299)  = \293(112) ,
  \3132(513)  = \3105(278)  & \315(117) ,
  \4786(421)  = ~\4780(230) ,
  \3540(2164)  = ~\3538(2117) ,
  \1849(1148)  = \1742(992)  & \1712(1065) ,
  \4068(1980)  = \4056(366)  & (\4030(183)  & \1916(1940) ),
  \5034(2203)  = ~\5032(2147)  | ~\5029(1668) ,
  \3125(485)  = \3092(279)  & \348(126) ,
  \4956(2267)  = ~\4954(2204)  | ~\4951(1200) ,
  \3476(1399)  = ~\5177(1265)  | ~\5170(1107) ,
  \2811(1298)  = ~\3021(1123) ,
  \1224(1777)  = \4(1)  & \1179(1552) ,
  \773(2194)  = \3696(378)  & (\3672(380)  & \4084(2180) ),
  \5340(318)  = \265(104) ,
  \2906(525)  = \2886(297)  & \2393(328) ,
  \1237(1818)  = ~\4251(1720)  | ~\4244(1739) ,
  \5331(1387)  = ~\5329(1232)  | ~\5322(932) ,
  \733(2197)  = \3594(384)  & (\3570(382)  & \4084(2180) ),
  \2875(956)  = \2857(844)  & (\2828(206)  & \81(29) ),
  \807(2480)  = \[120] ,
  \3965(2153)  = ~\3964(2042)  | ~\3963(2107) ,
  \5366(598)  = \2816(353) ,
  \633(365)  = ~\1(0)  | ~\373(133) ,
  \767(2479)  = \[119] ,
  \2809(1234)  = ~\2936(1072) ,
  \4507(1571)  = \1390(1443) ,
  \2871(957)  = \2857(844)  & (\2828(206)  & \80(28) ),
  \4503(2288)  = ~\4501(1745)  | ~\4494(2266) ,
  \4086(2231)  = \4081(810)  | (\4080(2134)  | \4079(1119) ),
  \2361(325)  = \254(101) ,
  \5285(1424)  = ~\5283(1338)  | ~\5276(1154) ,
  \4481(1904)  = ~\4477(1825) ,
  \2454(385)  = ~\2442(195) ,
  \3475(1398)  = ~\5176(1268)  | ~\5173(1104) ,
  \3358(350)  = \210(89) ,
  \5096(491)  = ~\5090(274) ,
  \4207(1545)  = \1023(1432) ,
  \3497(1626)  = \3463(1456) ,
  \1889(1850)  = ~\4707(1377)  | ~\4700(1685) ,
  \1660(799)  = \1633(212)  & (\1621(405)  & \176(77) ),
  \4199(1544)  = \1023(1432) ,
  \4432(2210)  = ~\4426(2155) ,
  \4991(1414)  = \2021(1306) ,
  \1948(1993)  = \1898(1946)  & \1903(1793) ,
  \3466(1395)  = ~\5168(1261)  | ~\5165(1097) ,
  \3891(1305)  = ~\5311(976)  | ~\5304(1133) ,
  \1729(1146)  = ~\4635(433)  | ~\4628(1063) ,
  \1287(1160)  = ~\4290(441)  | ~\4287(1108) ,
  \3305(476)  = ~\3302(261) ,
  \5108(300)  = \293(112) ,
  \4840(2262)  = ~\4838(2218)  | ~\4835(1502) ,
  \2337(2033)  = \2316(399)  & (\2281(210)  & \3790(2025) ),
  \5196(1092)  = \2780(940) ,
  \600(259)  = \[5] ,
  \4660(1050)  = \3143(919) ,
  \4284(240)  = \457(142) ,
  \5348(335)  = \234(95) ,
  \2572(436)  = \2545(345)  & (\468(143)  & \3553(198) ),
  \1151(1195)  = ~\4187(469)  | ~\4180(1083) ,
  \3542(2023)  = ~\5259(1931)  | ~\5252(1976) ,
  \5165(1097)  = \2784(944) ,
  \5151(1375)  = ~\5149(1217)  | ~\5142(1062) ,
  \3215(487)  = ~\3212(270) ,
  \2566(440)  = \2537(352)  & (\457(142)  & \3553(198) ),
  \4492(2215)  = ~\4490(2159)  | ~\4487(1743) ,
  \1388(1181)  = ~\4330(456)  | ~\4327(1086) ,
  \3219(488)  = ~\3216(271) ,
  \1033(1161)  = ~\4131(442)  | ~\4124(1109) ,
  \4899(2207)  = ~\4897(1678)  | ~\4890(2165) ,
  \3136(529)  = \3105(278)  & \299(113) ,
  \4591(2287)  = ~\4589(1744)  | ~\4582(2265) ,
  \4527(1582)  = \1365(1445) ,
  \4085(2232)  = \4078(812)  | (\4077(2135)  | \4076(1118) ),
  \779(2139)  = \3696(378)  & (\3660(190)  & \4025(2129) ),
  \1225(1819)  = \1224(1777)  | \1185(1721) ,
  \1776(1131)  = ~\4658(1051)  | ~\4655(231) ,
  \5399(946)  = ~\5365(775)  | ~\5364(772) ,
  \3837(1653)  = \3823(369)  & (\3795(185)  & \1878(1647) ),
  \3555(332)  = \242(97) ,
  \3289(871)  = \3288(693)  | \3287(427) ,
  \5150(1373)  = ~\5148(1221)  | ~\5145(1058) ,
  \1204(1813)  = ~\4203(1708)  | ~\4196(1707) ,
  \3485(1388)  = ~\5185(1272)  | ~\5178(934) ,
  \2081(970)  = \3139(917)  & \534(149) ,
  \1022(1164)  = ~\4123(443)  | ~\4116(1112) ,
  \1276(1165)  = ~\4282(444)  | ~\4279(1113) ,
  \3458(1607)  = ~\3454(1453) ,
  \1766(1135)  = ~\4651(426)  | ~\4644(1055) ,
  \1846(1147)  = \1742(992)  & (\1704(1073)  & \1712(1065) ),
  \689(2482)  = \2279(625)  & \2333(2478) ,
  \1222(1820)  = ~\4243(1690)  | ~\4236(1173) ,
  \1757(1141)  = ~\4643(430)  | ~\4636(1060) ,
  \4183(257)  = \374(134) ,
  \4935(1917)  = ~\4931(1842) ,
  \2430(383)  = ~\2418(193) ,
  \5161(1385)  = ~\5159(1230)  | ~\5152(1075) ,
  \4215(1541)  = \1034(1429) ,
  \4615(1581)  = \1365(1445) ,
  \778(2138)  = \3696(378)  & (\3672(380)  & \4083(2130) ),
  \3472(1641)  = ~\3468(1469) ,
  \659(2121)  = \1668(599)  | (\1667(797)  | (\1666(2035)  | \1664(1870) )),
  \3887(1654)  = ~\3883(1473) ,
  \4822(1995)  = ~\4821(1943)  | ~\4820(1879) ,
  \3972(184)  = \4091(175) ,
  \3285(876)  = \3284(696)  | \3283(432) ,
  \4780(230)  = \514(147) ,
  \2991(857)  = \2990(686)  | \2988(410) ,
  \4595(1574)  = \1390(1443) ,
  \4957(2216)  = ~\4955(1366)  | ~\4948(2149) ,
  \1242(1829)  = ~\4259(1738)  | ~\4252(1737) ,
  \658(2483)  = \[121] ,
  \3962(2154)  = ~\3961(2116)  | ~\3960(2108) ,
  \5090(274)  = \341(125) ,
  \4500(2286)  = ~\4494(2266) ,
  \1252(1824)  = ~\4275(1728)  | ~\4268(1747) ,
  \4569(1905)  = ~\4565(1826) ,
  \4537(1592)  = \1344(1449) ,
  \4788(229)  = \523(148) ,
  \5286(1431)  = \3350(1331) ,
  \4231(1521)  = \1052(1426) ,
  \5160(1380)  = ~\5158(1239)  | ~\5155(1069) ,
  \4937(1938)  = ~\4935(1917)  | ~\4928(1665) ,
  \4547(1591)  = \1344(1449) ,
  \1935(1994)  = \1883(1974)  & \1903(1793) ,
  \739(2140)  = \3594(384)  & (\3558(192)  & \4025(2129) ),
  \1885(1858)  = ~\4699(1382)  | ~\4692(1758) ,
  \2344(795)  = \2304(208)  & (\2293(401)  & \188(81) ),
  \764(2471)  = \2454(385)  & (\2418(193)  & \3655(2465) ),
  \2985(858)  = \2984(687)  | \2982(413) ,
  \4167(251)  = \400(137) ,
  \879(2452)  = \3765(371)  & (\3737(186)  & \1521(2450) ),
  \657(2481)  = \1606(623)  & \1662(2477) ,
  \4148(1098)  = \2784(944) ,
  \2639(316)  = \265(104) ,
  \2631(323)  = \257(102) ,
  \1775(983)  = \503(146)  & \3151(923) ,
  \4764(237)  = \479(144) ,
  \3481(1643)  = ~\3477(1471) ,
  \1789(865)  = \514(147)  & \3147(723) ,
  \5429(1642)  = ~\5425(1470) ,
  \2635(317)  = \265(104) ,
  \1051(1156)  = ~\4139(437)  | ~\4132(1105) ,
  \3231(981)  = ~\3230(868) ,
  \859(2132)  = \[63] ,
  \804(2470)  = \2512(379)  & (\2476(191)  & \3655(2465) ),
  \1919(1874)  = ~\4746(1782)  | ~\4743(1415) ,
  \5015(1915)  = ~\5013(1783)  | ~\5006(1198) ,
  \4306(447)  = ~\4300(244) ,
  \4879(1944)  = ~\4877(1884)  | ~\4870(1140) ,
  \1954(1997)  = \1953(1881)  | \1952(1945) ,
  \2561(336)  = \234(95) ,
  \4223(1540)  = \1034(1429) ,
  \738(2141)  = \3594(384)  & (\3570(382)  & \4083(2130) ),
  \5284(1437)  = ~\5282(1322)  | ~\5279(1170) ,
  \3387(699)  = \3361(590)  & (\2370(326)  & \457(142) ),
  \2059(975)  = \3143(919)  & \523(148) ,
  \4391(1547)  = \1278(1433) ,
  \4880(1996)  = ~\4879(1944)  | ~\4878(1880) ,
  \3232(418)  = \514(147)  & \2405(329) ,
  \763(2472)  = \2454(385)  & (\2430(383)  & \3656(2467) ),
  \2541(346)  = \218(91) ,
  \4104(1462)  = \4103(1386)  | \4099(1240) ,
  \1852(1149)  = \1742(992)  & \1712(1065) ,
  \1886(1975)  = ~\1885(1858)  | ~\1884(1928) ,
  \1909(1876)  = ~\1903(1793) ,
  \4401(1537)  = \1289(1428) ,
  \5098(290)  = \308(116) ,
  \1749(988)  = \3155(924)  & \490(145) ,
  \4558(1359)  = ~\4552(1194) ,
  \4859(1384)  = ~\4855(1238) ,
  \3651(2193)  = \3632(377)  & \3965(2153) ,
  \5328(1077)  = ~\5322(932) ,
  \1664(1870)  = \1645(403)  & (\1621(405)  & \3848(1864) ),
  \4319(1091)  = \2776(939) ,
  \2549(341)  = \226(93) ,
  \2338(796)  = \2304(208)  & (\2293(401)  & \182(79) ),
  \2597(667)  = \2544(585)  & \3549(200) ,
  \2600(388)  = \2549(341)  & \3547(201) ,
  \2066(1299)  = ~\4803(1205)  | ~\4796(226) ,
  \1943(1992)  = \1890(1973)  & \1903(1793) ,
  \1305(1157)  = ~\4298(438)  | ~\4295(1106) ,
  \4869(1378)  = ~\4865(1227) ,
  \568(2008)  = ~\1248(1959) ,
  \4156(1094)  = \2780(940) ,
  \2193(2403)  = \2174(161)  & (\2163(1969)  & \2166(2399) ),
  \2709(1183)  = \2692(902)  & \2670(1023) ,
  \2545(345)  = \218(91) ,
  \4585(1594)  = \1430(1451) ,
  \2776(939)  = \2754(551)  | \2753(743) ,
  \3346(943)  = \3321(780)  & \2361(325) ,
  \5209(925)  = ~\5107(729)  | ~\5106(728) ,
  \1462(1817)  = ~\1458(1719) ,
  \3342(942)  = \3309(778)  & \2361(325) ,
  \1882(1857)  = ~\4691(1381)  | ~\4684(1759) ,
  \3926(1667)  = \3892(1490) ,
  \2575(881)  = \2574(698)  | \2572(436) ,
  \4010(1981)  = \3998(367)  & (\3972(184)  & \1238(1953) ),
  \2772(937)  = \2752(544)  | \2751(741) ,
  \844(657)  = \27(10)  & \2825(204) ,
  \1115(1185)  = ~\4171(460)  | ~\4164(1090) ,
  \2405(329)  = \248(99) ,
  \719(2030)  = \2454(385)  & (\2418(193)  & \3790(2025) ),
  \2341(2032)  = \2316(399)  & (\2293(401)  & \3849(2024) ),
  \1363(1184)  = ~\4322(459)  | ~\4319(1091) ,
  \567(2009)  = ~\1253(1960) ,
  \3895(738)  = ~\5338(543)  | ~\5335(303) ,
  \5025(1987)  = ~\5023(1871)  | ~\5016(1968) ,
  \877(2126)  = \[67] ,
  \1489(2393)  = ~\1488(2372)  | ~\1487(2384) ,
  \4743(1415)  = \1778(1307) ,
  \3282(928)  = \3281(767)  | \3280(522) ,
  \3845(963)  = \3823(369)  & (\3803(375)  & \3015(863) ),
  \4707(1377)  = ~\4703(1225) ,
  \3790(2025)  = \3780(816)  | (\3779(1936)  | \3778(1293) ),
  \3090(753)  = \3051(540)  & \3556(324) ,
  \4114(359)  = \4115(177)  & \135(61) ,
  \3444(1368)  = ~\5125(1207)  | ~\5118(1046) ,
  \5069(1487)  = \2042(1408) ,
  \2192(2404)  = \2174(161)  & (\2160(1916)  & \2171(2400) ),
  \5409(1998)  = ~\5385(1885)  | ~\5384(1947) ,
  \3241(968)  = ~\3240(855) ,
  \582(2106)  = ~\1949(2040) ,
  \634(665)  = \[17] ,
  \4381(1529)  = \1307(1427) ,
  \1528(215)  = \1689(157) ,
  \2139(1792)  = ~\2135(1673) ,
  \4324(249)  = \411(138) ,
  \569(2012)  = ~\1243(1961) ,
  \3080(751)  = \3035(554)  & \3556(324) ,
  \1342(1189)  = ~\4314(464)  | ~\4311(1093) ,
  \803(2469)  = \2512(379)  & (\2488(381)  & \3656(2467) ),
  \1893(1972)  = ~\1892(1848)  | ~\1891(1923) ,
  \2569(884)  = \2568(700)  | \2566(440) ,
  \4164(1090)  = \2776(939) ,
  \2766(593)  = \2734(276)  & \209(88) ,
  \1215(1948)  = ~\1214(1801)  | ~\1213(1889) ,
  \4699(1382)  = ~\4695(1236) ,
  \3255(854)  = \534(149)  | (\3254(759)  | \3253(480) ),
  \4652(920)  = \3147(723) ,
  \3453(1361)  = ~\5133(1201)  | ~\5126(912) ,
  \5325(1070)  = ~\3282(928) ,
  \5321(1421)  = ~\5319(1312)  | ~\5312(1145) ,
  \2191(2402)  = \2179(207)  & (\2135(1673)  & \2166(2399) ),
  \2171(2400)  = ~\2170(2379)  | ~\2169(2389) ,
  \3443(1369)  = ~\5124(1206)  | ~\5121(1048) ,
  \2328(2473)  = \2316(399)  & (\2293(401)  & \3654(2468) ),
  \1883(1974)  = ~\1882(1857)  | ~\1881(1927) ,
  \4900(2281)  = ~\4899(2207)  | ~\4898(2261) ,
  \758(2031)  = \2454(385)  & (\2430(383)  & \3849(2024) ),
  \5134(1054)  = \3151(923) ,
  \5320(1418)  = ~\5318(1319)  | ~\5315(1136) ,
  \843(2455)  = \[117] ,
  \3461(1370)  = ~\5140(1211)  | ~\5137(922) ,
  \4300(244)  = \435(140) ,
  \4357(1957)  = ~\4355(1886)  | ~\4348(1016) ,
  \1420(1175)  = ~\4338(452)  | ~\4335(1101) ,
  \5145(1058)  = \3155(924) ,
  \5199(1089)  = \2776(939) ,
  \4802(411)  = ~\4796(226) ,
  \3616(182)  = \4092(176) ,
  \5049(1475)  = \2067(1403) ,
  \836(2128)  = \[62] ,
  \1133(1180)  = ~\4179(455)  | ~\4172(1087) ,
  \3961(2116)  = ~\5413(2046)  | ~\5406(2013) ,
  \1793(1128)  = ~\4667(415)  | ~\4660(1050) ,
  \3906(938)  = ~\3905(744)  | ~\3904(742) ,
  \722(2131)  = \[59] ,
  \5155(1069)  = \3165(927) ,
  \2019(978)  = ~\4786(421)  | ~\4783(921) ,
  \5016(1968)  = ~\5015(1915)  | ~\5014(1841) ,
  \1811(1125)  = ~\4675(412)  | ~\4668(1044) ,
  \1924(1872)  = ~\4754(1781)  | ~\4751(1485) ,
  \4715(1376)  = ~\4711(1224) ,
  \2001(987)  = \3155(924)  & \490(145) ,
  \1219(1900)  = ~\1218(1821)  | ~\1217(1723) ,
  \1914(1875)  = ~\4738(1791)  | ~\4735(1498) ,
  \2619(1171)  = \2603(895)  & \2582(1013) ,
  \5189(1082)  = \2767(936) ,
  \4072(821)  = \4049(178)  & (\4037(373)  & \112(42) ),
  \3538(2117)  = ~\3537(2019)  | ~\3536(2059) ,
  \882(2456)  = \[118] ,
  \1875(1279)  = \1829(1037)  & \54(20) ,
  \2190(2401)  = \2179(207)  & (\2139(1792)  & \2171(2400) ),
  \1214(1801)  = ~\4227(1704)  | ~\4220(1693) ,
  \2615(1155)  = \2598(880)  & \2576(995) ,
  \707(1277)  = \[41] ,
  \671(966)  = \2877(679)  | (\2876(683)  | (\2875(956)  | \2874(959) )),
  \875(2125)  = \[66] ,
  \834(2123)  = \[61] ,
  \5213(1061)  = ~\5209(925) ,
  \572(2113)  = ~\1268(2050) ,
  \3411(878)  = \468(143)  | (\3410(755)  | \3408(566) ),
  \3251(861)  = \523(148)  | (\3250(760)  | \3249(486) ),
  \2655(306)  = \281(108) ,
  \1598(610)  = \1552(213)  & (\1528(215)  & \164(73) ),
  \4841(2208)  = ~\4839(1679)  | ~\4832(2166) ,
  \3301(870)  = \490(145)  | (\3300(762)  | \3299(507) ),
  \2651(307)  = \281(108) ,
  \3076(907)  = \389(136)  | (\3075(750)  | \3073(560) ),
  \5299(1122)  = \3255(854)  & \3241(968) ,
  \691(2122)  = \2339(600)  | (\2338(796)  | (\2337(2033)  | \2335(1869) )),
  \1487(2384)  = ~\4404(2375)  | ~\4401(1537) ,
  \5389(1499)  = ~\5321(1421)  | ~\5320(1418) ,
  \4436(2283)  = ~\4435(2212)  | ~\4434(2263) ,
  \2692(902)  = \400(137)  | (\2691(671)  | \2689(391) ),
  \832(2133)  = \[60] ,
  \2536(591)  = ~\2533(351) ,
  \717(1282)  = \[37] ,
  \2148(1615)  = \2021(1306)  & (\2089(1039)  & (\2042(1408)  & \2067(1403) )),
  \3192(829)  = \3187(397)  & \83(31) ,
  \3062(901)  = \3061(709)  | \3060(457) ,
  \4799(1045)  = \3139(917) ,
  \3421(888)  = \435(140)  | (\3420(757)  | \3418(568) ),
  \2705(1186)  = \2687(905)  & \2664(1026) ,
  \690(2484)  = \[122] ,
  \4378(2284)  = ~\4377(2213)  | ~\4376(2264) ,
  \1890(1973)  = ~\1889(1850)  | ~\1888(1924) ,
  \1212(1949)  = ~\1211(1803)  | ~\1210(1890) ,
  \4804(234)  = \490(145) ,
  \1488(2372)  = ~\4405(1700)  | ~\4398(2362) ,
  \2702(910)  = \374(134)  | (\2701(673)  | \2699(393) ),
  \4412(1343)  = ~\4406(1177) ,
  \2623(1167)  = \2608(890)  & \2588(1009) ,
  \4821(1943)  = ~\4819(1878)  | ~\4812(986) ,
  \4878(1880)  = ~\4876(1315)  | ~\4873(1799) ,
  \2713(1178)  = \2697(897)  & \2676(1018) ,
  \5223(1629)  = ~\5219(1458) ,
  \4835(1502)  = \2099(1419) ,
  \4683(1362)  = ~\4679(1197) ,
  \1494(2394)  = ~\1493(2373)  | ~\1492(2385) ,
  \5141(1053)  = ~\5137(922) ,
  \5045(2289)  = ~\5043(1365)  | ~\5036(2259) ,
  \3245(869)  = \503(146)  | (\3244(758)  | \3243(498) ),
  \2699(393)  = \2651(307)  & \3547(201) ,
  \4303(1099)  = \2784(944) ,
  \3254(759)  = \3223(481)  & \2361(325) ,
  \589(1711)  = \1441(1563)  | (\1440(1534)  | (\1439(1539)  | \1286(1007) )),
  \3857(1450)  = ~\3853(1356) ,
  \840(2451)  = \3823(369)  & (\3795(185)  & \2198(2449) ),
  \639(1275)  = \[39] ,
  \2873(680)  = \2847(656)  & \2828(206) ,
  \3959(1466)  = ~\3958(1243)  & ~\3957(1389) ,
  \873(2124)  = \[65] ,
  \851(218)  = \[16] ,
  \2128(1619)  = \2009(1416)  & (\2021(1306)  & (\2042(1408)  & (\2067(1403)  & \2106(1040) ))),
  \1680(615)  = \1633(212)  & (\1609(214)  & \152(69) ),
  \5392(1635)  = ~\5386(1461) ,
  \5142(1062)  = \3161(926) ,
  \5186(1085)  = \2772(937) ,
  \2877(679)  = \2847(656)  & \2828(206) ,
  \2159(1621)  = \2067(1403)  & \2106(1040) ,
  \1211(1803)  = ~\4219(1705)  | ~\4212(1694) ,
  \599(269)  = \[4] ,
  \4561(1911)  = ~\4559(1827)  | ~\4552(1194) ,
  \849(219)  = \[14] ,
  \3529(1767)  = \3509(1637)  & (\3472(1641)  & \3481(1643) ),
  \5242(1628)  = ~\5236(1457) ,
  \715(1278)  = \[42] ,
  \2847(656)  = ~\2822(361) ,
  \1439(1539)  = \1301(1000)  & \1278(1433) ,
  \2689(391)  = \2635(317)  & \3547(201) ,
  \1206(1892)  = ~\4210(1812)  | ~\4207(1545) ,
  \798(2028)  = \2512(379)  & (\2488(381)  & \3849(2024) ),
  \4819(1878)  = ~\4815(1794) ,
  \1169(1525)  = \1064(996)  & (\1023(1432)  & \1034(1429) ),
  \3914(771)  = ~\5355(559)  | ~\5348(335) ,
  \4474(1964)  = ~\4473(1910)  | ~\4472(1836) ,
  \2897(520)  = ~\2894(294) ,
  \856(2029)  = \2512(379)  & (\2476(191)  & \3790(2025) ),
  \1330(1168)  = ~\4306(447)  | ~\4303(1099) ,
  \848(330)  = \[13] ,
  \3244(758)  = \3207(499)  & \2361(325) ,
  \4877(1884)  = ~\4873(1799) ,
  \1953(1881)  = \1764(1508)  & \1903(1793) ,
  \3250(760)  = \3215(487)  & \2361(325) ,
  \4327(1086)  = \2772(937) ,
  \2278(612)  = \2226(209)  & (\2203(211)  & \161(72) ),
  \3735(2142)  = \3717(169)  & (\3724(170)  & \1936(2105) ),
  \1674(614)  = \1633(212)  & (\1609(214)  & \158(71) ),
  \3930(1666)  = \3892(1490) ,
  \4311(1093)  = \2780(940) ,
  \3883(1473)  = ~\3882(1405)  | ~\3881(1402) ,
  \3786(808)  = \3757(181)  & (\3745(376)  & \127(55) ),
  \871(2127)  = \[64] ,
  \4756(1363)  = \1875(1279)  | \1837(1038) ,
  \5365(775)  = ~\5363(576)  | ~\5356(347) ,
  \619(1710)  = \1170(1555)  | (\1169(1525)  | (\1168(1542)  | \1031(1006) )),
  \5296(1127)  = \3251(861)  & \3237(973) ,
  \1236(1896)  = ~\4250(1831)  | ~\4247(1553) ,
  \3508(1766)  = ~\3505(1636) ,
  \1246(1906)  = ~\4266(1823)  | ~\4263(1586) ,
  \3069(713)  = \3055(538)  & (\2370(326)  & \374(134) ),
  \5375(776)  = ~\5373(588)  | ~\5366(598) ,
  \2925(875)  = \479(144)  | (\2924(748)  | \2922(518) ),
  \4415(1958)  = ~\4413(1887)  | ~\4406(1177) ,
  \636(1280)  = \[35] ,
  \3009(856)  = \534(149)  | (\3008(676)  | \3006(396) ),
  \704(1281)  = \[36] ,
  \1437(1530)  = \1278(1433)  & (\1289(1428)  & (\1307(1427)  & \1422(1439) )),
  \4668(1044)  = \3139(917) ,
  \2893(519)  = ~\2890(293) ,
  \1200(1934)  = ~\1199(1865)  | ~\1198(1778) ,
  \4698(1851)  = ~\4692(1758) ,
  \3131(730)  = \3112(495)  & \308(116) ,
  \2756(558)  = \2721(277)  & \264(103) ,
  \3322(597)  = \2816(353) ,
  \4266(1823)  = ~\4260(1727) ,
  \3015(863)  = \2999(419)  & \2980(690) ,
  \5042(2280)  = ~\5036(2259) ,
  \5184(1080)  = ~\5178(934) ,
  \3334(765)  = \3317(474)  & \2382(327) ,
  \4838(2218)  = ~\4832(2166) ,
  \3135(736)  = \3112(495)  & \293(112) ,
  \3306(594)  = \2816(353) ,
  \5422(1638)  = ~\3956(1465)  | ~\3959(1466) ,
  \2915(873)  = \2914(694)  | \2913(428) ,
  \2755(746)  = \2728(494)  & \257(102) ,
  \4903(1517)  = \1984(1423) ,
  \5001(1413)  = \2021(1306) ,
  \2333(2478)  = \2332(602)  | (\2331(798)  | (\2330(2474)  | \2328(2473) )),
  \1177(1524)  = \1052(1426)  & \1080(1438) ,
  \2007(1134)  = ~\4778(425)  | ~\4775(1056) ,
  \1901(1882)  = ~\1900(1795)  | ~\1899(1680) ,
  \5244(1966)  = ~\3521(1912)  | ~\3524(1913) ,
  \2349(2092)  = \2316(399)  & (\2281(210)  & \3792(2066) ),
  \2097(1138)  = ~\4810(429)  | ~\4807(1059) ,
  \4829(1855)  = ~\4825(1761) ,
  \2911(874)  = \2910(695)  | \2909(431) ,
  \3410(755)  = \3365(583)  & \3556(324) ,
  \570(2001)  = ~\1238(1953) ,
  \2894(294)  = \308(116) ,
  \4242(1341)  = ~\4236(1173) ,
  \5232(1640)  = ~\5226(1468) ,
  \2134(1614)  = \2021(1306)  & (\2089(1039)  & (\2009(1416)  & (\2042(1408)  & \2067(1403) ))),
  \4893(1500)  = \2099(1419) ,
  \3399(703)  = \3385(570)  & (\2370(326)  & \435(140) ),
  \3640(637)  = \3616(182)  & \94(36) ,
  \5229(1467)  = ~\5195(1391)  | ~\5194(1390) ,
  \2154(1617)  = \2089(1039)  & \2067(1403) ,
  \3233(689)  = ~\3232(418) ,
  \3395(705)  = \3377(578)  & (\2370(326)  & \422(139) ),
  \2607(669)  = \2560(574)  & \3549(200) ,
  \5315(1136)  = \3301(870)  & \3290(984) ,
  \2144(1613)  = \2021(1306)  & (\2089(1039)  & (\2042(1408)  & \2067(1403) )),
  \1203(1891)  = ~\4202(1814)  | ~\4199(1544) ,
  \3420(757)  = \3381(571)  & \3556(324) ,
  \2890(293)  = \308(116) ,
  \5152(1075)  = \3167(931) ,
  \3083(545)  = \3040(309)  & \3554(331) ,
  \4497(1595)  = \1430(1451) ,
  \2751(741)  = \2728(494)  & \273(106) ,
  \3504(1754)  = ~\3501(1625) ,
  \2611(1159)  = \2593(885)  & \2570(999) ,
  \3003(675)  = \2959(489)  & \3549(200) ,
  \3543(2120)  = ~\3542(2023)  | ~\3541(2062) ,
  \5304(1133)  = \3245(869)  & \3231(981) ,
  \1492(2385)  = ~\4462(2374)  | ~\4459(1538) ,
  \4896(2217)  = ~\4890(2165) ,
  \1445(1533)  = \1318(997)  & \1289(1428) ,
  \5036(2259)  = ~\5035(2148)  | ~\5034(2203) ,
  \2762(581)  = \2734(276)  & \225(92) ,
  \771(649)  = \3684(188)  & (\3660(190)  & \49(17) ),
  \1166(1522)  = \1023(1432)  & (\1052(1426)  & (\1080(1438)  & \1034(1429) )),
  \4434(2263)  = ~\4432(2210)  | ~\4429(1560) ,
  \1493(2373)  = ~\4463(1701)  | ~\4456(2361) ,
  \4494(2266)  = ~\4493(2162)  | ~\4492(2215) ,
  \2145(1620)  = \2067(1403)  & (\2021(1306)  & (\2042(1408)  & \2106(1040) )),
  \4343(1084)  = \2767(936) ,
  \2828(206)  = \2358(162) ,
  \5212(1071)  = ~\5206(929) ,
  \3526(1773)  = \3505(1636)  & (\3468(1469)  & \3477(1471) ),
  \2153(1618)  = \2089(1039)  & (\2042(1408)  & \2067(1403) ),
  \1272(1898)  = \1086(1554)  & \1225(1819) ,
  \4955(1366)  = ~\4951(1200) ,
  \1002(1920)  = \3533(1846) ,
  \820(1283)  = \[38] ,
  \4376(2264)  = ~\4374(2211)  | ~\4371(1561) ,
  \4477(1825)  = \1482(1575)  | \1478(1731) ,
  \5233(1639)  = ~\5229(1467) ,
  \5222(1634)  = ~\5216(1460) ,
  \2330(2474)  = \2316(399)  & (\2281(210)  & \3653(2466) ),
  \2717(1191)  = \2702(910)  & \2682(1031) ,
  \1199(1865)  = ~\4195(1746)  | ~\4188(363) ,
  \1223(1899)  = ~\1222(1820)  | ~\1221(1722) ,
  \2556(580)  = ~\2553(342) ,
  \4258(1830)  = ~\4252(1737) ,
  \2642(555)  = ~\2639(316) ,
  \601(220)  = \[6] ,
  \2749(739)  = \2728(494)  & \281(108) ,
  \3956(1465)  = ~\3955(1242)  & ~\3954(1392) ,
  \5219(1458)  = ~\5151(1375)  | ~\5150(1373) ,
  \1174(1527)  = \1064(996)  & \1034(1429) ,
  \1444(1531)  = \1289(1428)  & (\1307(1427)  & \1422(1439) ),
  \1168(1542)  = \1046(1001)  & \1023(1432) ,
  \3938(1096)  = \3915(941) ,
  \3126(492)  = \3092(279)  & \338(124) ,
  \4691(1381)  = ~\4687(1235) ,
  \4578(2160)  = ~\4572(2115) ,
  \3286(991)  = ~\3285(876) ,
  \4927(1379)  = ~\4923(1228) ,
  \4409(1807)  = ~\1448(1698) ,
  \4719(1515)  = \1730(1422) ,
  \3348(1043)  = ~\3328(916) ,
  \2576(995)  = ~\2575(881) ,
  \5396(1110)  = ~\5375(776)  | ~\5374(949) ,
  \5216(1460)  = ~\5161(1385)  | ~\5160(1380) ,
  \4917(1383)  = ~\4913(1237) ,
  \5347(550)  = ~\5343(313) ,
  \2201(2453)  = ~\2198(2449) ,
  \4247(1553)  = \1089(1436) ,
  \3300(762)  = \3275(508)  & \2361(325) ,
  \4429(1560)  = \1422(1439) ,
  \2552(579)  = ~\2549(341) ,
  \2929(749)  = \2901(511)  & \3556(324) ,
  \4580(2214)  = ~\4578(2160)  | ~\4575(1742) ,
  \4887(1854)  = ~\4883(1760) ,
  \3509(1637)  = \3486(1464) ,
  \2666(458)  = \2639(316)  & (\400(137)  & \3553(198) ),
  \3437(1047)  = ~\3433(918) ,
  \3268(292)  = \308(116) ,
  \2672(453)  = \2647(312)  & (\411(138)  & \3553(198) ),
  \3283(432)  = \3268(292)  & (\479(144)  & \2405(329) ),
  \761(643)  = \2442(195)  & (\2418(193)  & \70(24) ),
  \705(964)  = \2869(677)  | (\2868(681)  | (\2867(962)  | \2866(958) )),
  \4365(1810)  = ~\4361(1703) ,
  \3963(2107)  = ~\5420(2058)  | ~\5417(1877) ,
  \673(1276)  = \[40] ,
  \2356(803)  = \2304(208)  & (\2293(401)  & \149(68) ),
  \1216(1999)  = ~\1215(1948) ,
  \5226(1468)  = ~\5205(1394)  | ~\5204(1393) ,
  \1659(2476)  = \1645(403)  & (\1609(214)  & \3653(2466) ),
  \1251(1903)  = ~\4274(1838)  | ~\4271(1570) ,
  \3428(1036)  = ~\3424(913) ,
  \3979(374)  = ~\3972(184) ,
  \1442(1535)  = \1318(997)  & \1289(1428) ,
  \1241(1907)  = ~\4258(1830)  | ~\4255(1589) ,
  \4954(2204)  = ~\4948(2149) ,
  \3112(495)  = ~\3105(278) ,
  \5059(1496)  = \2009(1416) ,
  \3431(720)  = ~\5096(491)  | ~\5093(268) ,
  \4791(1049)  = \3143(919) ,
  \1231(1897)  = ~\1225(1819) ,
  \3260(295)  = \302(114) ,
  \3905(744)  = ~\5347(550)  | ~\5340(318) ,
  \4472(1836)  = ~\4470(1193)  | ~\4467(1735) ,
  \5181(1111)  = \2802(950) ,
  \1210(1890)  = ~\4218(1804)  | ~\4215(1541) ,
  \5312(1145)  = \3297(877)  & \3286(991) ,
  \3264(291)  = \308(116) ,
  \3065(708)  = \3047(547)  & (\2370(326)  & \411(138) ),
  \2150(1616)  = \2089(1039)  & (\2042(1408)  & \2067(1403) ),
  \2595(387)  = \2541(346)  & \3547(201) ,
  \1173(1523)  = \1034(1429)  & (\1052(1426)  & \1080(1438) ),
  \4202(1814)  = ~\4196(1707) ,
  \3061(709)  = \3039(552)  & (\2370(326)  & \400(137) ),
  \1524(2454)  = ~\1521(2450) ,
  \1742(992)  = \479(144)  & \3161(926) ,
  \2113(1632)  = \1958(1074)  & (\1966(1067)  & (\1984(1423)  & \2099(1419) )),
  \2304(208)  = \1694(160) ,
  \2065(1124)  = ~\4802(411)  | ~\4799(1045) ,
  \4727(1514)  = \1730(1422) ,
  \3500(1755)  = ~\3497(1626) ,
  \1947(1941)  = \1909(1876)  & \1901(1882) ,
  \3531(1757)  = ~\5242(1628)  | ~\5239(1374) ,
  \[10]  = ~\338(124) ,
  \1483(1895)  = \1453(1718)  & \1462(1817) ,
  \3267(516)  = ~\3264(291) ,
  \[11]  = ~\358(128) ,
  \1926(1937)  = ~\1925(1780)  | ~\1924(1872) ,
  \2992(969)  = ~\2991(857) ,
  \2355(2091)  = \2316(399)  & (\2281(210)  & \3793(2065) ),
  \3765(371)  = ~\3757(181) ,
  \4274(1838)  = ~\4268(1747) ,
  \[12]  = \145(66)  & \141(65) ,
  \3047(547)  = ~\3044(310) ,
  \3934(1095)  = \3915(941) ,
  \1171(1526)  = \1064(996)  & \1034(1429) ,
  \1604(611)  = \1552(213)  & (\1528(215)  & \161(72) ),
  \[13]  = ~\245(98) ,
  \1004(1977)  = \3968(1930) ,
  \[14]  = ~\552(152) ,
  \5363(576)  = ~\5359(338) ,
  \3129(727)  = \3112(495)  & \316(118) ,
  \3512(1768)  = ~\3509(1637) ,
  \5236(1457)  = ~\3515(1372)  | ~\3518(1371) ,
  \2973(423)  = \2952(283)  & (\503(146)  & \3553(198) ),
  \1898(1946)  = ~\1897(1883) ,
  \[15]  = ~\562(155) ,
  \3967(1769)  = ~\5429(1642)  | ~\5422(1638) ,
  \3043(546)  = ~\3040(309) ,
  \5252(1976)  = ~\3527(1932)  | ~\3530(1929) ,
  \[16]  = ~\559(154) ,
  \3263(523)  = ~\3260(295) ,
  \5425(1470)  = ~\5405(1264)  | ~\5404(1397) ,
  \[17]  = ~\633(365) ,
  \3326(475)  = \3302(261)  & \2405(329) ,
  \5373(588)  = ~\5369(348) ,
  \[18]  = \814(203)  & \136(62) ,
  \1931(1914)  = ~\1930(1840)  | ~\1929(1751) ,
  \4172(1087)  = \2772(937) ,
  \[19]  = ~\844(657) ,
  \3396(892)  = \3395(705)  | \3394(449) ,
  \3493(503)  = \3440(284) ,
  \4491(1833)  = ~\4487(1743) ,
  \581(2045)  = ~\1954(1997) ,
  \5335(303)  = \289(110) ,
  \3397(1012)  = ~\3396(892) ,
  \4210(1812)  = ~\4204(1706) ,
  \4218(1804)  = ~\4212(1694) ,
  \5009(1664)  = ~\2153(1618)  & (~\2152(1479)  & ~\2059(975) ),
  \1916(1940)  = ~\1915(1790)  | ~\1914(1875) ,
  \3734(629)  = \3717(169)  & (\3728(196)  & \123(53) ),
  \1440(1534)  = \1318(997)  & (\1278(1433)  & \1289(1428) ),
  \611(275)  = \[10] ,
  \2151(1622)  = \2067(1403)  & (\2042(1408)  & \2106(1040) ),
  \2343(2093)  = \2316(399)  & (\2281(210)  & \3791(2067) ),
  \721(646)  = \2442(195)  & (\2418(193)  & \61(21) ),
  \3514(1057)  = \3489(504)  & (\3424(913)  & \3433(918) ),
  \4366(2110)  = ~\4364(2053)  | ~\4361(1703) ,
  \3382(333)  = \234(95) ,
  \3745(376)  = ~\3737(186) ,
  \[20]  = ~\846(254) ,
  \4471(1828)  = ~\4467(1735) ,
  \2121(1633)  = \1966(1067)  & (\1984(1423)  & \2099(1419) ),
  \1481(1528)  = \1307(1427)  & \1422(1439) ,
  \1208(1950)  = ~\1207(1811)  | ~\1206(1892) ,
  \5351(319)  = \257(102) ,
  \4255(1589)  = \1100(1448) ,
  \4690(1852)  = ~\4684(1759) ,
  \2898(288)  = \316(118) ,
  \2252(2094)  = \2238(400)  & (\2203(211)  & \4024(2068) ),
  \1238(1953)  = ~\1237(1818)  | ~\1236(1896) ,
  \3960(2108)  = ~\5412(2057)  | ~\5409(1998) ,
  \1892(1848)  = ~\4715(1376)  | ~\4708(1684) ,
  \2968(266)  = \351(127) ,
  \5029(1668)  = ~\2148(1615)  & (~\2147(1476)  & (~\2146(1409)  & ~\2036(864) )),
  \2939(1144)  = \2925(875)  & \2912(990) ,
  \[26]  = ~\3175(221) ,
  \1930(1840)  = ~\4763(1659)  | ~\4756(1363) ,
  \[27]  = ~\140(64)  | ~\2822(361) ,
  \4605(1549)  = \1332(1435) ,
  \[28]  = ~\2822(361) ,
  \2964(267)  = \351(127) ,
  \1657(2475)  = \1645(403)  & (\1621(405)  & \3654(2468) ),
  \4820(1879)  = ~\4818(1139)  | ~\4815(1794) ,
  \2020(1130)  = ~\4787(1052)  | ~\4780(230) ,
  \3329(702)  = \3310(595)  & (\446(141)  & \2405(329) ),
  \5097(484)  = ~\5093(268) ,
  \3086(899)  = \411(138)  | (\3085(752)  | \3083(545) ),
  \144(354)  = \141(65) ,
  \3553(198)  = ~\3552(168) ,
  \2927(510)  = \2898(288)  & \3554(331) ,
  \3505(1636)  = \3486(1464) ,
  \2382(327)  = \251(100) ,
  \3929(1786)  = ~\3926(1667) ,
  \1248(1959)  = ~\1247(1822)  | ~\1246(1906) ,
  \3001(395)  = \2956(272)  & \3547(201) ,
  \5386(1461)  = ~\5331(1387)  | ~\5330(1231) ,
  \857(849)  = \2500(189)  & (\2488(381)  & \11(2) ),
  \2260(603)  = \2226(209)  & (\2203(211)  & \173(76) ),
  \1521(2450)  = ~\1520(2448)  | ~\1519(2445) ,
  \4226(1802)  = ~\4220(1693) ,
  \4346(468)  = ~\4340(256) ,
  \2347(2088)  = \2316(399)  & (\2293(401)  & \3850(2069) ),
  \3056(462)  = \3028(321)  & (\389(136)  & \2393(328) ),
  \5005(1491)  = ~\5001(1413) ,
  \5243(1459)  = ~\5239(1374) ,
  \4936(1873)  = ~\4934(1784)  | ~\4931(1842) ,
  \5403(1103)  = ~\5399(946) ,
  \4019(2137)  = \3998(367)  & (\3972(184)  & \1263(2111) ),
  \2250(2090)  = \2238(400)  & (\2215(402)  & \4082(2071) ),
  \[34]  = ~\4094(527) ,
  \[35]  = ~\635(1114) ,
  \4263(1586)  = \1116(1446) ,
  \2130(1753)  = ~\2128(1619) ,
  \3869(1447)  = ~\5274(1334)  | ~\5271(1187) ,
  \[36]  = ~\703(1115) ,
  \2119(1153)  = \1995(993)  & \1966(1067) ,
  \[37]  = ~\716(1116) ,
  \2866(958)  = \2857(844)  & (\2838(398)  & \79(27) ),
  \[38]  = ~\819(1117) ,
  \4180(1083)  = \2767(936) ,
  \1580(605)  = \1552(213)  & (\1528(215)  & \170(75) ),
  \[39]  = \2827(620)  & \637(965) ,
  \3897(935)  = ~\3896(740)  | ~\3895(738) ,
  \4423(1809)  = ~\4419(1702) ,
  \2912(990)  = ~\2911(874) ,
  \3287(427)  = \3276(285)  & (\490(145)  & \2405(329) ),
  \3338(1003)  = \3337(886)  | \3336(701) ,
  \3892(1490)  = ~\3891(1305)  | ~\3890(1411) ,
  \3918(1715)  = \3871(1548) ,
  \847(465)  = \[20] ,
  \5359(338)  = \226(93) ,
  \3501(1625)  = \3463(1456) ,
  \5085(258)  = \369(131) ,
  \3532(1627)  = ~\5243(1459)  | ~\5236(1457) ,
  \1888(1924)  = ~\4706(1798)  | ~\4703(1225) ,
  \2040(1129)  = ~\4794(416)  | ~\4791(1049) ,
  \711(630)  = \3684(188)  & (\3660(190)  & \106(40) ),
  \4845(1516)  = \1984(1423) ,
  \3066(898)  = \3065(708)  | \3064(454) ,
  \3059(1027)  = ~\3058(906) ,
  \4581(2161)  = ~\4579(1832)  | ~\4572(2115) ,
  \1205(1951)  = ~\1204(1813)  | ~\1203(1891) ,
  \4123(443)  = ~\4119(242) ,
  \801(642)  = \2500(189)  & (\2476(191)  & \70(24) ),
  \[40]  = \2827(620)  & \671(966) ,
  \2271(790)  = \2226(209)  & (\2215(402)  & \194(83) ),
  \5294(1699)  = ~\5292(1543)  | ~\5289(1158) ,
  \3362(344)  = \218(91) ,
  \3366(343)  = \218(91) ,
  \[41]  = \2827(620)  & \705(964) ,
  \3352(1042)  = ~\3335(915) ,
  \[42]  = \2827(620)  & \713(967) ,
  \5369(348)  = \210(89) ,
  \2254(606)  = \2226(209)  & (\2203(211)  & \170(75) ),
  \[43]  = \597(1202)  & (\596(1412)  & \595(1463) ),
  \1213(1889)  = ~\4226(1802)  | ~\4223(1540) ,
  \[44]  = \609(1430)  & (\608(1440)  & \607(1425) ),
  \1266(1954)  = \1231(1897)  & \1223(1899) ,
  \791(658)  = \2500(189)  & (\2476(191)  & \20(5) ),
  \[45]  = \1451(1551)  & \1437(1530) ,
  \4643(430)  = ~\4639(235) ,
  \4484(2114)  = ~\4483(2010)  | ~\4482(2055) ,
  \3347(1002)  = \446(141)  | (\3346(943)  | \3345(769) ),
  \4250(1831)  = ~\4244(1739) ,
  \[46]  = \1857(1608)  & \1843(1630) ,
  \815(627)  = \[18] ,
  \1921(1939)  = ~\1920(1789)  | ~\1919(1874) ,
  \4077(2135)  = \4056(366)  & (\4030(183)  & \1944(2104) ),
  \3392(879)  = \3391(697)  | \3390(435) ,
  \[47]  = \2128(1619)  & \2113(1632) ,
  \1243(1961)  = ~\1242(1829)  | ~\1241(1907) ,
  \[48]  = \1179(1552)  & \1166(1522) ,
  \588(1696)  = \[45] ,
  \3882(1405)  = ~\5303(1297)  | ~\5296(1127) ,
  \2986(972)  = ~\2985(858) ,
  \4832(2166)  = ~\4831(2061)  | ~\4830(2119) ,
  \3440(284)  = ~\324(120) ,
  \810(356)  = \[12] ,
  \4175(248)  = \411(138) ,
  \1662(2477)  = \1661(601)  | (\1660(799)  | (\1659(2476)  | \1657(2475) )),
  \1952(1945)  = \1909(1876)  & \1758(1420) ,
  \5063(1671)  = ~\5059(1496) ,
  \2281(210)  = \1691(159) ,
  \1253(1960)  = ~\1252(1824)  | ~\1251(1903) ,
  \2353(2089)  = \2316(399)  & (\2293(401)  & \3851(2063) ),
  \2913(428)  = \2902(287)  & (\490(145)  & \2393(328) ),
  \1847(1509)  = \1712(1065)  & (\1749(988)  & (\1704(1073)  & \1730(1422) )),
  \5126(912)  = \3119(470)  | \3118(715) ,
  \2976(866)  = \2975(691)  | \2973(423) ,
  \[51]  = \590(1806)  | \589(1711) ,
  \4667(415)  = ~\4663(228) ,
  \[52]  = \617(1849)  | \616(1763) ,
  \3167(931)  = \3136(529)  | \3135(736) ,
  \[53]  = \620(1800)  | \619(1710) ,
  \2574(698)  = \2548(584)  & (\3551(199)  & \468(143) ),
  \3247(417)  = \514(147)  | \3555(332) ,
  \[54]  = \628(1853)  | \627(1764) ,
  \3288(693)  = \3279(506)  & (\2382(327)  & \490(145) ),
  \2116(1152)  = \1995(993)  & (\1958(1074)  & \1966(1067) ),
  \[55]  = ~\3848(1864) ,
  \1701(355)  = \141(65) ,
  \[56]  = ~\3849(2024) ,
  \4322(459)  = ~\4316(250) ,
  \4424(2109)  = ~\4422(2054)  | ~\4419(1702) ,
  \3881(1402)  = ~\5302(1302)  | ~\5299(1122) ,
  \[57]  = ~\3790(2025) ,
  \4110(298)  = \299(113) ,
  \2980(690)  = ~\2979(420) ,
  \[58]  = ~\1936(2105) ,
  \4151(245)  = \435(140) ,
  \1855(1507)  = \1730(1422)  & \1758(1420) ,
  \[59]  = \721(646)  | (\720(848)  | (\719(2030)  | \718(1867) )),
  \1884(1928)  = ~\4698(1851)  | ~\4695(1236) ,
  \4716(989)  = ~\3155(924)  & ~\490(145) ,
  \4890(2165)  = ~\4889(2060)  | ~\4888(2118) ,
  \781(652)  = \3684(188)  & (\3660(190)  & \40(14) ),
  \3933(1785)  = ~\3930(1666) ,
  \2293(401)  = ~\2281(210) ,
  \2948(282)  = \324(120) ,
  \3757(181)  = \4092(176) ,
  \2960(273)  = \341(125) ,
  \4812(986)  = ~\3155(924)  & ~\490(145) ,
  \4351(1805)  = \1481(1528)  | \1448(1698) ,
  \[60]  = ~\4082(2071) ,
  \597(1202)  = ~\3348(1043) ,
  \4271(1570)  = \1134(1442) ,
  \4671(227)  = \534(149) ,
  \[61]  = ~\3851(2063) ,
  \5073(1662)  = ~\5069(1487) ,
  \4371(1561)  = \1422(1439) ,
  \[62]  = ~\3850(2069) ,
  \3468(1469)  = ~\3467(1396)  | ~\3466(1395) ,
  \4783(921)  = \3147(723) ,
  \[63]  = \858(647)  | (\857(849)  | (\856(2029)  | \855(1866) )),
  \5053(1656)  = ~\5049(1475) ,
  \3477(1471)  = ~\3476(1399)  | ~\3475(1398) ,
  \3284(696)  = \3271(517)  & (\2382(327)  & \479(144) ),
  \[64]  = ~\4024(2068) ,
  \1486(1952)  = ~\1483(1895) ,
  \3067(1019)  = ~\3066(898) ,
  \[65]  = ~\3793(2065) ,
  \[66]  = ~\3792(2066) ,
  \[67]  = ~\3791(2067) ,
  \5173(1104)  = \2794(947) ,
  \2605(389)  = \2557(337)  & \3547(201) ,
  \3416(893)  = \422(139)  | (\3415(756)  | \3413(567) ),
  \2942(1137)  = \2930(872)  & \2916(985) ,
  \4083(2130)  = \4072(821)  | (\4071(2026)  | \4070(1285) ),
  \3737(186)  = \4091(175) ,
  \4025(2129)  = \4014(820)  | (\4013(2027)  | \4012(1288) ),
  \3343(1004)  = \446(141)  | (\3342(942)  | \3341(768) ),
  \4655(231)  = \514(147) ,
  \5394(1676)  = ~\5392(1635)  | ~\5389(1499) ,
  \2331(798)  = \2304(208)  & (\2293(401)  & \176(77) ),
  \751(659)  = \2442(195)  & (\2418(193)  & \20(5) ),
  \[70]  = \574(2158)  & (\573(2157)  & (\572(2113)  & (\571(2052)  & (\570(2001)  & (\569(2012)  & (\568(2008)  & (\567(2009)  & \566(1979) ))))))),
  \[71]  = \584(2151)  & (\583(2150)  & (\582(2106)  & (\581(2045)  & (\580(1991)  & (\579(1990)  & (\578(1988)  & (\577(1967)  & \576(1776) ))))))),
  \5162(1100)  = \2788(945) ,
  \3036(314)  = \265(104) ,
  \[72]  = \1606(623)  & \659(2121) ,
  \[73]  = \2279(625)  & \691(2122) ,
  \3032(315)  = \265(104) ,
  \[74]  = \746(654)  | (\745(841)  | (\744(2081)  | \743(2082) )),
  \5322(932)  = \3293(761)  | \3292(531) ,
  \2734(276)  = \335(123) ,
  \1467(1596)  = \1344(1449)  & (\1412(1033)  & (\1365(1445)  & \1390(1443) )),
  \1457(1597)  = \1344(1449)  & (\1412(1033)  & (\1332(1435)  & (\1365(1445)  & \1390(1443) ))),
  \3208(281)  = \324(120) ,
  \1764(1508)  = ~\1758(1420) ,
  \[75]  = \751(659)  | (\750(831)  | (\749(2083)  | \748(2086) )),
  \1271(1955)  = \1231(1897)  & \1080(1438) ,
  \3175(221)  = \549(151) ,
  \2166(2399)  = ~\2165(2378)  | ~\2164(2388) ,
  \4026(2185)  = \4017(836)  | (\4016(2073)  | \4015(1289) ),
  \[76]  = \756(660)  | (\755(832)  | (\754(2084)  | \753(2087) )),
  \3556(324)  = \254(101) ,
  \[77]  = \761(643)  | (\760(835)  | (\759(2085)  | \758(2031) )),
  \3204(280)  = \324(120) ,
  \[78]  = \786(653)  | (\785(840)  | (\784(2077)  | \783(2074) )),
  \4340(256)  = \374(134) ,
  \5393(1677)  = ~\5389(1499) ,
  \[79]  = \791(658)  | (\790(830)  | (\789(2078)  | \788(2075) )),
  \3401(1008)  = ~\3400(889) ,
  \3922(1714)  = \3871(1548) ,
  \4119(242)  = \446(141) ,
  \5268(1166)  = \3421(888)  & \3401(1008) ,
  \1178(1559)  = \1071(1014)  & \1052(1426) ,
  \2036(864)  = \3147(723)  & \514(147) ,
  \4022(2136)  = \3998(367)  & (\3972(184)  & \1258(2112) ),
  \1881(1927)  = ~\4690(1852)  | ~\4687(1235) ,
  \1469(1583)  = \1382(1024)  & \1344(1449) ,
  \3777(2209)  = ~\3962(2154) ,
  \4631(236)  = \479(144) ,
  \1179(1552)  = \1134(1442)  & (\1089(1436)  & (\1116(1446)  & (\1152(1452)  & \1100(1448) ))),
  \5170(1107)  = \2798(948) ,
  \2767(936)  = \2750(537)  | \2749(739) ,
  \1256(2049)  = \1231(1897)  & \1209(2000) ,
  \3224(264)  = \351(127) ,
  \2802(950)  = \2766(593)  | \2765(783) ,
  \4559(1827)  = ~\4555(1734) ,
  \5289(1158)  = \3406(883)  & \3389(998) ,
  \1220(1956)  = ~\1219(1900) ,
  \[80]  = \796(661)  | (\795(833)  | (\794(2079)  | \793(2076) )),
  \1189(1567)  = \1100(1448)  & (\1145(1020)  & \1116(1446) ),
  \3220(265)  = \351(127) ,
  \741(651)  = \3582(194)  & (\3558(192)  & \40(14) ),
  \[81]  = \801(642)  | (\800(834)  | (\799(2080)  | \798(2028) )),
  \3331(1005)  = \3330(887)  | \3329(702) ,
  \1288(1328)  = ~\4291(1269)  | ~\4284(240) ,
  \1891(1923)  = ~\4714(1797)  | ~\4711(1224) ,
  \3486(1464)  = ~\3485(1388)  | ~\3484(1241) ,
  \5206(929)  = ~\5117(735)  | ~\5116(731) ,
  \[82]  = \1526(622)  & \640(2170) ,
  \4639(235)  = \490(145) ,
  \[83]  = \1606(623)  & \662(2173) ,
  \3085(752)  = \3043(546)  & \3556(324) ,
  \5383(1689)  = ~\5379(1518) ,
  \2122(1151)  = \1995(993)  & \1966(1067) ,
  \[84]  = \1606(623)  & \665(2174) ,
  \2916(985)  = ~\2915(873) ,
  \[85]  = \1606(623)  & \668(2177) ,
  \4135(238)  = \468(143) ,
  \993(850)  = \1688(663) ,
  \[86]  = \2202(626)  & \674(2171) ,
  \921(664)  = \2826(364) ,
  \[87]  = \2279(625)  & \694(2172) ,
  \3075(750)  = \3027(561)  & \3556(324) ,
  \1591(789)  = \1552(213)  & (\1540(406)  & \197(84) ),
  \1389(1347)  = ~\4331(1248)  | ~\4324(249) ,
  \[88]  = \2279(625)  & \697(2175) ,
  \3071(1030)  = ~\3070(909) ,
  \3063(1022)  = ~\3062(901) ,
  \[89]  = \2279(625)  & \700(2176) ,
  \1181(1590)  = \1111(1028)  & \1089(1436) ,
  \3181(205)  = ~\2358(162) ,
  \731(650)  = \3582(194)  & (\3558(192)  & \49(17) ),
  \1086(1554)  = ~\1080(1438) ,
  \3314(260)  = \361(129) ,
  \2882(302)  = \293(112) ,
  \3835(2206)  = ~\3965(2153) ,
  \3137(914)  = \3121(472)  | \3120(717) ,
  \5046(2325)  = ~\5045(2289)  | ~\5044(2312) ,
  \4194(662)  = ~\4188(363) ,
  \1176(1558)  = \1071(1014)  & \1052(1426) ,
  \1845(1226)  = \1724(1066)  & \1704(1073) ,
  \3256(301)  = \293(112) ,
  \4080(2134)  = \4056(366)  & (\4030(183)  & \1936(2105) ),
  \3445(1455)  = ~\3444(1368)  | ~\3443(1369) ,
  \3052(304)  = \281(108) ,
  \[90]  = \817(2230)  & \816(628) ,
  \3896(740)  = ~\5339(536)  | ~\5332(308) ,
  \1688(663)  = \2826(364) ,
  \1806(974)  = \523(148)  & \3143(919) ,
  \[91]  = \812(2205)  | \811(2219) ,
  \4308(253)  = \389(136) ,
  \4084(2180)  = \4075(817)  | (\4074(2072)  | \4073(1286) ),
  \4876(1315)  = ~\4870(1140) ,
  \3143(919)  = \3125(485)  | \3124(721) ,
  \[92]  = ~\4086(2231) ,
  \1609(214)  = \1689(157) ,
  \[93]  = ~\4085(2232) ,
  \5054(2338)  = ~\5052(2336)  | ~\5049(1475) ,
  \1258(2112)  = \1257(2004)  | \1256(2049) ,
  \2990(686)  = \2971(482)  & (\3551(199)  & \534(149) ),
  \[94]  = ~\4084(2180) ,
  \1579(787)  = \1552(213)  & (\1540(406)  & \200(85) ),
  \[95]  = ~\4083(2130) ,
  \632(1692)  = \[48] ,
  \1468(1572)  = \1390(1443)  & (\1344(1449)  & (\1365(1445)  & \1430(1451) )),
  \[96]  = \245(98)  & (\853(2202)  & \852(255) ),
  \2067(1403)  = ~\2066(1299)  | ~\2065(1124) ,
  \3861(1444)  = ~\5267(1345)  | ~\5260(1182) ,
  \[97]  = ~\4028(2234) ,
  \5055(2327)  = ~\5053(1656)  | ~\5046(2325) ,
  \[98]  = ~\4027(2235) ,
  \2155(1657)  = \2154(1617)  | \2081(970) ,
  \1678(2099)  = \1645(403)  & (\1609(214)  & \3792(2066) ),
  \2914(694)  = \2905(509)  & (\2370(326)  & \490(145) ),
  \4096(2167)  = ~\1936(2105)  | ~\4113(1859) ,
  \[99]  = ~\4026(2185) ,
  \1175(1556)  = \1034(1429)  & (\1052(1426)  & \1071(1014) ),
  \3433(918)  = ~\3432(722)  | ~\3431(720) ,
  \3281(767)  = \3263(523)  & \2382(327) ,
  \1585(785)  = \1552(213)  & (\1540(406)  & \203(86) ),
  \2259(784)  = \2226(209)  & (\2215(402)  & \203(86) ),
  \4948(2149)  = ~\4947(2038)  | ~\4946(2103) ,
  \2984(687)  = \2963(490)  & (\3551(199)  & \523(148) ),
  \3860(1441)  = ~\5266(1348)  | ~\5263(1179) ,
  \2910(695)  = \2897(520)  & (\2370(326)  & \479(144) ),
  \4579(1832)  = ~\4575(1742) ,
  \1473(1599)  = \1412(1033)  & (\1365(1445)  & \1390(1443) ),
  \1466(1577)  = \1344(1449)  & (\1404(1021)  & \1365(1445) ),
  \1209(2000)  = ~\1208(1950) ,
  \3199(639)  = \3181(205)  & \88(34) ,
  \1454(1593)  = \1359(1029)  & \1332(1435) ,
  \1576(2097)  = \1564(404)  & (\1540(406)  & \4082(2071) ),
  \1456(1578)  = \1344(1449)  & (\1404(1021)  & (\1332(1435)  & \1365(1445) )),
  \2765(783)  = \2741(493)  & \206(87) ,
  \2265(788)  = \2226(209)  & (\2215(402)  & \197(84) ),
  \3901(1081)  = ~\3897(935) ,
  \1447(1565)  = \1324(1017)  & \1307(1427) ,
  \2160(1916)  = \2130(1753)  & \2139(1792) ,
  \3463(1456)  = ~\3462(1210)  | ~\3461(1370) ,
  \2687(905)  = \389(136)  | (\2686(670)  | \2684(390) ),
  \3377(578)  = ~\3374(340) ,
  \5052(2336)  = ~\5046(2325) ,
  \3406(883)  = \457(142)  | (\3405(754)  | \3403(565) ),
  \2279(625)  = \1698(358) ,
  \2933(933)  = \2920(747)  | \2918(533) ,
  \3454(1453)  = ~\3453(1361)  | ~\3452(1196) ,
  \1465(1584)  = \1382(1024)  & \1344(1449) ,
  \1455(1585)  = \1382(1024)  & (\1332(1435)  & \1344(1449) ),
  \2880(684)  = \2847(656)  & \2838(398) ,
  \5279(1170)  = \3416(893)  & \3397(1012) ,
  \3496(725)  = ~\3493(503) ,
  \4355(1886)  = ~\4351(1805) ,
  \809(655)  = \[28] ,
  \4565(1826)  = ~\1478(1731) ,
  \1475(1579)  = \1404(1021)  & \1365(1445) ,
  \2179(207)  = ~\2174(161) ,
  \5276(1154)  = \3411(878)  & \3393(994) ,
  \4347(1246)  = ~\4343(1084) ,
  \1188(1587)  = \1128(1025)  & \1100(1448) ,
  \3373(577)  = ~\3370(339) ,
  \5039(1199)  = \2106(1040) ,
  \3236(860)  = \3235(688)  | \3234(414) ,
  \3870(1434)  = ~\5275(1353)  | ~\5268(1166) ,
  \1446(1564)  = \1289(1428)  & (\1324(1017)  & \1307(1427) ),
  \3866(1726)  = ~\3862(1566) ,
  \4103(1386)  = \3170(1076)  & \4099(1240) ,
  \3325(781)  = ~\3322(597) ,
  \2761(774)  = \2741(493)  & \218(91) ,
  \5329(1232)  = ~\5325(1070) ,
  \3321(780)  = ~\3318(596) ,
  \1471(1598)  = \1344(1449)  & (\1412(1033)  & (\1365(1445)  & \1390(1443) )),
  \2868(681)  = \2847(656)  & \2838(398) ,
  \1516(2407)  = \1497(156)  & (\1486(1952)  & \1489(2393) ),
  \4178(1249)  = ~\4172(1087) ,
  \4931(1842)  = \2159(1621)  | \2155(1657) ,
  \2857(844)  = ~\2847(656) ,
  \2662(711)  = \2634(564)  & (\3551(199)  & \389(136) ),
  \2963(490)  = ~\2960(273) ,
  \5044(2312)  = ~\5042(2280)  | ~\5039(1199) ,
  \3549(200)  = ~\3548(166) ,
  \1509(2431)  = ~\4550(2425)  | ~\4547(1591) ,
  \2759(773)  = \2741(493)  & \226(93) ,
  \3309(778)  = ~\3306(594) ,
  \3910(1088)  = ~\3906(938) ,
  \5066(2383)  = ~\5065(2359)  | ~\5064(2370) ,
  \3492(726)  = ~\3489(504) ,
  \4413(1887)  = ~\4409(1807) ,
  \1676(2095)  = \1645(403)  & (\1621(405)  & \3850(2069) ),
  \1172(1557)  = \1034(1429)  & (\1071(1014)  & \1052(1426) ),
  \3783(809)  = \3757(181)  & (\3745(376)  & \126(54) ),
  \2135(1673)  = \2134(1614)  | (\2133(1478)  | (\2132(1489)  | (\2131(1493)  | \2018(982) ))),
  \4113(1859)  = \4112(1774)  | \4111(1765) ,
  \5258(2022)  = ~\5252(1976) ,
  \1515(2408)  = \1497(156)  & (\1483(1895)  & \1494(2394) ),
  \3088(539)  = \3048(305)  & \3554(331) ,
  \5149(1217)  = ~\5145(1058) ,
  \1899(1680)  = ~\4730(1317)  | ~\4727(1514) ,
  \1183(1568)  = \1100(1448)  & (\1145(1020)  & (\1089(1436)  & \1116(1446) )),
  \2663(904)  = \2662(711)  | \2660(461) ,
  \1267(2003)  = \1220(1956)  & \1225(1819) ,
  \1472(1580)  = \1404(1021)  & \1365(1445) ,
  \1257(2004)  = \1205(1951)  & \1225(1819) ,
  \5372(782)  = ~\5366(598) ,
  \4368(2156)  = ~\4367(2048)  | ~\4366(2110) ,
  \1474(1573)  = \1390(1443)  & (\1365(1445)  & \1430(1451) ),
  \4730(1317)  = ~\4724(1142) ,
  \1684(2098)  = \1645(403)  & (\1609(214)  & \3793(2065) ),
  \3345(769)  = \3318(596)  & \3555(332) ,
  \2142(1410)  = \2059(975)  & \2021(1306) ,
  \1507(2428)  = ~\4541(1741)  | ~\4534(2419) ,
  \1508(2435)  = ~\1507(2428)  | ~\1506(2432) ,
  \3341(768)  = \3306(594)  & \3555(332) ,
  \4099(1240)  = ~\3170(1076) ,
  \1514(2406)  = \1502(216)  & (\1458(1719)  & \1489(2393) ),
  \1263(2111)  = \1262(2002)  | \1261(2051) ,
  \1513(2405)  = \1502(216)  & (\1462(1817)  & \1494(2394) ),
  \5006(1198)  = \2089(1039) ,
  \2169(2389)  = ~\4926(2380)  | ~\4923(1228) ,
  \5101(289)  = \316(118) ,
  \887(528)  = \4110(298) ,
  \1078(1340)  = ~\4146(1263)  | ~\4143(246) ,
  \1519(2445)  = ~\4626(2421)  | ~\4623(2442) ,
  \1306(1325)  = ~\4299(1267)  | ~\4292(239) ,
  \1421(1342)  = ~\4339(1262)  | ~\4332(247) ,
  \1277(1333)  = ~\4283(1274)  | ~\4276(243) ,
  \4017(836)  = \3991(179)  & (\3979(374)  & \53(19) ),
  \1856(1513)  = \1749(988)  & \1730(1422) ,
  \5111(296)  = \302(114) ,
  \2042(1408)  = ~\2041(1304)  | ~\2040(1129) ,
  \3357(589)  = ~\3354(349) ,
  \5307(862)  = \3247(417)  & \3233(689) ,
  \1518(2436)  = \1508(2435)  & \1497(156) ,
  \5148(1221)  = ~\5142(1062) ,
  \3073(560)  = \3024(320)  & \3554(331) ,
  \1192(1569)  = \1116(1446)  & \1145(1020) ,
  \3528(1861)  = \3512(1768)  & (\3481(1643)  & \3468(1469) ),
  \1443(1562)  = \1289(1428)  & (\1324(1017)  & \1307(1427) ),
  \3405(754)  = \3357(589)  & \3556(324) ,
  \3393(994)  = ~\3392(879) ,
  \881(370)  = \3757(181)  & \3737(186) ,
  \4888(2118)  = ~\4886(2044)  | ~\4883(1760) ,
  \4186(1245)  = ~\4180(1083) ,
  \4487(1743)  = \1468(1572)  | (\1467(1596)  | (\1466(1577)  | (\1465(1584)  | \1359(1029) ))),
  \3890(1411)  = ~\5310(1309)  | ~\5307(862) ,
  \3008(676)  = \2967(483)  & \3549(200) ,
  \3696(378)  = ~\3684(188) ,
  \1482(1575)  = \1390(1443)  & \1430(1451) ,
  \3415(756)  = \3373(577)  & \3556(324) ,
  \1331(1336)  = ~\4307(1260)  | ~\4300(244) ,
  \2125(1688)  = \2124(1506)  | \1995(993) ,
  \4094(527)  = \4110(298) ,
  \4275(1728)  = ~\4271(1570) ,
  \1170(1555)  = \1034(1429)  & (\1071(1014)  & (\1023(1432)  & \1052(1426) )),
  \1682(2096)  = \1645(403)  & (\1621(405)  & \3851(2063) ),
  \2345(613)  = \2304(208)  & (\2281(210)  & \158(71) ),
  \5159(1230)  = ~\5155(1069) ,
  \4268(1747)  = \1197(1650)  | \1160(1034) ,
  \3243(498)  = \3204(280)  & \3555(332) ,
  \3848(1864)  = \3838(804)  | (\3837(1653)  | \3836(1120) ),
  \602(222)  = \[7] ,
  \1506(2432)  = ~\4540(2426)  | ~\4537(1592) ,
  \2351(616)  = \2304(208)  & (\2281(210)  & \152(69) ),
  \5158(1239)  = ~\5152(1075) ,
  \5064(2370)  = ~\5062(2358)  | ~\5059(1496) ,
  \1087(1337)  = ~\4154(1259)  | ~\4151(245) ,
  \1470(1576)  = \1344(1449)  & (\1404(1021)  & \1365(1445) ),
  \1854(1512)  = \1749(988)  & \1730(1422) ,
  \5263(1179)  = \3086(899)  & \3067(1019) ,
  \2825(204)  = ~\2824(163) ,
  \598(1623)  = \[43] ,
  \1517(2440)  = \1502(216)  & \1512(2438) ,
  \3390(435)  = \3366(343)  & (\468(143)  & \2393(328) ),
  \4023(818)  = \3991(179)  & (\3979(374)  & \115(45) ),
  \4746(1782)  = ~\4740(1661) ,
  \4259(1738)  = ~\4255(1589) ,
  \4467(1735)  = \1474(1573)  | (\1473(1599)  | (\1472(1580)  | \1382(1024) )),
  \2165(2378)  = ~\4869(1378)  | ~\4862(2368) ,
  \766(644)  = \2442(195)  & (\2418(193)  & \64(22) ),
  \1441(1563)  = \1289(1428)  & (\1324(1017)  & (\1278(1433)  & \1307(1427) )),
  \5271(1187)  = \3076(907)  & \3059(1027) ,
  \4331(1248)  = ~\4327(1086) ,
  \4290(441)  = ~\4284(240) ,
  \4426(2155)  = ~\4425(2047)  | ~\4424(2109) ,
  \4946(2103)  = ~\4944(2037)  | ~\4941(1669) ,
  \1853(1510)  = \1712(1065)  & (\1730(1422)  & \1749(988) ),
  \1895(1681)  = ~\4722(1143)  | ~\4719(1515) ,
  \5056(2350)  = ~\5055(2327)  | ~\5054(2338) ,
  \1182(1588)  = \1128(1025)  & (\1089(1436)  & \1100(1448) ),
  \3525(1863)  = \3508(1766)  & (\3477(1471)  & \3472(1641) ),
  \5214(1220)  = ~\5212(1071)  | ~\5209(925) ,
  \1273(2005)  = \1272(1898)  | \1271(1955) ,
  \5065(2359)  = ~\5063(1671)  | ~\5056(2350) ,
  \776(632)  = \3684(188)  & (\3660(190)  & \103(39) ),
  \4572(2115)  = ~\4571(2011)  | ~\4570(2056) ,
  \3523(1749)  = \3501(1625)  & (\3449(1624)  & \3458(1607) ),
  \3432(722)  = ~\5097(484)  | ~\5090(274) ,
  \3280(522)  = \3260(295)  & \2405(329) ,
  \4560(1837)  = ~\4558(1359)  | ~\4555(1734) ,
  \3398(445)  = \3382(333)  & (\435(140)  & \2393(328) ),
  \3847(805)  = \3815(180)  & (\3803(375)  & \130(58) ),
  \3018(1126)  = \3004(859)  & \2986(972) ,
  \2697(897)  = \411(138)  | (\2696(672)  | \2694(392) ),
  \2099(1419)  = ~\2098(1314)  | ~\2097(1138) ,
  \4187(469)  = ~\4183(257) ,
  \4419(1702)  = ~\1446(1564)  & (~\1445(1533)  & ~\1301(1000) ),
  \5413(2046)  = ~\5409(1998) ,
  \2586(704)  = \2564(573)  & (\3551(199)  & \435(140) ),
  \3122(719)  = \3099(496)  & \351(127) ,
  \3422(716)  = ~\5088(477)  | ~\5085(258) ,
  \2009(1416)  = ~\2008(1310)  | ~\2007(1134) ,
  \4684(1759)  = \1851(1631)  | (\1850(1511)  | (\1849(1148)  | \1724(1066) )),
  \1262(2002)  = \1212(1949)  & \1225(1819) ,
  \1949(2040)  = \1948(1993)  | \1947(1941) ,
  \4267(1736)  = ~\4263(1586) ,
  \852(255)  = \552(152)  & (\556(153)  & (\559(154)  & \386(135) )),
  \889(734)  = \4094(527) ,
  \4163(463)  = ~\4159(252) ,
  \3253(480)  = \3220(265)  & \3555(332) ,
  \3333(473)  = \3314(260)  & \2405(329) ,
  \5354(572)  = ~\5348(335) ,
  \5260(1182)  = \3081(900)  & \3063(1022) ,
  \4298(438)  = ~\4292(239) ,
  \3394(449)  = \3374(340)  & (\422(139)  & \2393(328) ),
  \2650(549)  = ~\2647(312) ,
  \5406(2013)  = ~\3944(1962)  | ~\3947(1963) ,
  \4493(2162)  = ~\4491(1833)  | ~\4484(2114) ,
  \4998(2416)  = ~\4997(2390)  | ~\4996(2409) ,
  \2164(2388)  = ~\4868(2381)  | ~\4865(1227) ,
  \1451(1551)  = \1332(1435)  & (\1344(1449)  & (\1365(1445)  & (\1390(1443)  & \1430(1451) ))),
  \1132(1346)  = ~\4178(1249)  | ~\4175(248) ,
  \2967(483)  = ~\2964(267) ,
  \3027(561)  = ~\3024(320) ,
  \4367(2048)  = ~\4365(1810)  | ~\4358(2006) ,
  \4754(1781)  = ~\4748(1658) ,
  \2658(541)  = ~\2655(306) ,
  \4825(1761)  = \2121(1633)  | (\2120(1503)  | (\2119(1153)  | \1978(1068) )),
  \2316(399)  = ~\2304(208) ,
  \4889(2060)  = ~\4887(1854)  | ~\4880(1996) ,
  \3207(499)  = ~\3204(280) ,
  \846(254)  = \556(153)  & \386(135) ,
  \4009(1287)  = \3998(367)  & (\3979(374)  & \2623(1167) ),
  \4395(1713)  = ~\4391(1547) ,
  \3672(380)  = ~\3660(190) ,
  \2587(891)  = \2586(704)  | \2584(446) ,
  \2988(410)  = \2968(266)  & (\534(149)  & \3553(198) ),
  \2654(542)  = ~\2651(307) ,
  \2393(328)  = \248(99) ,
  \1850(1511)  = \1712(1065)  & (\1749(988)  & \1730(1422) ),
  \3317(474)  = ~\3314(260) ,
  \2584(446)  = \2561(336)  & (\435(140)  & \3553(198) ),
  \790(830)  = \2500(189)  & (\2488(381)  & \76(26) ),
  \5062(2358)  = ~\5056(2350) ,
  \5215(1233)  = ~\5213(1061)  | ~\5206(929) ,
  \1511(2434)  = ~\1510(2427)  | ~\1509(2431) ,
  \3520(1748)  = \3497(1626)  & (\3445(1455)  & \3454(1453) ),
  \3336(701)  = \3322(597)  & (\446(141)  & \2405(329) ),
  \1863(1675)  = \1862(1610)  | (\1861(1482)  | (\1860(1486)  | (\1859(1495)  | \1775(983) ))),
  \3227(479)  = ~\3224(264) ,
  \4425(2047)  = ~\4423(1809)  | ~\4416(2007) ,
  \656(621)  = \[27] ,
  \4251(1720)  = ~\4247(1553) ,
  \4260(1727)  = \1196(1651)  | (\1195(1605)  | \1145(1020) ),
  \1512(2438)  = ~\1511(2434) ,
  \1477(1600)  = \1412(1033)  & \1390(1443) ,
  \5332(308)  = \281(108) ,
  \2750(537)  = \2721(277)  & \288(109) ,
  \4195(1746)  = ~\4191(1602) ,
  \4433(1724)  = ~\4429(1560) ,
  \4692(1758)  = ~\1853(1510)  & (~\1852(1149)  & ~\1724(1066) ),
  \3123(478)  = \3092(279)  & \358(128) ,
  \3012(1132)  = \2997(867)  & \2977(980) ,
  \5088(477)  = ~\5082(262) ,
  \3197(953)  = \3196(640)  | \3195(828) ,
  \4794(416)  = ~\4788(229) ,
  \1510(2427)  = ~\4551(1740)  | ~\4544(2418) ,
  \4676(360)  = \54(20) ,
  \5140(1211)  = ~\5134(1054) ,
  \3632(377)  = ~\3628(187) ,
  \4770(434)  = ~\4764(237) ,
  \612(263)  = \[11] ,
  \5330(1231)  = ~\5328(1077)  | ~\5325(1070) ,
  \732(2300)  = \[103] ,
  \2146(1409)  = \2059(975)  & \2021(1306) ,
  \688(2317)  = \[116] ,
  \3660(190)  = \4089(173) ,
  \4219(1705)  = ~\4215(1541) ,
  \5250(2016)  = ~\5244(1966) ,
  \2170(2379)  = ~\4927(1379)  | ~\4920(2367) ,
  \1778(1307)  = ~\1777(979)  | ~\1776(1131) ,
  \973(202)  = \3173(164) ,
  \3403(565)  = \3354(349)  & \3554(331) ,
  \3176(362)  = \27(10)  & \31(11) ,
  \770(838)  = \3684(188)  & (\3672(380)  & \46(16) ),
  \736(633)  = \3582(194)  & (\3558(192)  & \103(39) ),
  \4375(1725)  = ~\4371(1561) ,
  \3223(481)  = ~\3220(265) ,
  \5019(1779)  = ~\2155(1657) ,
  \4883(1760)  = ~\2123(1505)  & (~\2122(1151)  & ~\1978(1068) ),
  \1476(1601)  = \1412(1033)  & (\1365(1445)  & \1390(1443) ),
  \3006(396)  = \2964(267)  & \3547(201) ,
  \5414(2018)  = ~\3950(1970)  | ~\3953(1971) ,
  \3558(192)  = \4088(172) ,
  \3413(567)  = \3370(339)  & \3554(331) ,
  \726(631)  = \3582(194)  & (\3558(192)  & \106(40) ),
  \4405(1700)  = ~\4401(1537) ,
  \1021(1332)  = ~\4122(1273)  | ~\4119(242) ,
  \4067(1284)  = \4056(366)  & (\4037(373)  & \3012(1132) ),
  \2748(535)  = \2721(277)  & \292(111) ,
  \2867(962)  = \2857(844)  & (\2828(206)  & \23(6) ),
  \4778(425)  = ~\4772(232) ,
  \780(826)  = \3684(188)  & (\3672(380)  & \91(35) ),
  \3170(1076)  = \3167(931) ,
  \1934(2039)  = \1909(1876)  & \1887(2021) ,
  \4244(1739)  = \1191(1649)  | (\1190(1603)  | (\1189(1567)  | (\1188(1587)  | \1111(1028) ))),
  \4738(1791)  = ~\4732(1670) ,
  \4147(451)  = ~\4143(246) ,
  \806(645)  = \2500(189)  & (\2476(191)  & \64(22) ),
  \796(661)  = \2500(189)  & (\2476(191)  & \17(4) ),
  \3134(521)  = \3105(278)  & \307(115) ,
  \2822(361)  = \31(11)  & \27(10) ,
  \2997(867)  = \503(146)  | (\2996(674)  | \2994(394) ),
  \3684(188)  = \4090(174) ,
  \1777(979)  = ~\4659(422)  | ~\4652(920) ,
  \1268(2050)  = \1267(2003)  | \1266(1954) ,
  \4056(366)  = ~\4049(178) ,
  \4276(243)  = \446(141) ,
  \2826(364)  = \1(0) ,
  \2418(193)  = \4088(172) ,
  \5193(1244)  = ~\5189(1082) ,
  \4227(1704)  = ~\4223(1540) ,
  \3622(372)  = ~\3616(182) ,
  \4252(1737)  = \1194(1652)  | (\1193(1606)  | (\1192(1569)  | \1128(1025) )),
  \3021(1123)  = \3009(856)  & \2992(969) ,
  \3733(1868)  = \3721(197)  & (\3724(170)  & \4113(1859) ),
  \4453(1712)  = ~\4449(1546) ,
  \4490(2159)  = ~\4484(2114) ,
  \3297(877)  = \479(144)  | (\3296(763)  | \3295(515) ),
  \926(624)  = \1697(357) ,
  \3966(1862)  = ~\5428(1770)  | ~\5425(1470) ,
  \816(628)  = ~\4114(359) ,
  \3237(973)  = ~\3236(860) ,
  \1032(1329)  = ~\4130(1270)  | ~\4127(241) ,
  \760(835)  = \2442(195)  & (\2430(383)  & \67(23) ),
  \5192(1247)  = ~\5186(1085) ,
  \3728(196)  = ~\3724(170) ,
  \1661(601)  = \1633(212)  & (\1609(214)  & \179(78) ),
  \2106(1040)  = ~\3137(914) ,
  \4015(1289)  = \3998(367)  & (\3979(374)  & \2615(1155) ),
  \2089(1039)  = \3137(914) ,
  \4994(2410)  = ~\4988(2391) ,
  \4830(2119)  = ~\4828(2043)  | ~\4825(1761) ,
  \4358(2006)  = ~\4357(1957)  | ~\4356(1901) ,
  \2977(980)  = ~\2976(866) ,
  \4292(239)  = \468(143) ,
  \1578(2101)  = \1564(404)  & (\1528(215)  & \4024(2068) ),
  \1520(2448)  = ~\4627(2446)  | ~\4620(2415) ,
  \685(2316)  = \[115] ,
  \2339(600)  = \2304(208)  & (\2281(210)  & \185(80) ),
  \4796(226)  = \534(149) ,
  \750(831)  = \2442(195)  & (\2430(383)  & \76(26) ),
  \2798(948)  = \2764(587)  | \2763(777) ,
  \5082(262)  = \361(129) ,
  \4570(2056)  = ~\4568(2015)  | ~\4565(1826) ,
  \2158(1501)  = \1984(1423)  & \2099(1419) ,
  \5013(1783)  = ~\5009(1664) ,
  \4795(1208)  = ~\4791(1049) ,
  \2117(1504)  = \1966(1067)  & (\2001(987)  & (\1958(1074)  & \1984(1423) )),
  \2918(533)  = \2882(302)  & \3554(331) ,
  \4073(1286)  = \4056(366)  & (\4037(373)  & \2939(1144) ),
  \880(815)  = \3757(181)  & (\3745(376)  & \118(48) ),
  \5024(2036)  = ~\5022(2017)  | ~\5019(1779) ,
  \4463(1701)  = ~\4459(1538) ,
  \4706(1798)  = ~\4700(1685) ,
  \4666(1209)  = ~\4660(1050) ,
  \720(848)  = \2442(195)  & (\2430(383)  & \11(2) ),
  \5356(347)  = \218(91) ,
  \4803(1205)  = ~\4799(1045) ,
  \1191(1649)  = \1100(1448)  & (\1134(1442)  & (\1116(1446)  & (\1152(1452)  & \4(1) ))),
  \3852(1190)  = \3091(908)  & \3071(1030) ,
  \2794(947)  = \2762(581)  | \2761(774) ,
  \1942(2041)  = \1909(1876)  & \1894(2020) ,
  \1887(2021)  = ~\1886(1975) ,
  \1098(1354)  = ~\4162(1255)  | ~\4159(252) ,
  \5137(922)  = \3147(723) ,
  \1868(1609)  = \1778(1307)  & (\1837(1038)  & (\1794(1406)  & \1812(1404) )),
  \4299(1267)  = ~\4295(1106) ,
  \3234(414)  = \3216(271)  & (\523(148)  & \2405(329) ),
  \730(839)  = \3582(194)  & (\3570(382)  & \46(16) ),
  \2816(353)  = \206(87) ,
  \3130(505)  = \3105(278)  & \323(119) ,
  \1050(1324)  = ~\4138(1266)  | ~\4135(238) ,
  \4159(252)  = \389(136) ,
  \786(653)  = \3684(188)  & (\3660(190)  & \37(13) ),
  \4416(2007)  = ~\4415(1958)  | ~\4414(1902) ,
  \4196(1707)  = \1173(1523)  | (\1172(1557)  | (\1171(1526)  | \1046(1001) )),
  \5033(1787)  = ~\5029(1668) ,
  \3391(697)  = \3369(582)  & (\2370(326)  & \468(143) ),
  \4772(232)  = \503(146) ,
  \2643(311)  = \273(106) ,
  \2647(312)  = \273(106) ,
  \1857(1608)  = \1812(1404)  & (\1767(1417)  & (\1794(1406)  & (\1829(1037)  & \1778(1307) ))),
  \740(827)  = \3582(194)  & (\3570(382)  & \91(35) ),
  \2975(691)  = \2955(502)  & (\3551(199)  & \503(146) ),
  \654(2315)  = \[112] ,
  \1552(213)  = \1690(158) ,
  \756(660)  = \2442(195)  & (\2418(193)  & \17(4) ),
  \777(2278)  = \[107] ,
  \2627(322)  = \257(102) ,
  \4815(1794)  = \2158(1501)  | \2125(1688) ,
  \2788(945)  = \2760(575)  | \2759(773) ,
  \2780(940)  = \2756(558)  | \2755(746) ,
  \4030(183)  = \4091(175) ,
  \1668(599)  = \1633(212)  & (\1609(214)  & \185(80) ),
  \2131(1493)  = \2036(864)  & \2009(1416) ,
  \2784(944)  = \2758(569)  | \2757(770) ,
  \1983(1321)  = ~\4771(1223)  | ~\4764(237) ,
  \4012(1288)  = \3998(367)  & (\3979(374)  & \2619(1171) ),
  \4483(2010)  = ~\4481(1904)  | ~\4474(1964) ,
  \2553(342)  = \226(93) ,
  \4831(2061)  = ~\4829(1855)  | ~\4822(1995) ,
  \4204(1706)  = ~\1175(1556)  & (~\1174(1527)  & ~\1046(1001) ),
  \2593(885)  = \457(142)  | (\2592(666)  | \2590(386) ),
  \2557(337)  = \234(95) ,
  \4714(1797)  = ~\4708(1684) ,
  \818(2273)  = \[90] ,
  \4810(429)  = ~\4804(234) ,
  \2268(2251)  = \2238(400)  & (\2215(402)  & \4085(2232) ),
  \4934(1784)  = ~\4928(1665) ,
  \4626(2421)  = ~\4620(2415) ,
  \4923(1228)  = \1966(1067) ,
  \1195(1605)  = \1160(1034)  & \1134(1442) ,
  \3198(843)  = \3187(397)  & \34(12) ,
  \5072(2392)  = ~\5066(2383) ,
  \5125(1207)  = ~\5121(1048) ,
  \3105(278)  = \332(122) ,
  \3228(424)  = \3208(281)  & (\503(146)  & \2405(329) ),
  \4945(1788)  = ~\4941(1669) ,
  \4203(1708)  = ~\4199(1544) ,
  \4674(1204)  = ~\4668(1044) ,
  \2163(1969)  = ~\2160(1916) ,
  \737(2279)  = \[104] ,
  \2512(379)  = ~\2500(189) ,
  \1792(1303)  = ~\4666(1209)  | ~\4663(228) ,
  \5428(1770)  = ~\5422(1638) ,
  \1810(1300)  = ~\4674(1204)  | ~\4671(227) ,
  \2810(1078)  = ~\2933(933) ,
  \2603(895)  = \422(139)  | (\2602(668)  | \2600(388) ),
  \3925(1815)  = ~\3922(1714) ,
  \3628(187)  = \4091(175) ,
  \1666(2035)  = \1645(403)  & (\1609(214)  & \3790(2025) ),
  \4361(1703)  = \1444(1531)  | (\1443(1562)  | (\1442(1535)  | \1301(1000) )),
  \1672(2100)  = \1645(403)  & (\1609(214)  & \3791(2067) ),
  \4873(1799)  = ~\2125(1688) ,
  \2123(1505)  = \1966(1067)  & (\2001(987)  & \1984(1423) ),
  \4332(247)  = \422(139) ,
  \4138(1266)  = ~\4132(1105) ,
  \1894(2020)  = ~\1893(1972) ,
  \5124(1206)  = ~\5118(1046) ,
  \2124(1506)  = \2001(987)  & \1984(1423) ,
  \1184(1604)  = \1100(1448)  & (\1160(1034)  & (\1089(1436)  & (\1116(1446)  & \1134(1442) ))),
  \2936(1072)  = ~\2908(930) ,
  \4070(1285)  = \4056(366)  & (\4037(373)  & \2942(1137) ),
  \646(2269)  = \1592(607)  | (\1591(789)  | (\1590(2201)  | \1588(2200) )),
  \1823(971)  = \534(149)  & \3139(917) ,
  \5225(1762)  = ~\5223(1629)  | ~\5216(1460) ,
  \1193(1606)  = \1160(1034)  & (\1116(1446)  & \1134(1442) ),
  \4913(1237)  = \1958(1074) ,
  \3949(1843)  = \3926(1667)  & (\3874(1203)  & \3883(1473) ),
  \5133(1201)  = ~\5129(1041) ,
  \651(2314)  = \[111] ,
  \4779(1213)  = ~\4775(1056) ,
  \826(2275)  = \[93] ,
  \728(2250)  = \3594(384)  & (\3570(382)  & \4085(2232) ),
  \746(654)  = \3582(194)  & (\3558(192)  & \37(13) ),
  \4146(1263)  = ~\4140(1102) ,
  \2721(277)  = \335(123) ,
  \3296(763)  = \3267(516)  & \2361(325) ,
  \3339(1162)  = ~\3338(1003) ,
  \4339(1262)  = ~\4335(1101) ,
  \3846(1982)  = \3823(369)  & (\3795(185)  & \1921(1939) ),
  \800(834)  = \2500(189)  & (\2488(381)  & \67(23) ),
  \5022(2017)  = ~\5016(1968) ,
  \1261(2051)  = \1231(1897)  & \1216(1999) ,
  \2276(2253)  = \2238(400)  & (\2203(211)  & \4028(2234) ),
  \2149(1480)  = \2081(970)  & \2042(1408) ,
  \4634(1222)  = ~\4628(1063) ,
  \5077(2441)  = \2195(2429)  | \2194(2439) ,
  \4154(1259)  = ~\4148(1098) ,
  \4534(2419)  = ~\4533(2398)  | ~\4532(2413) ,
  \4544(2418)  = ~\4543(2397)  | ~\4542(2412) ,
  \3946(1835)  = \3922(1714)  & (\3857(1450)  & \3866(1726) ),
  \865(2277)  = \[98] ,
  \595(1463)  = \2810(1078)  & (\2809(1234)  & (\2808(1318)  & \2807(1313) )),
  \3788(1984)  = \3765(371)  & (\3737(186)  & \1243(1961) ),
  \3452(1196)  = ~\5132(1035)  | ~\5129(1041) ,
  \1502(216)  = ~\1497(156) ,
  \4480(2014)  = ~\4474(1964) ,
  \4627(2446)  = ~\4623(2442) ,
  \710(822)  = \3684(188)  & (\3672(380)  & \109(41) ),
  \4211(1709)  = ~\4207(1545) ,
  \3639(2463)  = \3622(372)  & \3658(2460) ,
  \1114(1351)  = ~\4170(1251)  | ~\4167(251) ,
  \4855(1238)  = \1958(1074) ,
  \5169(1258)  = ~\5165(1097) ,
  \3203(951)  = \3202(638)  | \3201(842) ,
  \1000(2168)  = \3543(2120) ,
  \679(2272)  = \[113] ,
  \2945(1079)  = \2933(933) ,
  \3780(816)  = \3757(181)  & (\3745(376)  & \117(47) ),
  \2813(977)  = ~\3015(863) ,
  \1756(1316)  = ~\4642(1219)  | ~\4639(235) ,
  \1429(1358)  = ~\4347(1246)  | ~\4340(256) ,
  \3238(409)  = \3224(264)  & (\534(149)  & \2405(329) ),
  \1448(1698)  = \1447(1565)  | \1318(997) ,
  \4018(1290)  = \3998(367)  & (\3979(374)  & \2611(1159) ),
  \1289(1428)  = ~\1288(1328)  | ~\1287(1160) ,
  \1728(1320)  = ~\4634(1222)  | ~\4631(236) ,
  \4532(2413)  = ~\4530(2396)  | ~\4527(1582) ,
  \4542(2412)  = ~\4618(2395)  | ~\4615(1581) ,
  \3337(886)  = \3325(781)  & (\2382(327)  & \446(141) ),
  \3229(692)  = \3211(500)  & (\2382(327)  & \503(146) ),
  \3836(1120)  = \3823(369)  & (\3803(375)  & \3352(1042) ),
  \1564(404)  = ~\1552(213) ,
  \2147(1476)  = \2021(1306)  & (\2081(970)  & \2042(1408) ),
  \824(2274)  = \[92] ,
  \2120(1503)  = \1966(1067)  & (\2001(987)  & \1984(1423) ),
  \4307(1260)  = ~\4303(1099) ,
  \1878(1647)  = ~\1877(1472)  | ~\1876(1400) ,
  \1869(1645)  = \1778(1307)  & (\1812(1404)  & (\1794(1406)  & (\1829(1037)  & \54(20) ))),
  \1936(2105)  = \1935(1994)  | \1934(2039) ,
  \978(851)  = \1688(663) ,
  \2238(400)  = ~\2226(209) ,
  \2274(2252)  = \2238(400)  & (\2215(402)  & \4086(2231) ),
  \2540(592)  = ~\2537(352) ,
  \3424(913)  = ~\3423(718)  | ~\3422(716) ,
  \4865(1227)  = \1966(1067) ,
  \4988(2391)  = ~\4987(2369)  | ~\4986(2382) ,
  \4013(2027)  = \3998(367)  & (\3972(184)  & \1273(2005) ),
  \4388(2330)  = ~\4387(2306)  | ~\4386(2321) ,
  \4315(1254)  = ~\4311(1093) ,
  \3658(2460)  = \3652(2457)  | \3651(2193) ,
  \4868(2381)  = ~\4862(2368) ,
  \1540(406)  = ~\1528(215) ,
  \4608(2366)  = ~\4602(2355) ,
  \4996(2409)  = ~\5072(2392)  | ~\5069(1487) ,
  \863(2276)  = \[97] ,
  \1190(1603)  = \1100(1448)  & (\1160(1034)  & (\1116(1446)  & \1134(1442) )),
  \3070(909)  = \3069(713)  | \3068(466) ,
  \1686(618)  = \1633(212)  & (\1609(214)  & \146(67) ),
  \4016(2073)  = \3998(367)  & (\3972(184)  & \1268(2050) ),
  \3843(1983)  = \3823(369)  & (\3795(185)  & \1926(1937) ),
  \5224(1756)  = ~\5222(1634)  | ~\5219(1458) ,
  \[3]  = ~\545(150) ,
  \2500(189)  = \4090(174) ,
  \4687(1235)  = \1704(1073) ,
  \4682(648)  = ~\4676(360) ,
  \[4]  = ~\348(126) ,
  \649(2292)  = \1598(610)  | (\1597(791)  | (\1596(2258)  | \1594(2255) )),
  \3328(916)  = \3327(766)  | \3326(475) ,
  \[5]  = ~\366(130) ,
  \1765(1311)  = ~\4650(1212)  | ~\4647(233) ,
  \4071(2026)  = \4056(366)  & (\4030(183)  & \1954(1997) ),
  \[6]  = \562(155)  & \552(152) ,
  \4609(1716)  = ~\4605(1549) ,
  \854(2268)  = \[96] ,
  \3649(2458)  = \3628(187)  & \1524(2454) ,
  \[7]  = ~\549(151) ,
  \[8]  = ~\545(150) ,
  \3785(1985)  = \3765(371)  & (\3737(186)  & \1248(1959) ),
  \4623(2442)  = \1518(2436)  | \1517(2440) ,
  \577(1967)  = ~\1931(1914) ,
  \4162(1255)  = ~\4156(1094) ,
  \[9]  = ~\545(150) ,
  \635(1114)  = \3176(362)  & \3197(953) ,
  \3656(2467)  = \3646(636)  | \3645(2464) ,
  \3943(1834)  = \3918(1715)  & (\3853(1356)  & \3862(1566) ),
  \3196(640)  = \3181(205)  & \86(32) ,
  \4078(812)  = \4049(178)  & (\4037(373)  & \121(51) ),
  \3921(1816)  = ~\3918(1715) ,
  \2691(671)  = \2638(556)  & \3549(200) ,
  \648(2295)  = \[110] ,
  \4291(1269)  = ~\4287(1108) ,
  \4997(2390)  = ~\5073(1662)  | ~\5066(2383) ,
  \2881(678)  = \2847(656)  & \2828(206) ,
  \819(1117)  = \3176(362)  & \3194(954) ,
  \3636(2461)  = \3622(372)  & \3657(2459) ,
  \5235(1772)  = ~\5233(1639)  | ~\5226(1468) ,
  \1197(1650)  = \1152(1452)  & \4(1) ,
  \1944(2104)  = \1943(1992)  | \1942(2041) ,
  \645(2271)  = \[109] ,
  \1596(2258)  = \1564(404)  & (\1528(215)  & \4027(2235) ),
  \5168(1261)  = ~\5162(1100) ,
  \4695(1236)  = \1704(1073) ,
  \1584(2146)  = \1564(404)  & (\1528(215)  & \4025(2129) ),
  \1343(1355)  = ~\4315(1254)  | ~\4308(253) ,
  \2758(569)  = \2734(276)  & \241(96) ,
  \1364(1350)  = ~\4323(1252)  | ~\4316(250) ,
  \4323(1252)  = ~\4319(1091) ,
  \1867(1481)  = \1778(1307)  & (\1823(971)  & \1794(1406) ),
  \3657(2459)  = \3649(2458)  | \3648(2192) ,
  \4116(1112)  = \2802(950) ,
  \4279(1113)  = \2802(950) ,
  \1670(2034)  = \1645(403)  & (\1621(405)  & \3849(2024) ),
  \5303(1297)  = ~\5299(1122) ,
  \3058(906)  = \3057(712)  | \3056(462) ,
  \4947(2038)  = ~\4945(1788)  | ~\4938(1989) ,
  \3645(2464)  = \3622(372)  & \3658(2460) ,
  \813(2260)  = \[91] ,
  \2588(1009)  = ~\2587(891) ,
  \4642(1219)  = ~\4636(1060) ,
  \4170(1251)  = ~\4164(1090) ,
  \4620(2415)  = \1516(2407)  | (\1515(2408)  | (\1514(2406)  | \1513(2405) )),
  \1196(1651)  = \1134(1442)  & (\1152(1452)  & \4(1) ),
  \4397(2345)  = ~\4395(1713)  | ~\4388(2330) ,
  \4599(1730)  = ~\4595(1574) ,
  \3133(732)  = \3112(495)  & \302(114) ,
  \2889(526)  = ~\2886(297) ,
  \5176(1268)  = ~\5170(1107) ,
  \3519(1839)  = \3500(1755)  & (\3454(1453)  & \3449(1624) ),
  \4122(1273)  = ~\4116(1112) ,
  \5234(1771)  = ~\5232(1640)  | ~\5229(1467) ,
  \578(1988)  = ~\1926(1937) ,
  \716(1116)  = \3176(362)  & \3203(951) ,
  \4619(1732)  = ~\4615(1581) ,
  \3239(685)  = \3227(479)  & (\2382(327)  & \534(149) ),
  \2133(1478)  = \2021(1306)  & (\2081(970)  & (\2009(1416)  & \2042(1408) )),
  \4828(2043)  = ~\4822(1995) ,
  \4446(2331)  = ~\4445(2307)  | ~\4444(2322) ,
  \5177(1265)  = ~\5173(1104) ,
  \2869(677)  = \2847(656)  & \2828(206) ,
  \2152(1479)  = \2081(970)  & \2042(1408) ,
  \3782(1986)  = \3765(371)  & (\3737(186)  & \1253(1960) ),
  \2143(1477)  = \2021(1306)  & (\2081(970)  & \2042(1408) ),
  \3310(595)  = \2816(353) ,
  \3654(2468)  = \3640(637)  | \3639(2463) ,
  \4514(2354)  = ~\4513(2332)  | ~\4512(2346) ,
  \1874(1646)  = \1812(1404)  & (\1829(1037)  & \54(20) ),
  \4455(2344)  = ~\4453(1712)  | ~\4446(2331) ,
  \3078(553)  = \3032(315)  & \3554(331) ,
  \3844(814)  = \3815(180)  & (\3803(375)  & \119(49) ),
  \566(1979)  = ~\1200(1934) ,
  \3655(2465)  = \3643(634)  | \3642(2462) ,
  \2270(2254)  = \2238(400)  & (\2203(211)  & \4027(2235) ),
  \2258(2144)  = \2238(400)  & (\2203(211)  & \4025(2129) ),
  \4074(2072)  = \4056(366)  & (\4030(183)  & \1949(2040) ),
  \2708(1352)  = ~\2705(1186) ,
  \4703(1225)  = \1712(1065) ,
  \5004(2422)  = ~\4998(2416) ,
  \4540(2426)  = ~\4534(2419) ,
  \4550(2425)  = ~\4544(2418) ,
  \1877(1472)  = ~\4683(1362)  | ~\4676(360) ,
  \1194(1652)  = \1134(1442)  & (\1116(1446)  & (\1152(1452)  & \4(1) )),
  \3318(596)  = \2816(353) ,
  \3653(2466)  = \3637(635)  | \3636(2461) ,
  \1594(2255)  = \1564(404)  & (\1540(406)  & \4085(2232) ),
  \2886(297)  = \302(114) ,
  \4589(1744)  = ~\4585(1594) ,
  \3646(636)  = \3616(182)  & \94(36) ,
  \3187(397)  = ~\3181(205) ,
  \579(1990)  = ~\1921(1939) ,
  \1150(1360)  = ~\4186(1245)  | ~\4183(257) ,
  \2908(930)  = \2907(764)  | \2906(525) ,
  \3057(712)  = \3031(562)  & (\2370(326)  & \389(136) ),
  \5081(2444)  = ~\5077(2441) ,
  \3947(1963)  = ~\3946(1835)  & ~\3945(1908) ,
  \4568(2015)  = ~\4562(1965) ,
  \628(1853)  = \2135(1673)  & \2113(1632) ,
  \4650(1212)  = ~\4644(1055) ,
  \2678(467)  = \2655(306)  & (\374(134)  & \3553(198) ),
  \2764(587)  = \2734(276)  & \217(90) ,
  \3235(688)  = \3219(488)  & (\2382(327)  & \523(148) ),
  \4739(1674)  = ~\4735(1498) ,
  \2754(551)  = \2721(277)  & \272(105) ,
  \686(2294)  = \2278(612)  | (\2277(792)  | (\2276(2253)  | \2274(2252) )),
  \5116(731)  = ~\5114(530)  | ~\5111(296) ,
  \637(965)  = \2881(678)  | (\2880(684)  | (\2879(960)  | \2878(961) )),
  \4283(1274)  = ~\4279(1113) ,
  \3332(1163)  = ~\3331(1005) ,
  \1582(2145)  = \1564(404)  & (\1540(406)  & \4083(2130) ),
  \3484(1241)  = ~\5184(1080)  | ~\5181(1111) ,
  \5106(728)  = ~\5104(514)  | ~\5101(289) ,
  \3295(515)  = \3264(291)  & \3555(332) ,
  \3952(1844)  = \3930(1666)  & (\3878(1367)  & \3887(1654) ),
  \1697(357)  = \137(63) ,
  \4082(2071)  = \4069(837)  | (\4068(1980)  | \4067(1284) ),
  \703(1115)  = \3176(362)  & \3200(952) ,
  \4130(1270)  = ~\4124(1109) ,
  \1872(1648)  = \1812(1404)  & (\1794(1406)  & (\1829(1037)  & \54(20) )),
  \4944(2037)  = ~\4938(1989) ,
  \2753(743)  = \2728(494)  & \265(104) ,
  \4024(2068)  = \4011(811)  | (\4010(1981)  | \4009(1287) ),
  \4014(820)  = \3991(179)  & (\3979(374)  & \113(43) ),
  \3642(2462)  = \3622(372)  & \3657(2459) ,
  \727(2298)  = \[102] ,
  \4394(2342)  = ~\4388(2330) ,
  \5247(1847)  = ~\5225(1762)  | ~\5224(1756) ,
  \2638(556)  = ~\2635(317) ,
  \2630(563)  = ~\2627(322) ,
  \2256(2143)  = \2238(400)  & (\2215(402)  & \4083(2130) ),
  \2634(564)  = ~\2631(323) ,
  \3259(532)  = ~\3256(301) ,
  \4711(1224)  = \1712(1065) ,
  \2132(1489)  = \2059(975)  & (\2009(1416)  & \2021(1306) ),
  \713(967)  = \2873(680)  | (\2872(682)  | (\2871(957)  | \2870(955) )),
  \5405(1264)  = ~\5403(1103)  | ~\5396(1110) ,
  \3731(1121)  = \3721(197)  & (\3728(196)  & \2945(1079) ),
  \1365(1445)  = ~\1364(1350)  | ~\1363(1184) ,
  \5203(1250)  = ~\5199(1089) ,
  \5074(2414)  = \2193(2403)  | (\2192(2404)  | (\2191(2402)  | \2190(2401) )),
  \2728(494)  = ~\2721(277) ,
  \4523(2364)  = ~\4521(1717)  | ~\4514(2354) ,
  \4849(1686)  = ~\4845(1516) ,
  \1064(996)  = \468(143)  & \2794(947) ,
  \1332(1435)  = ~\1331(1336)  | ~\1330(1168) ,
  \2570(999)  = ~\2569(884) ,
  \1278(1433)  = ~\1277(1333)  | ~\1276(1165) ,
  \4611(2363)  = ~\4609(1716)  | ~\4602(2355) ,
  \3147(723)  = \3126(492)  | \3099(496) ,
  \4886(2044)  = ~\4880(1996) ,
  \1843(1630)  = \1704(1073)  & (\1730(1422)  & (\1758(1420)  & \1712(1065) )),
  \603(225)  = \[8] ,
  \4452(2343)  = ~\4446(2331) ,
  \4951(1200)  = \2106(1040) ,
  \2747(737)  = \2728(494)  & \289(110) ,
  \4444(2322)  = ~\4442(2308)  | ~\4439(1532) ,
  \4918(2356)  = ~\4916(2341)  | ~\4913(1237) ,
  \4386(2321)  = ~\4384(2309)  | ~\4381(1529) ,
  \3055(538)  = ~\3052(304) ,
  \1217(1723)  = ~\4234(1174)  | ~\4231(1521) ,
  \1307(1427)  = ~\1306(1325)  | ~\1305(1157) ,
  \2226(209)  = \1694(160) ,
  \1344(1449)  = ~\1343(1355)  | ~\1342(1189) ,
  \5026(2102)  = ~\5025(1987)  | ~\5024(2036) ,
  \4555(1734)  = ~\1476(1601)  & (~\1475(1579)  & ~\1382(1024) ),
  \3652(2457)  = \3628(187)  & \2201(2453) ,
  \4811(1218)  = ~\4807(1059) ,
  \5402(1271)  = ~\5396(1110) ,
  \5185(1272)  = ~\5181(1111) ,
  \4020(819)  = \3991(179)  & (\3979(374)  & \114(44) ),
  \4771(1223)  = ~\4767(1064) ,
  \2660(461)  = \2631(323)  & (\389(136)  & \3553(198) ),
  \5355(559)  = ~\5351(319) ,
  \2578(450)  = \2553(342)  & (\422(139)  & \3553(198) ),
  \2564(573)  = ~\2561(336) ,
  \4602(2355)  = ~\4601(2333)  | ~\4600(2347) ,
  \2041(1304)  = ~\4795(1208)  | ~\4788(229) ,
  \4679(1197)  = \1829(1037) ,
  \1089(1436)  = ~\1088(1169)  | ~\1087(1337) ,
  \680(2270)  = \2266(608)  | (\2265(788)  | (\2264(2199)  | \2262(2198) )),
  \683(2291)  = \2272(609)  | (\2271(790)  | (\2270(2254)  | \2268(2251) )),
  \4618(2395)  = ~\4612(2386) ,
  \5104(514)  = ~\5098(290) ,
  \2760(575)  = \2734(276)  & \233(94) ,
  \2548(584)  = ~\2545(345) ,
  \4839(1679)  = ~\4835(1502) ,
  \2560(574)  = ~\2557(337) ,
  \3913(745)  = ~\5354(572)  | ~\5351(319) ,
  \5202(1253)  = ~\5196(1092) ,
  \4521(1717)  = ~\4517(1550) ,
  \3944(1962)  = ~\3943(1834)  & ~\3942(1909) ,
  \2676(1018)  = ~\2675(896) ,
  \4708(1684)  = ~\1856(1513)  & ~\1742(992) ,
  \3128(497)  = \3105(278)  & \331(121) ,
  \5319(1312)  = ~\5315(1136) ,
  \3051(540)  = ~\3048(305) ,
  \1602(2257)  = \1564(404)  & (\1528(215)  & \4028(2234) ),
  \2544(585)  = ~\2541(346) ,
  \682(2296)  = \[114] ,
  \4978(2360)  = ~\4977(2339)  | ~\4976(2351) ,
  \1116(1446)  = ~\1115(1185)  | ~\1114(1351) ,
  \4987(2369)  = ~\4985(1663)  | ~\4978(2360) ,
  \1478(1731)  = \1477(1600)  | \1404(1021) ,
  \2664(1026)  = ~\2663(904) ,
  \5080(2420)  = ~\5074(2414) ,
  \1860(1486)  = \1806(974)  & (\1767(1417)  & \1778(1307) ),
  \4111(1765)  = \4107(1644)  & \4104(1462) ,
  \3423(718)  = ~\5089(471)  | ~\5082(262) ,
  \2350(800)  = \2304(208)  & (\2293(401)  & \155(70) ),
  \4387(2306)  = ~\4385(1695)  | ~\4378(2284) ,
  \4976(2351)  = ~\4974(2337)  | ~\4971(1497) ,
  \2021(1306)  = ~\2020(1130)  | ~\2019(978) ,
  \1861(1482)  = \1778(1307)  & (\1823(971)  & (\1767(1417)  & \1794(1406) )),
  \3271(517)  = ~\3268(292) ,
  \4575(1742)  = ~\1471(1598)  & (~\1470(1576)  & (~\1469(1583)  & ~\1359(1029) )),
  \2999(419)  = \514(147)  | \3547(201) ,
  \3127(724)  = \3112(495)  & \324(120) ,
  \4862(2368)  = ~\4861(2349)  | ~\4860(2357) ,
  \4112(1774)  = \132(60)  & \4107(1644) ,
  \3937(1256)  = ~\3934(1095) ,
  \4897(1678)  = ~\4893(1500) ,
  \652(2293)  = \1604(611)  | (\1603(793)  | (\1602(2257)  | \1600(2256) )),
  \2885(534)  = ~\2882(302) ,
  \3092(279)  = \332(122) ,
  \5338(543)  = ~\5332(308) ,
  \718(1867)  = \2454(385)  & (\2430(383)  & \3848(1864) ),
  \1526(622)  = \1697(357) ,
  \1134(1442)  = ~\1133(1180)  | ~\1132(1346) ,
  \4520(2365)  = ~\4514(2354) ,
  \1851(1631)  = \1712(1065)  & (\1730(1422)  & \1758(1420) ),
  \1422(1439)  = ~\1421(1342)  | ~\1420(1175) ,
  \4524(2387)  = ~\4523(2364)  | ~\4522(2377) ,
  \3838(804)  = \3815(180)  & (\3803(375)  & \131(59) ),
  \3948(1919)  = \3929(1786)  & (\3883(1473)  & \3878(1367) ),
  \855(1866)  = \2512(379)  & (\2488(381)  & \3848(1864) ),
  \772(2299)  = \[106] ,
  \1915(1790)  = ~\4739(1674)  | ~\4732(1670) ,
  \4511(1729)  = ~\4507(1571) ,
  \3064(454)  = \3044(310)  & (\411(138)  & \2393(328) ),
  \4612(2386)  = ~\4611(2363)  | ~\4610(2376) ,
  \4522(2377)  = ~\4520(2365)  | ~\4517(1550) ,
  \1870(1483)  = \1794(1406)  & \1823(971) ,
  \2979(420)  = \514(147)  & \3553(198) ,
  \2202(626)  = \1698(358) ,
  \4531(1733)  = ~\4527(1582) ,
  \4445(2307)  = ~\4443(1697)  | ~\4436(2283) ,
  \1600(2256)  = \1564(404)  & (\1540(406)  & \4086(2231) ),
  \785(840)  = \3684(188)  & (\3672(380)  & \43(15) ),
  \5114(530)  = ~\5108(300) ,
  \5376(1808)  = ~\5295(1536)  | ~\5294(1699) ,
  \1873(1611)  = \1837(1038)  & \1812(1404) ,
  \3202(638)  = \3181(205)  & \88(34) ,
  \4748(1658)  = \1874(1646)  | (\1873(1611)  | \1823(971) ),
  \842(368)  = \3815(180)  & \3795(185) ,
  \4079(1119)  = \4056(366)  & (\4037(373)  & \2945(1079) ),
  \3060(457)  = \3036(314)  & (\400(137)  & \2393(328) ),
  \1597(791)  = \1552(213)  & (\1540(406)  & \194(83) ),
  \5318(1319)  = ~\5312(1145) ,
  \3522(1845)  = \3504(1754)  & (\3458(1607)  & \3445(1455) ),
  \712(2297)  = \[101] ,
  \5089(471)  = ~\5085(258) ,
  \3533(1846)  = ~\3532(1627)  | ~\3531(1757) ,
  \5412(2057)  = ~\5406(2013) ,
  \3290(984)  = ~\3289(871) ,
  \3489(504)  = \3440(284) ,
  \1592(607)  = \1552(213)  & (\1528(215)  & \167(74) ),
  \3839(1291)  = \3823(369)  & (\3803(375)  & \3021(1123) ),
  \1390(1443)  = ~\1389(1347)  | ~\1388(1181) ,
  \4287(1108)  = \2798(948) ,
  \3299(507)  = \3272(286)  & \3555(332) ,
  \1458(1719)  = \1457(1597)  | (\1456(1578)  | (\1455(1585)  | (\1454(1593)  | \1341(1010) ))),
  \5343(313)  = \273(106) ,
  \3787(1296)  = \3765(371)  & (\3745(376)  & \2705(1186) ),
  \3378(334)  = \234(95) ,
  \3953(1971)  = ~\3952(1844)  & ~\3951(1918) ,
  \2878(961)  = \2857(844)  & (\2838(398)  & \24(7) ),
  \3778(1293)  = \3765(371)  & (\3745(376)  & \2717(1191) ),
  \1185(1721)  = \1184(1604)  | (\1183(1568)  | (\1182(1588)  | (\1181(1590)  | \1097(1011) ))),
  \1606(623)  = \1697(357) ,
  \2701(673)  = \2654(542)  & \3549(200) ,
  \5293(1326)  = ~\5289(1158) ,
  \4571(2011)  = ~\4569(1905)  | ~\4562(1965) ,
  \5014(1841)  = ~\5012(1364)  | ~\5009(1664) ,
  \4384(2309)  = ~\4378(2284) ,
  \5266(1348)  = ~\5260(1182) ,
  \5267(1345)  = ~\5263(1179) ,
  \795(833)  = \2500(189)  & (\2488(381)  & \73(25) ),
  \2008(1310)  = ~\4779(1213)  | ~\4772(232) ,
  \1862(1610)  = \1778(1307)  & (\1837(1038)  & (\1767(1417)  & (\1794(1406)  & \1812(1404) ))),
  \[100]  = ~\4025(2129) ,
  \1903(1793)  = \1902(1775)  | \1863(1675) ,
  \[101]  = \711(630)  | (\710(822)  | (\709(2245)  | \708(2243) )),
  \1318(997)  = \2794(947)  & \468(143) ,
  \3991(179)  = \4092(176) ,
  \3068(466)  = \3052(304)  & (\374(134)  & \2393(328) ),
  \[102]  = \726(631)  | (\725(823)  | (\724(2247)  | \723(2249) )),
  \765(847)  = \2442(195)  & (\2430(383)  & \14(3) ),
  \2582(1013)  = ~\2581(894) ,
  \4335(1101)  = \2788(945) ,
  \4364(2053)  = ~\4358(2006) ,
  \4541(1741)  = ~\4537(1592) ,
  \4501(1745)  = ~\4497(1595) ,
  \1929(1751)  = ~\4762(1454)  | ~\4759(1484) ,
  \[103]  = \731(650)  | (\730(839)  | (\729(2248)  | \728(2250) )),
  \1859(1495)  = \1789(865)  & \1767(1417) ,
  \3276(285)  = \316(118) ,
  \[104]  = \736(633)  | (\735(825)  | (\734(2196)  | \733(2197) )),
  \4533(2398)  = ~\4531(1733)  | ~\4524(2387) ,
  \[105]  = \741(651)  | (\740(827)  | (\739(2140)  | \738(2141) )),
  \3194(954)  = \3193(641)  | \3192(829) ,
  \[106]  = \771(649)  | (\770(838)  | (\769(2246)  | \768(2244) )),
  \4107(1644)  = ~\132(60)  | ~\4104(1462) ,
  \3551(199)  = ~\3550(167) ,
  \4543(2397)  = ~\4619(1732)  | ~\4612(2386) ,
  \4155(448)  = ~\4151(245) ,
  \[107]  = \776(632)  | (\775(824)  | (\774(2195)  | \773(2194) )),
  \3462(1210)  = ~\5141(1053)  | ~\5134(1054) ,
  \3418(568)  = \3378(334)  & \3554(331) ,
  \4860(2357)  = ~\4858(2340)  | ~\4855(1238) ,
  \4848(2303)  = ~\4842(2282) ,
  \2874(959)  = \2857(844)  & (\2838(398)  & \26(9) ),
  \839(2241)  = \3823(369)  & (\3803(375)  & \3835(2206) ),
  \699(2227)  = \[88] ,
  \[108]  = \781(652)  | (\780(826)  | (\779(2139)  | \778(2138) )),
  \2098(1314)  = ~\4811(1218)  | ~\4804(234) ,
  \4732(1670)  = \1869(1645)  | (\1868(1609)  | (\1867(1481)  | (\1866(1407)  | \1789(865) ))),
  \1128(1025)  = \400(137)  & \2776(939) ,
  \4551(1740)  = ~\4547(1591) ,
  \[109]  = \1526(622)  & \643(2221) ,
  \1667(797)  = \1633(212)  & (\1621(405)  & \182(79) ),
  \3968(1930)  = ~\3967(1769)  | ~\3966(1862) ,
  \4723(1683)  = ~\4719(1515) ,
  \2272(609)  = \2226(209)  & (\2203(211)  & \164(73) ),
  \853(2202)  = \3970(1978)  & (\3535(1921)  & (\3545(2169)  & (\3540(2164)  & \562(155) ))),
  \2720(1357)  = ~\2717(1191) ,
  \1871(1612)  = \1837(1038)  & (\1794(1406)  & \1812(1404) ),
  \812(2205)  = \1936(2105)  & \4096(2167) ,
  \1586(604)  = \1552(213)  & (\1528(215)  & \173(76) ),
  \3370(339)  = \226(93) ,
  \5420(2058)  = ~\5414(2018) ,
  \1046(1001)  = \457(142)  & \2798(948) ,
  \3536(2059)  = ~\5250(2016)  | ~\5247(1847) ,
  \3279(506)  = ~\3276(285) ,
  \2370(326)  = \251(100) ,
  \1221(1722)  = ~\4242(1341)  | ~\4239(1520) ,
  \[110]  = \1526(622)  & \646(2269) ,
  \4131(442)  = ~\4127(241) ,
  \4442(2308)  = ~\4436(2283) ,
  \2277(792)  = \2226(209)  & (\2215(402)  & \191(82) ),
  \3970(1978)  = ~\3968(1930) ,
  \[111]  = \1526(622)  & \649(2292) ,
  \1673(794)  = \1633(212)  & (\1621(405)  & \188(81) ),
  \4926(2380)  = ~\4920(2367) ,
  \4295(1106)  = \2794(947) ,
  \3272(286)  = \316(118) ,
  \[112]  = \1526(622)  & \652(2293) ,
  \607(1425)  = \2614(1327)  & (\2618(1323)  & (\2622(1339)  & \2626(1335) )),
  \1023(1432)  = ~\1022(1164)  | ~\1021(1332) ,
  \[113]  = \2202(626)  & \677(2220) ,
  \4076(1118)  = \4056(366)  & (\4037(373)  & \2936(1072) ),
  \3374(340)  = \226(93) ,
  \2266(608)  = \2226(209)  & (\2203(211)  & \167(74) ),
  \4610(2376)  = ~\4608(2366)  | ~\4605(1549) ,
  \5282(1322)  = ~\5276(1154) ,
  \3408(566)  = \3362(344)  & \3554(331) ,
  \769(2246)  = \3696(378)  & (\3660(190)  & \4027(2235) ),
  \3275(508)  = ~\3272(286) ,
  \[114]  = \2202(626)  & \680(2270) ,
  \[115]  = \2202(626)  & \683(2291) ,
  \3795(185)  = \4091(175) ,
  \[116]  = \2202(626)  & \686(2294) ,
  \4037(373)  = ~\4030(183) ,
  \2870(955)  = \2857(844)  & (\2838(398)  & \82(30) ),
  \4984(2371)  = ~\4978(2360) ,
  \4968(2326)  = ~\4967(2301)  | ~\4966(2318) ,
  \4908(2320)  = ~\4906(2302)  | ~\4903(1517) ,
  \580(1991)  = ~\1916(1940) ,
  \3779(1936)  = \3765(371)  & (\3737(186)  & \1200(1934) ),
  \709(2245)  = \3696(378)  & (\3660(190)  & \4028(2234) ),
  \[117]  = \842(368)  | (\841(813)  | (\840(2451)  | \839(2241) )),
  \5178(934)  = \2748(535)  | \2747(737) ,
  \4338(452)  = ~\4332(247) ,
  \2670(1023)  = ~\2669(903) ,
  \[118]  = \881(370)  | (\880(815)  | (\879(2452)  | \878(2242) )),
  \[119]  = \766(644)  | (\765(847)  | (\764(2471)  | \763(2472) )),
  \4986(2382)  = ~\4984(2371)  | ~\4981(1488) ,
  \4928(1665)  = \2151(1622)  | (\2150(1616)  | (\2149(1480)  | \2059(975) )),
  \1100(1448)  = ~\1099(1188)  | ~\1098(1354) ,
  \4552(1194)  = \1412(1033) ,
  \3950(1970)  = ~\3949(1843)  & ~\3948(1919) ,
  \878(2242)  = \3765(371)  & (\3745(376)  & \3777(2209) ),
  \2537(352)  = \210(89) ,
  \4763(1659)  = ~\4759(1484) ,
  \4651(426)  = ~\4647(233) ,
  \745(841)  = \3582(194)  & (\3570(382)  & \43(15) ),
  \4314(464)  = ~\4308(253) ,
  \828(2233)  = \[94] ,
  \1900(1795)  = ~\4731(1682)  | ~\4724(1142) ,
  \4966(2318)  = ~\4964(2313)  | ~\4961(1474) ,
  \2533(351)  = \210(89) ,
  \2901(511)  = ~\2898(288) ,
  \4422(2054)  = ~\4416(2007) ,
  \5093(268)  = \351(127) ,
  \3554(331)  = \242(97) ,
  \677(2220)  = \2260(603)  | (\2259(784)  | (\2258(2144)  | \2256(2143) )),
  \1359(1029)  = \2780(940)  & \389(136) ,
  \845(845)  = \[19] ,
  \4755(1660)  = ~\4751(1485) ,
  \[120]  = \806(645)  | (\805(846)  | (\804(2470)  | \803(2469) )),
  \596(1412)  = \2814(1308)  & (\2813(977)  & (\2812(1301)  & \2811(1298) )),
  \4731(1682)  = ~\4727(1514) ,
  \775(824)  = \3684(188)  & (\3672(380)  & \100(38) ),
  \[121]  = ~\657(2481) ,
  \892(408)  = \3175(221) ,
  \4675(412)  = ~\4671(227) ,
  \729(2248)  = \3594(384)  & (\3558(192)  & \4027(2235) ),
  \[122]  = ~\689(2482) ,
  \676(2229)  = \[86] ,
  \1866(1407)  = \1806(974)  & \1778(1307) ,
  \708(2243)  = \3696(378)  & (\3672(380)  & \4086(2231) ),
  \4659(422)  = ~\4655(231) ,
  \3784(1295)  = \3765(371)  & (\3745(376)  & \2709(1183) ),
  \3941(1257)  = ~\3938(1096) ,
  \1034(1429)  = ~\1033(1161)  | ~\1032(1329) ,
  \608(1440)  = \2708(1352)  & (\2712(1349)  & (\2716(1344)  & \2720(1357) )),
  \3721(197)  = ~\3717(169) ,
  \696(2226)  = \[87] ,
  \4530(2396)  = ~\4524(2387) ,
  \3862(1566)  = ~\3861(1444)  | ~\3860(1441) ,
  \1704(1073)  = ~\3167(931) ,
  \667(2224)  = \[84] ,
  \4482(2055)  = ~\4480(2014)  | ~\4477(1825) ,
  \867(2237)  = \[99] ,
  \755(832)  = \2442(195)  & (\2430(383)  & \73(25) ),
  \2332(602)  = \2304(208)  & (\2281(210)  & \179(78) ),
  \4139(437)  = ~\4135(238) ,
  \3951(1918)  = \3933(1785)  & (\3887(1654)  & \3874(1203) ),
  \4330(456)  = ~\4324(249) ,
  \5035(2148)  = ~\5033(1787)  | ~\5026(2102) ,
  \4635(433)  = ~\4631(236) ,
  \1145(1020)  = \411(138)  & \2772(937) ,
  \609(1430)  = ~\3350(1331) ,
  \1876(1400)  = ~\4682(648)  | ~\4679(1197) ,
  \5283(1338)  = ~\5279(1170) ,
  \1052(1426)  = ~\1051(1156)  | ~\1050(1324) ,
  \768(2244)  = \3696(378)  & (\3672(380)  & \4085(2232) ),
  \5274(1334)  = ~\5268(1166) ,
  \2682(1031)  = ~\2681(911) ,
  \923(619)  = \1701(355) ,
  \1453(1718)  = ~\1451(1551) ,
  \3388(882)  = \3387(699)  | \3386(439) ,
  \4700(1685)  = \1855(1507)  | (\1854(1512)  | \1742(992) ),
  \817(2230)  = \3735(2142)  | (\3734(629)  | (\3733(1868)  | \3731(1121) )),
  \3803(375)  = ~\3795(185) ,
  \2681(911)  = \2680(714)  | \2678(467) ,
  \3354(349)  = \210(89) ,
  \4977(2339)  = ~\4975(1672)  | ~\4968(2326) ,
  \2955(502)  = ~\2952(283) ,
  \1080(1438)  = ~\1079(1172)  | ~\1078(1340) ,
  \2952(283)  = \324(120) ,
  \4920(2367)  = ~\4919(2348)  | ~\4918(2356) ,
  \4965(1655)  = ~\4961(1474) ,
  \5374(949)  = ~\5372(782)  | ~\5369(348) ,
  \3216(271)  = \341(125) ,
  \4124(1109)  = \2798(948) ,
  \3212(270)  = \341(125) ,
  \4919(2348)  = ~\4917(1383)  | ~\4910(2329) ,
  \4759(1484)  = \1812(1404) ,
  \2598(880)  = \468(143)  | (\2597(667)  | \2595(387) ),
  \4964(2313)  = ~\4958(2290) ,
  \2951(501)  = ~\2948(282) ,
  \5379(1518)  = ~\5285(1424)  | ~\5284(1437) ,
  \4132(1105)  = \2794(947) ,
  \3823(369)  = ~\3815(180) ,
  \591(1894)  = \[51] ,
  \2956(272)  = \341(125) ,
  \1588(2200)  = \1564(404)  & (\1540(406)  & \4084(2180) ),
  \3044(310)  = \273(106) ,
  \3842(1292)  = \3823(369)  & (\3803(375)  & \3018(1126) ),
  \629(1926)  = \[54] ,
  \805(846)  = \2500(189)  & (\2488(381)  & \14(3) ),
  \618(1925)  = \[52] ,
  \1404(1021)  = \2772(937)  & \411(138) ,
  \2264(2199)  = \2238(400)  & (\2203(211)  & \4026(2185) ),
  \4049(178)  = \4092(176) ,
  \664(2223)  = \[83] ,
  \3781(1294)  = \3765(371)  & (\3745(376)  & \2713(1178) ),
  \4985(1663)  = ~\4981(1488) ,
  \621(1893)  = \[53] ,
  \643(2221)  = \1586(604)  | (\1585(785)  | (\1584(2146)  | \1582(2145) )),
  \4143(246)  = \422(139) ,
  \1412(1033)  = \2767(936)  & \374(134) ,
  \610(1519)  = \[44] ,
  \2814(1308)  = ~\3012(1132) ,
  \3874(1203)  = ~\3348(1043) ,
  \1978(1068)  = \3165(927) ,
  \4663(228)  = \523(148) ,
  \2608(890)  = \435(140)  | (\2607(669)  | \2605(389) ),
  \3524(1913)  = ~\3523(1749)  & ~\3522(1845) ,
  \2592(666)  = \2536(591)  & \3549(200) ,
  \3541(2062)  = ~\5258(2022)  | ~\5255(1860) ,
  \3878(1367)  = ~\3874(1203) ,
  \3527(1932)  = ~\3526(1773)  & ~\3525(1863) ,
  \782(2239)  = \[108] ,
  \814(203)  = ~\3173(164) ,
  \5032(2147)  = ~\5026(2102) ,
  \735(825)  = \3582(194)  & (\3570(382)  & \100(38) ),
  \4907(1687)  = ~\4903(1517) ,
  \1794(1406)  = ~\1793(1128)  | ~\1792(1303) ,
  \3958(1243)  = \3938(1096)  & (\3901(1081)  & \3910(1088) ),
  \1324(1017)  = \2788(945)  & \422(139) ,
  \3211(500)  = ~\3208(281) ,
  \1031(1006)  = \446(141)  & \2802(950) ,
  \869(2181)  = \[100] ,
  \4740(1661)  = \1872(1648)  | (\1871(1612)  | (\1870(1483)  | \1806(974) )),
  \4995(1492)  = ~\4991(1414) ,
  \3518(1371)  = ~\3517(1214)  & ~\3516(1215) ,
  \642(2222)  = \[82] ,
  \1812(1404)  = ~\1811(1125)  | ~\1810(1300) ,
  \585(2236)  = \[71] ,
  \2618(1323)  = ~\2615(1155) ,
  \1896(1796)  = ~\4723(1683)  | ~\4716(989) ,
  \4858(2340)  = ~\4852(2328) ,
  \1633(212)  = \1690(158) ,
  \4916(2341)  = ~\4910(2329) ,
  \4127(241)  = \457(142) ,
  \4974(2337)  = ~\4968(2326) ,
  \724(2247)  = \3594(384)  & (\3558(192)  & \4028(2234) ),
  \4647(233)  = \503(146) ,
  \3535(1921)  = ~\3533(1846) ,
  \2812(1301)  = ~\3018(1126) ,
  \4140(1102)  = \2788(945) ,
  \4975(1672)  = ~\4971(1497) ,
  \841(813)  = \3815(180)  & (\3803(375)  & \120(50) ),
  \1984(1423)  = ~\1983(1321)  | ~\1982(1150) ,
  \1603(793)  = \1552(213)  & (\1540(406)  & \191(82) ),
  \2262(2198)  = \2238(400)  & (\2215(402)  & \4084(2180) ),
  \725(823)  = \3582(194)  & (\3570(382)  & \109(41) ),
  \742(2238)  = \[105] ,
  \5023(1871)  = ~\5019(1779) ,
  \594(224)  = \[3] ,
  \2018(982)  = \3151(923)  & \503(146) ,
  \3517(1214)  = \3493(503)  & (\3428(1036)  & \3437(1047) ),
  \1966(1067)  = ~\3165(927) ,
  \4851(2304)  = ~\4849(1686)  | ~\4842(2282) ,
  \3954(1392)  = \3937(1256)  & (\3906(938)  & \3901(1081) ),
  \5302(1302)  = ~\5296(1127) ,
  \3793(2065)  = \3789(807)  | (\3788(1984)  | \3787(1296) ),
  \1111(1028)  = \389(136)  & \2780(940) ,
  \1724(1066)  = \3165(927) ,
  \1925(1780)  = ~\4755(1660)  | ~\4748(1658) ,
  \723(2249)  = \3594(384)  & (\3570(382)  & \4086(2231) ),
  \3792(2066)  = \3786(808)  | (\3785(1985)  | \3784(1295) ),
  \3028(321)  = \257(102) ,
  \2902(287)  = \316(118) ,
  \3851(2063)  = \3847(805)  | (\3846(1982)  | \3845(963) ),
  \3850(2069)  = \3844(814)  | (\3843(1983)  | \3842(1292) ),
  \3200(952)  = \3199(639)  | \3198(843) ,
  \3815(180)  = \4092(176) ,
  \3024(320)  = \257(102) ,
  \1341(1010)  = \2784(944)  & \435(140) ,
  \4316(250)  = \400(137) ,
  \3155(924)  = \3130(505)  | \3129(727) ,
  \3293(761)  = \3259(532)  & \2361(325) ,
  \2905(509)  = ~\2902(287) ,
  \3353(1330)  = \3347(1002)  & \3339(1162) ,
  \575(2240)  = \[70] ,
  \2115(1229)  = \1978(1068)  & \1958(1074) ,
  \3091(908)  = \374(134)  | (\3090(753)  | \3088(539) ),
  \3165(927)  = \3134(521)  | \3133(732) ,
  \1958(1074)  = ~\3167(931) ,
  \3515(1372)  = ~\3514(1057)  & ~\3513(1216) ,
  \3151(923)  = \3128(497)  | \3127(724) ,
  \3361(590)  = ~\3358(350) ,
  \3161(926)  = \3132(513)  | \3131(730) ,
  \3516(1215)  = \3496(725)  & (\3437(1047)  & \3424(913) ),
  \3081(900)  = \400(137)  | (\3080(751)  | \3078(553) ),
  \3335(915)  = \3334(765)  | \3333(473) ,
  \1712(1065)  = ~\3165(927) ,
  \3521(1912)  = ~\3520(1748)  & ~\3519(1839) ,
  \1902(1775)  = \54(20)  & \1857(1608) ,
  \2909(431)  = \2894(294)  & (\479(144)  & \2393(328) ),
  \3955(1242)  = \3934(1095)  & (\3897(935)  & \3906(938) ),
  \787(2186)  = \[78] ,
  \3791(2067)  = \3783(809)  | (\3782(1986)  | \3781(1294) ),
  \3240(855)  = \3239(685)  | \3238(409) ,
  \4941(1669)  = \2145(1620)  | (\2144(1613)  | (\2143(1477)  | (\2142(1410)  | \2036(864) ))),
  \670(2225)  = \[85] ,
  \1286(1007)  = \2802(950)  & \446(141) ,
  \4818(1139)  = ~\4812(986) ,
  \4069(837)  = \4049(178)  & (\4037(373)  & \52(18) ),
  \3385(570)  = ~\3382(333) ,
  \3048(305)  = \281(108) ,
  \4909(2305)  = ~\4907(1687)  | ~\4900(2281) ,
  \4598(2334)  = ~\4592(2323) ,
  \3139(917)  = \3123(478)  | \3122(719) ,
  \4971(1497)  = \2009(1416) ,
  \1382(1024)  = \2776(939)  & \400(137) ,
  \3302(261)  = \361(129) ,
  \3330(887)  = \3313(779)  & (\2382(327)  & \446(141) ),
  \3381(571)  = ~\3378(334) ,
  \789(2078)  = \2512(379)  & (\2476(191)  & \3793(2065) ),
  \4021(1401)  = \3998(367)  & (\3979(374)  & \3353(1330) ),
  \5195(1391)  = ~\5193(1244)  | ~\5186(1085) ,
  \2716(1344)  = ~\2713(1178) ,
  \747(2187)  = \[74] ,
  \5417(1877)  = ~\5395(1856)  | ~\5394(1676) ,
  \4081(810)  = \4049(178)  & (\4037(373)  & \123(53) ),
  \574(2158)  = ~\1258(2112) ,
  \3195(828)  = \3187(397)  & \87(33) ,
  \4910(2329)  = ~\4909(2305)  | ~\4908(2320) ,
  \5255(1860)  = ~\5235(1772)  | ~\5234(1771) ,
  \4354(1176)  = ~\4348(1016) ,
  \2203(211)  = \1691(159) ,
  \1160(1034)  = \374(134)  & \2767(936) ,
  \5310(1309)  = ~\5304(1133) ,
  \3099(496)  = ~\3092(279) ,
  \3040(309)  = \273(106) ,
  \1767(1417)  = ~\1766(1135)  | ~\1765(1311) ,
  \5295(1536)  = ~\5293(1326)  | ~\5286(1431) ,
  \3915(941)  = ~\3914(771)  | ~\3913(745) ,
  \606(407)  = \[26] ,
  \3945(1908)  = \3925(1815)  & (\3866(1726)  & \3853(1356) ),
  \5205(1394)  = ~\5203(1250)  | ~\5196(1092) ,
  \4235(1691)  = ~\4231(1521) ,
  \4406(1177)  = \1324(1017) ,
  \668(2177)  = \1686(618)  | (\1685(802)  | (\1684(2098)  | \1682(2096) )),
  \4398(2362)  = ~\4397(2345)  | ~\4396(2353) ,
  \584(2151)  = ~\1936(2105) ,
  \5194(1390)  = ~\5192(1247)  | ~\5189(1082) ,
  \2680(714)  = \2658(541)  & (\3551(199)  & \374(134) ),
  \1645(403)  = ~\1633(212) ,
  \2763(777)  = \2741(493)  & \210(89) ,
  \2996(674)  = \2951(501)  & \3549(200) ,
  \1097(1011)  = \435(140)  & \2784(944) ,
  \3840(1935)  = \3823(369)  & (\3795(185)  & \1931(1914) ),
  \4404(2375)  = ~\4398(2362) ,
  \2696(672)  = \2646(548)  & \3549(200) ,
  \2215(402)  = ~\2203(211) ,
  \4502(2311)  = ~\4500(2286)  | ~\4497(1595) ,
  \4396(2353)  = ~\4394(2342)  | ~\4391(1547) ,
  \573(2157)  = ~\1263(2111) ,
  \3350(1331)  = \3343(1004)  & \3332(1163) ,
  \702(2228)  = \[89] ,
  \2253(786)  = \2226(209)  & (\2215(402)  & \200(85) ),
  \4504(2324)  = ~\4503(2288)  | ~\4502(2311) ,
  \749(2083)  = \2454(385)  & (\2418(193)  & \3793(2065) ),
  \2614(1327)  = ~\2611(1159) ,
  \3193(641)  = \3181(205)  & \83(31) ,
  \2994(394)  = \2948(282)  & \3547(201) ,
  \4456(2361)  = ~\4455(2344)  | ~\4454(2352) ,
  \5204(1393)  = ~\5202(1253)  | ~\5199(1089) ,
  \4075(817)  = \4049(178)  & (\4037(373)  & \116(46) ),
  \4191(1602)  = \1152(1452) ,
  \2808(1318)  = ~\2939(1144) ,
  \2694(392)  = \2643(311)  & \3547(201) ,
  \2876(683)  = \2847(656)  & \2838(398) ,
  \850(217)  = \[15] ,
  \4724(1142)  = \1749(988) ,
  \1758(1420)  = ~\1757(1141)  | ~\1756(1316) ,
  \788(2075)  = \2512(379)  & (\2488(381)  & \3851(2063) ),
  \949(852)  = \1688(663) ,
  \583(2150)  = ~\1944(2104) ,
  \5385(1885)  = ~\5383(1689)  | ~\5376(1808) ,
  \3853(1356)  = ~\3852(1190) ,
  \4967(2301)  = ~\4965(1655)  | ~\4958(2290) ,
  \2668(710)  = \2642(555)  & (\3551(199)  & \400(137) ),
  \822(1933)  = \[55] ,
  \5129(1041)  = \3137(914) ,
  \2930(872)  = \490(145)  | (\2929(749)  | \2927(510) ),
  \2686(670)  = \2630(563)  & \3549(200) ,
  \5311(976)  = ~\5307(862) ,
  \2872(682)  = \2847(656)  & \2838(398) ,
  \2757(770)  = \2741(493)  & \234(95) ,
  \3313(779)  = ~\3310(595) ,
  \5292(1543)  = ~\5286(1431) ,
  \4751(1485)  = \1794(1406) ,
  \3400(889)  = \3399(703)  | \3398(445) ,
  \3513(1216)  = \3492(726)  & (\3433(918)  & \3428(1036) ),
  \3530(1929)  = ~\3529(1767)  & ~\3528(1861) ,
  \3292(531)  = \3256(301)  & \3555(332) ,
  \3369(582)  = ~\3366(343) ,
  \4628(1063)  = \3161(926) ,
  \2807(1313)  = ~\2942(1137) ,
  \4861(2349)  = ~\4859(1384)  | ~\4852(2328) ,
  \4243(1690)  = ~\4239(1520) ,
  \1301(1000)  = \2798(948)  & \457(142) ,
  \4958(2290)  = ~\4957(2216)  | ~\4956(2267) ,
  \2684(390)  = \2627(322)  & \3547(201) ,
  \799(2080)  = \2512(379)  & (\2476(191)  & \3791(2067) ),
  \802(2183)  = \[81] ,
  \2669(903)  = \2668(710)  | \2666(458) ,
  \3547(201)  = ~\3546(165) ,
  \4906(2302)  = ~\4900(2281) ,
  \2907(764)  = \2889(526)  & \2370(326) ,
  \623(2152)  = \[58] ,
  \5395(1856)  = ~\5393(1677)  | ~\5386(1461) ,
  \759(2085)  = \2454(385)  & (\2418(193)  & \3791(2067) ),
  \1995(993)  = \3161(926)  & \479(144) ,
  \4747(1494)  = ~\4743(1415) ,
  \4385(1695)  = ~\4381(1529) ,
  \3230(868)  = \3229(692)  | \3228(424) ,
  \3365(583)  = ~\3362(344) ,
  \697(2175)  = \2351(616)  | (\2350(800)  | (\2349(2092)  | \2347(2088) )),
  \4762(1454)  = ~\4756(1363) ,
  \3789(807)  = \3757(181)  & (\3745(376)  & \128(56) ),
  \5364(772)  = ~\5362(586)  | ~\5359(338) ,
  \811(2219)  = \4096(2167)  & \4113(1859) ,
  \939(853)  = \1688(663) ,
  \2626(1335)  = ~\2623(1167) ,
  \4236(1173)  = \1071(1014) ,
  \1590(2201)  = \1564(404)  & (\1528(215)  & \4026(2185) ),
  \4212(1694)  = \1177(1524)  | (\1176(1558)  | \1064(996) ),
  \1920(1789)  = ~\4747(1494)  | ~\4740(1661) ,
  \3004(859)  = \523(148)  | (\3003(675)  | \3001(395) ),
  \1152(1452)  = ~\1151(1195)  | ~\1150(1360) ,
  \1621(405)  = ~\1609(214) ,
  \3942(1909)  = \3921(1816)  & (\3862(1566)  & \3857(1450) ),
  \4513(2332)  = ~\4511(1729)  | ~\4504(2324) ,
  \5043(1365)  = ~\5039(1199) ,
  \5118(1046)  = \3139(917) ,
  \748(2086)  = \2454(385)  & (\2430(383)  & \3851(2063) ),
  \4722(1143)  = ~\4716(989) ,
  \4592(2323)  = ~\4591(2287)  | ~\4590(2310) ,
  \838(2064)  = \[56] ,
  \5382(1888)  = ~\5376(1808) ,
  \2189(2437)  = ~\2188(2433) ,
  \752(2189)  = \[75] ,
  \4470(1193)  = ~\4464(1032) ,
  \5117(735)  = ~\5115(524)  | ~\5108(300) ,
  \792(2188)  = \[79] ,
  \4228(1015)  = ~\2788(945)  & ~\422(139) ,
  \830(2182)  = \[95] ,
  \4462(2374)  = ~\4456(2361) ,
  \1099(1188)  = ~\4163(463)  | ~\4156(1094) ,
  \3957(1389)  = \3941(1257)  & (\3910(1088)  & \3897(935) ),
  \2741(493)  = ~\2734(276) ,
  \4852(2328)  = ~\4851(2304)  | ~\4850(2319) ,
  \620(1800)  = \1166(1522)  & \1185(1721) ,
  \617(1849)  = \1843(1630)  & \1863(1675) ,
  \4590(2310)  = ~\4588(2285)  | ~\4585(1594) ,
  \998(2163)  = \3538(2117) ,
  \5107(729)  = ~\5105(512)  | ~\5098(290) ,
  \5012(1364)  = ~\5006(1198) ,
  \4636(1060)  = \3155(924) ,
  \2602(668)  = \2552(579)  & \3549(200) ,
  \4234(1174)  = ~\4228(1015) ,
  \784(2077)  = \3696(378)  & (\3660(190)  & \4024(2068) ),
  \3201(842)  = \3187(397)  & \34(12) ,
  \4870(1140)  = \2001(987) ,
  \4220(1693)  = ~\1178(1559)  & ~\1064(996) ,
  \762(2184)  = \[77] ,
  \4658(1051)  = ~\4652(920) ,
  \700(2176)  = \2357(617)  | (\2356(803)  | (\2355(2091)  | \2353(2089) )),
  \5404(1397)  = ~\5402(1271)  | ~\5399(946) ,
  \4454(2352)  = ~\4452(2343)  | ~\4449(1546) ,
  \665(2174)  = \1680(615)  | (\1679(801)  | (\1678(2099)  | \1676(2095) )),
  \2712(1349)  = ~\2709(1183) ,
  \1698(358)  = \137(63) ,
  \794(2079)  = \2512(379)  & (\2476(191)  & \3792(2066) ),
  \1982(1150)  = ~\4770(434)  | ~\4767(1064) ,
  \5239(1374)  = ~\5215(1233)  | ~\5214(1220) ,
  \1198(1778)  = ~\4194(662)  | ~\4191(1602) ,
  \2187(2423)  = ~\5005(1491)  | ~\4998(2416) ,
  \694(2172)  = \2345(613)  | (\2344(795)  | (\2343(2093)  | \2341(2032) )),
  \674(2171)  = \2254(606)  | (\2253(786)  | (\2252(2094)  | \2250(2090) )),
  \3643(634)  = \3616(182)  & \97(37) ,
  \3327(766)  = \3305(476)  & \2382(327) ,
  \4735(1498)  = \1767(1417) ,
  \590(1806)  = \1458(1719)  & \1437(1530) ,
  \604(223)  = \[9] ,
  \2357(617)  = \2304(208)  & (\2281(210)  & \146(67) ),
  \2188(2433)  = ~\2187(2423)  | ~\2186(2430) ,
  \793(2076)  = \2512(379)  & (\2488(381)  & \3850(2069) ),
  \4898(2261)  = ~\4896(2217)  | ~\4893(1500) ,
  \3637(635)  = \3616(182)  & \97(37) ,
  \2838(398)  = ~\2828(206) ,
  \2184(2411)  = ~\4995(1492)  | ~\4988(2391) ,
  \693(2179)  = \[73] ,
  \4443(1697)  = ~\4439(1532) ,
  \627(1764)  = \2117(1504)  | (\2116(1152)  | (\2115(1229)  | \3167(931) )),
  \744(2081)  = \3594(384)  & (\3558(192)  & \4024(2068) ),
  \1079(1172)  = ~\4147(451)  | ~\4140(1102) ,
  \4562(1965)  = ~\4561(1911)  | ~\4560(1837) ,
  \1071(1014)  = \2788(945)  & \422(139) ,
  \4510(2335)  = ~\4504(2324) ,
  \2183(2417)  = ~\4994(2410)  | ~\4991(1414) ,
  \858(647)  = \2500(189)  & (\2476(191)  & \61(21) ),
  \2195(2429)  = \2185(2424)  & \2174(161) ,
  \2827(620)  = \1701(355) ,
  \3389(998)  = ~\3388(882) ,
  \5105(512)  = ~\5101(289) ,
  \2198(2449)  = ~\2197(2447)  | ~\2196(2443) ,
  \4011(811)  = \3991(179)  & (\3979(374)  & \122(52) ),
  \783(2074)  = \3696(378)  & (\3672(380)  & \4082(2071) ),
  \5132(1035)  = ~\5126(912) ,
  \4348(1016)  = ~\2788(945)  & ~\422(139) ,
  \4377(2213)  = ~\4375(1725)  | ~\4368(2156) ,
  \4512(2346)  = ~\4510(2335)  | ~\4507(1571) ,
  \5259(1931)  = ~\5255(1860) ,
  \1685(802)  = \1633(212)  & (\1621(405)  & \149(68) ),
  \2580(706)  = \2556(580)  & (\3551(199)  & \422(139) ),
  \3545(2169)  = ~\3543(2120) ,
  \2924(748)  = \2893(519)  & \3556(324) ,
  \4239(1520)  = \1052(1426) ,
  \753(2087)  = \2454(385)  & (\2430(383)  & \3850(2069) ),
  \3841(806)  = \3815(180)  & (\3803(375)  & \129(57) ),
  \757(2190)  = \[76] ,
  \2185(2424)  = ~\2184(2411)  | ~\2183(2417) ,
  \4600(2347)  = ~\4598(2334)  | ~\4595(1574) ,
  \4588(2285)  = ~\4582(2265) ,
  \616(1763)  = \1847(1509)  | (\1846(1147)  | (\1845(1226)  | \3167(931) )),
  \2920(747)  = \2885(534)  & \3556(324) ,
  \3039(552)  = ~\3036(314) ,
  \3035(554)  = ~\3032(315) ,
  \743(2082)  = \3594(384)  & (\3570(382)  & \4082(2071) ),
  \2186(2430)  = ~\5004(2422)  | ~\5001(1413) ,
  \4601(2333)  = ~\4599(1730)  | ~\4592(2323) ,
  \754(2084)  = \2454(385)  & (\2418(193)  & \3792(2066) ),
  \1679(801)  = \1633(212)  & (\1621(405)  & \155(70) ),
  \5115(524)  = ~\5111(296) ,
  \3849(2024)  = \3841(806)  | (\3840(1935)  | \3839(1291) ),
  \5275(1353)  = ~\5271(1187) ,
  \2197(2447)  = ~\5081(2444)  | ~\5074(2414) ,
  \3537(2019)  = ~\5251(1922)  | ~\5244(1966) ,
  \4282(444)  = ~\4276(243) ,
  \3118(715)  = \3099(496)  & \369(131) ,
  \2476(191)  = \4089(173) ,
  \4842(2282)  = ~\4841(2208)  | ~\4840(2262) ,
  \797(2191)  = \[80] ,
  \1088(1169)  = ~\4155(448)  | ~\4148(1098) ,
  \662(2173)  = \1674(614)  | (\1673(794)  | (\1672(2100)  | \1670(2034) )),
  \3904(742)  = ~\5346(557)  | ~\5343(313) ,
  \2674(707)  = \2650(549)  & (\3551(199)  & \411(138) ),
  \4644(1055)  = \3151(923) ,
  \661(2178)  = \[72] ,
  \4787(1052)  = ~\4783(921) ,
  \4414(1902)  = ~\4412(1343)  | ~\4409(1807) ,
  \5346(557)  = ~\5340(318) ,
  \1829(1037)  = ~\3137(914) ,
  \3594(384)  = ~\3582(194) ,
  \5339(536)  = ~\5335(303) ,
  \5384(1947)  = ~\5382(1888)  | ~\5379(1518) ,
  \2622(1339)  = ~\2619(1171) ,
  \3120(717)  = \3099(496)  & \361(129) ,
  \4473(1910)  = ~\4471(1828)  | ~\4464(1032) ,
  \593(733)  = \[34] ,
  \4850(2319)  = ~\4848(2303)  | ~\4845(1516) ,
  \4449(1546)  = \1278(1433) ,
  \3386(439)  = \3358(350)  & (\457(142)  & \2393(328) ),
  \4171(460)  = ~\4167(251) ,
  \2590(386)  = \2533(351)  & \3547(201) ,
  \1218(1821)  = ~\4235(1691)  | ~\4228(1015) ,
  \4356(1901)  = ~\4354(1176)  | ~\4351(1805) ,
  \3871(1548)  = ~\3870(1434)  | ~\3869(1447) ,
  \4439(1532)  = \1307(1427) ,
  \4459(1538)  = \1289(1428) ,
  \2971(482)  = ~\2968(266) ,
  \4775(1056)  = \3151(923) ,
  \4807(1059)  = \3155(924) ,
  \3124(721)  = \3099(496)  & \341(125) ,
  \626(1752)  = \[47] ,
  \571(2052)  = ~\1273(2005) ,
  \1730(1422)  = ~\1729(1146)  | ~\1728(1320) ,
  \2196(2443)  = ~\5080(2420)  | ~\5077(2441) ,
  \4188(363)  = \4(1) ,
  \3964(2042)  = ~\5421(1942)  | ~\5414(2018) ,
  \640(2170)  = \1580(605)  | (\1579(787)  | (\1578(2101)  | \1576(2097) )),
  \1247(1822)  = ~\4267(1736)  | ~\4260(1727) ,
  \4464(1032)  = ~\2767(936)  & ~\374(134) ,
  \4179(455)  = ~\4175(248) ,
  \1430(1451)  = ~\1429(1358)  | ~\1428(1192) ,
  \2194(2439)  = \2179(207)  & \2189(2437) ,
  \4435(2212)  = ~\4433(1724)  | ~\4426(2155) ,
  \2488(381)  = ~\2476(191) ,
  \5421(1942)  = ~\5417(1877) ,
  \4517(1550)  = \1332(1435) ,
  \1428(1192)  = ~\4346(468)  | ~\4343(1084) ,
  \3031(562)  = ~\3028(321) ,
  \4374(2211)  = ~\4368(2156) ,
  \4767(1064)  = \3161(926) ,
  \3582(194)  = \4087(171) ,
  \4028(2234)  = \4023(818)  | (\4022(2136)  | \4021(1401) ),
  \3648(2192)  = \3632(377)  & \3962(2154) ,
  \2568(700)  = \2540(592)  & (\3551(199)  & \457(142) ),
  \3121(472)  = \3092(279)  & \366(130) ,
  \1897(1883)  = ~\1896(1796)  | ~\1895(1681) ,
  \2982(413)  = \2960(273)  & (\523(148)  & \3553(198) );
endmodule

