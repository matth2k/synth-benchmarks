module s15850 (
  CK,
  g100,
  g101,
  g102,
  g103,
  g104,
  g109,
  g1170,
  g1173,
  g1176,
  g1179,
  g1182,
  g1185,
  g1188,
  g1191,
  g1194,
  g1197,
  g1200,
  g1203,
  g1696,
  g1700,
  g1712,
  g18,
  g1960,
  g1961,
  g23,
  g27,
  g28,
  g29,
  g30,
  g31,
  g41,
  g42,
  g43,
  g44,
  g45,
  g46,
  g47,
  g48,
  g741,
  g742,
  g743,
  g744,
  g750,
  g82,
  g83,
  g84,
  g85,
  g86,
  g87,
  g872,
  g873,
  g877,
  g88,
  g881,
  g886,
  g889,
  g89,
  g892,
  g895,
  g898,
  g90,
  g901,
  g904,
  g907,
  g91,
  g910,
  g913,
  g916,
  g919,
  g92,
  g922,
  g925,
  g93,
  g94,
  g95,
  g96,
  g99,
  g7744,
  g6926,
  g8562,
  g6282,
  g4888,
  g6264,
  g4193,
  g6284,
  g2601,
  g2610,
  g2602,
  g2607,
  g4194,
  g6280,
  g8982,
  g4176,
  g11163,
  g2604,
  g2609,
  g4215,
  g10465,
  g4198,
  g4201,
  g10459,
  g8328,
  g10461,
  g8984,
  g4211,
  g6920,
  g8561,
  g6270,
  g8979,
  g10457,
  g4210,
  g8313,
  g4214,
  g6279,
  g4887,
  g6257,
  g8323,
  g8318,
  g4180,
  g4192,
  g8349,
  g8335,
  g4195,
  g4202,
  g4207,
  g3069,
  g6259,
  g8977,
  g4203,
  g6281,
  g6254,
  g6258,
  g4178,
  g6268,
  g4191,
  g4177,
  g4205,
  g6267,
  g10377,
  g2648,
  g6942,
  g8564,
  g2355,
  g4171,
  g6932,
  g8563,
  g10463,
  g4208,
  g8340,
  g6260,
  g6277,
  g6255,
  g11489,
  g4172,
  g3007,
  g10455,
  g4173,
  g5816,
  g8271,
  g6275,
  g6265,
  g4209,
  g6283,
  g6949,
  g8565,
  g8316,
  g6278,
  g8352,
  g9451,
  g9961,
  g4216,
  g6276,
  g6263,
  g8985,
  g11206,
  g2986,
  g6285,
  g6842,
  g4179,
  g4204,
  g10801,
  g8986,
  g6273,
  g8347,
  g6262,
  g5101,
  g8061,
  g4212,
  g10379,
  g5659,
  g6253,
  g4206,
  g6271,
  g5105,
  g8062,
  g8331,
  g4196,
  g6266,
  g6272,
  g6955,
  g8566,
  g5658,
  g6261,
  g4181,
  g4213,
  g8980,
  g4200,
  g3327,
  g1957,
  g4174,
  g6274,
  g8978,
  g8981,
  g2603,
  g2608,
  g8976,
  g2606,
  g2612,
  g2605,
  g2611,
  g6269,
  g10628,
  g4175,
  g6256,
  g8983,
  g4197,
  g4199
);
  input CK;
  wire CK;
  input g100;
  wire g100;
  input g101;
  wire g101;
  input g102;
  wire g102;
  input g103;
  wire g103;
  input g104;
  wire g104;
  input g109;
  wire g109;
  input g1170;
  wire g1170;
  input g1173;
  wire g1173;
  input g1176;
  wire g1176;
  input g1179;
  wire g1179;
  input g1182;
  wire g1182;
  input g1185;
  wire g1185;
  input g1188;
  wire g1188;
  input g1191;
  wire g1191;
  input g1194;
  wire g1194;
  input g1197;
  wire g1197;
  input g1200;
  wire g1200;
  input g1203;
  wire g1203;
  input g1696;
  wire g1696;
  input g1700;
  wire g1700;
  input g1712;
  wire g1712;
  input g18;
  wire g18;
  input g1960;
  wire g1960;
  input g1961;
  wire g1961;
  input g23;
  wire g23;
  input g27;
  wire g27;
  input g28;
  wire g28;
  input g29;
  wire g29;
  input g30;
  wire g30;
  input g31;
  wire g31;
  input g41;
  wire g41;
  input g42;
  wire g42;
  input g43;
  wire g43;
  input g44;
  wire g44;
  input g45;
  wire g45;
  input g46;
  wire g46;
  input g47;
  wire g47;
  input g48;
  wire g48;
  input g741;
  wire g741;
  input g742;
  wire g742;
  input g743;
  wire g743;
  input g744;
  wire g744;
  input g750;
  wire g750;
  input g82;
  wire g82;
  input g83;
  wire g83;
  input g84;
  wire g84;
  input g85;
  wire g85;
  input g86;
  wire g86;
  input g87;
  wire g87;
  input g872;
  wire g872;
  input g873;
  wire g873;
  input g877;
  wire g877;
  input g88;
  wire g88;
  input g881;
  wire g881;
  input g886;
  wire g886;
  input g889;
  wire g889;
  input g89;
  wire g89;
  input g892;
  wire g892;
  input g895;
  wire g895;
  input g898;
  wire g898;
  input g90;
  wire g90;
  input g901;
  wire g901;
  input g904;
  wire g904;
  input g907;
  wire g907;
  input g91;
  wire g91;
  input g910;
  wire g910;
  input g913;
  wire g913;
  input g916;
  wire g916;
  input g919;
  wire g919;
  input g92;
  wire g92;
  input g922;
  wire g922;
  input g925;
  wire g925;
  input g93;
  wire g93;
  input g94;
  wire g94;
  input g95;
  wire g95;
  input g96;
  wire g96;
  input g99;
  wire g99;
  output g7744;
  wire g7744;
  output g6926;
  wire g6926;
  output g8562;
  wire g8562;
  output g6282;
  wire g6282;
  output g4888;
  wire g4888;
  output g6264;
  wire g6264;
  output g4193;
  wire g4193;
  output g6284;
  wire g6284;
  output g2601;
  wire g2601;
  output g2610;
  wire g2610;
  output g2602;
  wire g2602;
  output g2607;
  wire g2607;
  output g4194;
  wire g4194;
  output g6280;
  wire g6280;
  output g8982;
  wire g8982;
  output g4176;
  wire g4176;
  output g11163;
  wire g11163;
  output g2604;
  wire g2604;
  output g2609;
  wire g2609;
  output g4215;
  wire g4215;
  output g10465;
  wire g10465;
  output g4198;
  wire g4198;
  output g4201;
  wire g4201;
  output g10459;
  wire g10459;
  output g8328;
  wire g8328;
  output g10461;
  wire g10461;
  output g8984;
  wire g8984;
  output g4211;
  wire g4211;
  output g6920;
  wire g6920;
  output g8561;
  wire g8561;
  output g6270;
  wire g6270;
  output g8979;
  wire g8979;
  output g10457;
  wire g10457;
  output g4210;
  wire g4210;
  output g8313;
  wire g8313;
  output g4214;
  wire g4214;
  output g6279;
  wire g6279;
  output g4887;
  wire g4887;
  output g6257;
  wire g6257;
  output g8323;
  wire g8323;
  output g8318;
  wire g8318;
  output g4180;
  wire g4180;
  output g4192;
  wire g4192;
  output g8349;
  wire g8349;
  output g8335;
  wire g8335;
  output g4195;
  wire g4195;
  output g4202;
  wire g4202;
  output g4207;
  wire g4207;
  output g3069;
  wire g3069;
  output g6259;
  wire g6259;
  output g8977;
  wire g8977;
  output g4203;
  wire g4203;
  output g6281;
  wire g6281;
  output g6254;
  wire g6254;
  output g6258;
  wire g6258;
  output g4178;
  wire g4178;
  output g6268;
  wire g6268;
  output g4191;
  wire g4191;
  output g4177;
  wire g4177;
  output g4205;
  wire g4205;
  output g6267;
  wire g6267;
  output g10377;
  wire g10377;
  output g2648;
  wire g2648;
  output g6942;
  wire g6942;
  output g8564;
  wire g8564;
  output g2355;
  wire g2355;
  output g4171;
  wire g4171;
  output g6932;
  wire g6932;
  output g8563;
  wire g8563;
  output g10463;
  wire g10463;
  output g4208;
  wire g4208;
  output g8340;
  wire g8340;
  output g6260;
  wire g6260;
  output g6277;
  wire g6277;
  output g6255;
  wire g6255;
  output g11489;
  wire g11489;
  output g4172;
  wire g4172;
  output g3007;
  wire g3007;
  output g10455;
  wire g10455;
  output g4173;
  wire g4173;
  output g5816;
  wire g5816;
  output g8271;
  wire g8271;
  output g6275;
  wire g6275;
  output g6265;
  wire g6265;
  output g4209;
  wire g4209;
  output g6283;
  wire g6283;
  output g6949;
  wire g6949;
  output g8565;
  wire g8565;
  output g8316;
  wire g8316;
  output g6278;
  wire g6278;
  output g8352;
  wire g8352;
  output g9451;
  wire g9451;
  output g9961;
  wire g9961;
  output g4216;
  wire g4216;
  output g6276;
  wire g6276;
  output g6263;
  wire g6263;
  output g8985;
  wire g8985;
  output g11206;
  wire g11206;
  output g2986;
  wire g2986;
  output g6285;
  wire g6285;
  output g6842;
  wire g6842;
  output g4179;
  wire g4179;
  output g4204;
  wire g4204;
  output g10801;
  wire g10801;
  output g8986;
  wire g8986;
  output g6273;
  wire g6273;
  output g8347;
  wire g8347;
  output g6262;
  wire g6262;
  output g5101;
  wire g5101;
  output g8061;
  wire g8061;
  output g4212;
  wire g4212;
  output g10379;
  wire g10379;
  output g5659;
  wire g5659;
  output g6253;
  wire g6253;
  output g4206;
  wire g4206;
  output g6271;
  wire g6271;
  output g5105;
  wire g5105;
  output g8062;
  wire g8062;
  output g8331;
  wire g8331;
  output g4196;
  wire g4196;
  output g6266;
  wire g6266;
  output g6272;
  wire g6272;
  output g6955;
  wire g6955;
  output g8566;
  wire g8566;
  output g5658;
  wire g5658;
  output g6261;
  wire g6261;
  output g4181;
  wire g4181;
  output g4213;
  wire g4213;
  output g8980;
  wire g8980;
  output g4200;
  wire g4200;
  output g3327;
  wire g3327;
  output g1957;
  wire g1957;
  output g4174;
  wire g4174;
  output g6274;
  wire g6274;
  output g8978;
  wire g8978;
  output g8981;
  wire g8981;
  output g2603;
  wire g2603;
  output g2608;
  wire g2608;
  output g8976;
  wire g8976;
  output g2606;
  wire g2606;
  output g2612;
  wire g2612;
  output g2605;
  wire g2605;
  output g2611;
  wire g2611;
  output g6269;
  wire g6269;
  output g10628;
  wire g10628;
  output g4175;
  wire g4175;
  output g6256;
  wire g6256;
  output g8983;
  wire g8983;
  output g4197;
  wire g4197;
  output g4199;
  wire g4199;
  wire __0__;
  wire __1__;
  wire __2__;
  wire __3__;
  wire __4__;
  wire __5__;
  wire __6__;
  wire __7__;
  wire __8__;
  wire __9__;
  wire __10__;
  wire __11__;
  wire __12__;
  wire __13__;
  wire __14__;
  wire __15__;
  wire __16__;
  wire __17__;
  wire __18__;
  wire __19__;
  wire __20__;
  wire __21__;
  wire __22__;
  wire __23__;
  wire __24__;
  wire __25__;
  wire __26__;
  wire __27__;
  wire __28__;
  wire __29__;
  wire __30__;
  wire __31__;
  wire __32__;
  wire __33__;
  wire __34__;
  wire __35__;
  wire __36__;
  wire __37__;
  wire __38__;
  wire __39__;
  wire __40__;
  wire __41__;
  wire __42__;
  wire __43__;
  wire __44__;
  wire __45__;
  wire __46__;
  wire __47__;
  wire __48__;
  wire __49__;
  wire __50__;
  wire __51__;
  wire __52__;
  wire __53__;
  wire __54__;
  wire __55__;
  wire __56__;
  wire __57__;
  wire __58__;
  wire __59__;
  wire __60__;
  wire __61__;
  wire __62__;
  wire __63__;
  wire __64__;
  wire __65__;
  wire __66__;
  wire __67__;
  wire __68__;
  wire __69__;
  wire __70__;
  wire __71__;
  wire __72__;
  wire __73__;
  wire __74__;
  wire __75__;
  wire __76__;
  wire __77__;
  wire __78__;
  wire __79__;
  wire __80__;
  wire __81__;
  wire __82__;
  wire __83__;
  wire __84__;
  wire __85__;
  wire __86__;
  wire __87__;
  wire __88__;
  wire __89__;
  wire __90__;
  wire __91__;
  wire __92__;
  wire __93__;
  wire __94__;
  wire __95__;
  wire __96__;
  wire __97__;
  wire __98__;
  wire __99__;
  wire __100__;
  wire __101__;
  wire __102__;
  wire __103__;
  wire __104__;
  wire __105__;
  wire __106__;
  wire __107__;
  wire __108__;
  wire __109__;
  wire __110__;
  wire __111__;
  wire __112__;
  wire __113__;
  wire __114__;
  wire __115__;
  wire __116__;
  wire __117__;
  wire __118__;
  wire __119__;
  wire __120__;
  wire __121__;
  wire __122__;
  wire __123__;
  wire __124__;
  wire __125__;
  wire __126__;
  wire __127__;
  wire __128__;
  wire __129__;
  wire __130__;
  wire __131__;
  wire __132__;
  wire __133__;
  wire __134__;
  wire __135__;
  wire __136__;
  wire __137__;
  wire __138__;
  wire __139__;
  wire __140__;
  wire __141__;
  wire __142__;
  wire __143__;
  wire __144__;
  wire __145__;
  wire __146__;
  wire __147__;
  wire __148__;
  wire __149__;
  wire __150__;
  wire __151__;
  wire __152__;
  wire __153__;
  wire __154__;
  wire __155__;
  wire __156__;
  wire __157__;
  wire __158__;
  wire __159__;
  wire __160__;
  wire __161__;
  wire __162__;
  wire __163__;
  wire __164__;
  wire __165__;
  wire __166__;
  wire __167__;
  wire __168__;
  wire __169__;
  wire __170__;
  wire __171__;
  wire __172__;
  wire __173__;
  wire __174__;
  wire __175__;
  wire __176__;
  wire __177__;
  wire __178__;
  wire __179__;
  wire __180__;
  wire __181__;
  wire __182__;
  wire __183__;
  wire __184__;
  wire __185__;
  wire __186__;
  wire __187__;
  wire __188__;
  wire __189__;
  wire __190__;
  wire __191__;
  wire __192__;
  wire __193__;
  wire __194__;
  wire __195__;
  wire __196__;
  wire __197__;
  wire __198__;
  wire __199__;
  wire __200__;
  wire __201__;
  wire __202__;
  wire __203__;
  wire __204__;
  wire __205__;
  wire __206__;
  wire __207__;
  wire __208__;
  wire __209__;
  wire __210__;
  wire __211__;
  wire __212__;
  wire __213__;
  wire __214__;
  wire __215__;
  wire __216__;
  wire __217__;
  wire __218__;
  wire __219__;
  wire __220__;
  wire __221__;
  wire __222__;
  wire __223__;
  wire __224__;
  wire __225__;
  wire __226__;
  wire __227__;
  wire __228__;
  wire __229__;
  wire __230__;
  wire __231__;
  wire __232__;
  wire __233__;
  wire __234__;
  wire __235__;
  wire __236__;
  wire __237__;
  wire __238__;
  wire __239__;
  wire __240__;
  wire __241__;
  wire __242__;
  wire __243__;
  wire __244__;
  wire __245__;
  wire __246__;
  wire __247__;
  wire __248__;
  wire __249__;
  wire __250__;
  wire __251__;
  wire __252__;
  wire __253__;
  wire __254__;
  wire __255__;
  wire __256__;
  wire __257__;
  wire __258__;
  wire __259__;
  wire __260__;
  wire __261__;
  wire __262__;
  wire __263__;
  wire __264__;
  wire __265__;
  wire __266__;
  wire __267__;
  wire __268__;
  wire __269__;
  wire __270__;
  wire __271__;
  wire __272__;
  wire __273__;
  wire __274__;
  wire __275__;
  wire __276__;
  wire __277__;
  wire __278__;
  wire __279__;
  wire __280__;
  wire __281__;
  wire __282__;
  wire __283__;
  wire __284__;
  wire __285__;
  wire __286__;
  wire __287__;
  wire __288__;
  wire __289__;
  wire __290__;
  wire __291__;
  wire __292__;
  wire __293__;
  wire __294__;
  wire __295__;
  wire __296__;
  wire __297__;
  wire __298__;
  wire __299__;
  wire __300__;
  wire __301__;
  wire __302__;
  wire __303__;
  wire __304__;
  wire __305__;
  wire __306__;
  wire __307__;
  wire __308__;
  wire __309__;
  wire __310__;
  wire __311__;
  wire __312__;
  wire __313__;
  wire __314__;
  wire __315__;
  wire __316__;
  wire __317__;
  wire __318__;
  wire __319__;
  wire __320__;
  wire __321__;
  wire __322__;
  wire __323__;
  wire __324__;
  wire __325__;
  wire __326__;
  wire __327__;
  wire __328__;
  wire __329__;
  wire __330__;
  wire __331__;
  wire __332__;
  wire __333__;
  wire __334__;
  wire __335__;
  wire __336__;
  wire __337__;
  wire __338__;
  wire __339__;
  wire __340__;
  wire __341__;
  wire __342__;
  wire __343__;
  wire __344__;
  wire __345__;
  wire __346__;
  wire __347__;
  wire __348__;
  wire __349__;
  wire __350__;
  wire __351__;
  wire __352__;
  wire __353__;
  wire __354__;
  wire __355__;
  wire __356__;
  wire __357__;
  wire __358__;
  wire __359__;
  wire __360__;
  wire __361__;
  wire __362__;
  wire __363__;
  wire __364__;
  wire __365__;
  wire __366__;
  wire __367__;
  wire __368__;
  wire __369__;
  wire __370__;
  wire __371__;
  wire __372__;
  wire __373__;
  wire __374__;
  wire __375__;
  wire __376__;
  wire __377__;
  wire __378__;
  wire __379__;
  wire __380__;
  wire __381__;
  wire __382__;
  wire __383__;
  wire __384__;
  wire __385__;
  wire __386__;
  wire __387__;
  wire __388__;
  wire __389__;
  wire __390__;
  wire __391__;
  wire __392__;
  wire __393__;
  wire __394__;
  wire __395__;
  wire __396__;
  wire __397__;
  wire __398__;
  wire __399__;
  wire __400__;
  wire __401__;
  wire __402__;
  wire __403__;
  wire __404__;
  wire __405__;
  wire __406__;
  wire __407__;
  wire __408__;
  wire __409__;
  wire __410__;
  wire __411__;
  wire __412__;
  wire __413__;
  wire __414__;
  wire __415__;
  wire __416__;
  wire __417__;
  wire __418__;
  wire __419__;
  wire __420__;
  wire __421__;
  wire __422__;
  wire __423__;
  wire __424__;
  wire __425__;
  wire __426__;
  wire __427__;
  wire __428__;
  wire __429__;
  wire __430__;
  wire __431__;
  wire __432__;
  wire __433__;
  wire __434__;
  wire __435__;
  wire __436__;
  wire __437__;
  wire __438__;
  wire __439__;
  wire __440__;
  wire __441__;
  wire __442__;
  wire __443__;
  wire __444__;
  wire __445__;
  wire __446__;
  wire __447__;
  wire __448__;
  wire __449__;
  wire __450__;
  wire __451__;
  wire __452__;
  wire __453__;
  wire __454__;
  wire __455__;
  wire __456__;
  wire __457__;
  wire __458__;
  wire __459__;
  wire __460__;
  wire __461__;
  wire __462__;
  wire __463__;
  wire __464__;
  wire __465__;
  wire __466__;
  wire __467__;
  wire __468__;
  wire __469__;
  wire __470__;
  wire __471__;
  wire __472__;
  wire __473__;
  wire __474__;
  wire __475__;
  wire __476__;
  wire __477__;
  wire __478__;
  wire __479__;
  wire __480__;
  wire __481__;
  wire __482__;
  wire __483__;
  wire __484__;
  wire __485__;
  wire __486__;
  wire __487__;
  wire __488__;
  wire __489__;
  wire __490__;
  wire __491__;
  wire __492__;
  wire __493__;
  wire __494__;
  wire __495__;
  wire __496__;
  wire __497__;
  wire __498__;
  wire __499__;
  wire __500__;
  wire __501__;
  wire __502__;
  wire __503__;
  wire __504__;
  wire __505__;
  wire __506__;
  wire __508__;
  wire __509__;
  wire __511__;
  wire __512__;
  wire __513__;
  wire __514__;
  wire __515__;
  wire __516__;
  wire __517__;
  wire __518__;
  wire __519__;
  wire __520__;
  wire __521__;
  wire __522__;
  wire __523__;
  wire __524__;
  wire __525__;
  wire __526__;
  wire __527__;
  wire __528__;
  wire __529__;
  wire __530__;
  wire __531__;
  wire __532__;
  wire __533__;
  wire __534__;
  wire __535__;
  wire __536__;
  wire __537__;
  wire __538__;
  wire __539__;
  wire __540__;
  wire __541__;
  wire __542__;
  wire __543__;
  wire __544__;
  wire __545__;
  wire __546__;
  wire __547__;
  wire __548__;
  wire __549__;
  wire __550__;
  wire __551__;
  wire __552__;
  wire __553__;
  wire __554__;
  wire __555__;
  wire __556__;
  wire __557__;
  wire __558__;
  wire __559__;
  wire __560__;
  wire __561__;
  wire __562__;
  wire __563__;
  wire __564__;
  wire __565__;
  wire __566__;
  wire __567__;
  wire __568__;
  wire __569__;
  wire __570__;
  wire __571__;
  wire __572__;
  wire __573__;
  wire __574__;
  wire __575__;
  wire __576__;
  wire __577__;
  wire __578__;
  wire __579__;
  wire __580__;
  wire __581__;
  wire __582__;
  wire __583__;
  wire __584__;
  wire __585__;
  wire __586__;
  wire __587__;
  wire __588__;
  wire __589__;
  wire __590__;
  wire __591__;
  wire __592__;
  wire __593__;
  wire __594__;
  wire __595__;
  wire __596__;
  wire __597__;
  wire __598__;
  wire __599__;
  wire __600__;
  wire __601__;
  wire __602__;
  wire __603__;
  wire __604__;
  wire __605__;
  wire __606__;
  wire __607__;
  wire __608__;
  wire __609__;
  wire __610__;
  wire __611__;
  wire __612__;
  wire __613__;
  wire __614__;
  wire __615__;
  wire __616__;
  wire __617__;
  wire __618__;
  wire __619__;
  wire __620__;
  wire __621__;
  wire __622__;
  wire __623__;
  wire __624__;
  wire __625__;
  wire __626__;
  wire __627__;
  wire __628__;
  wire __629__;
  wire __630__;
  wire __631__;
  wire __632__;
  wire __633__;
  wire __634__;
  wire __635__;
  wire __636__;
  wire __637__;
  wire __638__;
  wire __639__;
  wire __640__;
  wire __641__;
  wire __642__;
  wire __643__;
  wire __644__;
  wire __645__;
  wire __646__;
  wire __647__;
  wire __648__;
  wire __649__;
  wire __650__;
  wire __651__;
  wire __652__;
  wire __653__;
  wire __654__;
  wire __655__;
  wire __656__;
  wire __657__;
  wire __658__;
  wire __659__;
  wire __660__;
  wire __661__;
  wire __662__;
  wire __663__;
  wire __664__;
  wire __665__;
  wire __666__;
  wire __667__;
  wire __668__;
  wire __669__;
  wire __670__;
  wire __671__;
  wire __672__;
  wire __673__;
  wire __674__;
  wire __675__;
  wire __676__;
  wire __677__;
  wire __678__;
  wire __679__;
  wire __680__;
  wire __681__;
  wire __682__;
  wire __683__;
  wire __684__;
  wire __685__;
  wire __686__;
  wire __687__;
  wire __688__;
  wire __689__;
  wire __690__;
  wire __691__;
  wire __692__;
  wire __693__;
  wire __694__;
  wire __695__;
  wire __696__;
  wire __697__;
  wire __698__;
  wire __699__;
  wire __700__;
  wire __701__;
  wire __702__;
  wire __703__;
  wire __704__;
  wire __705__;
  wire __706__;
  wire __707__;
  wire __708__;
  wire __709__;
  wire __710__;
  wire __711__;
  wire __712__;
  wire __713__;
  wire __714__;
  wire __715__;
  wire __716__;
  wire __717__;
  wire __718__;
  wire __719__;
  wire __720__;
  wire __721__;
  wire __722__;
  wire __723__;
  wire __724__;
  wire __725__;
  wire __726__;
  wire __727__;
  wire __728__;
  wire __729__;
  wire __730__;
  wire __731__;
  wire __732__;
  wire __733__;
  wire __734__;
  wire __735__;
  wire __736__;
  wire __737__;
  wire __738__;
  wire __739__;
  wire __740__;
  wire __741__;
  wire __742__;
  wire __743__;
  wire __744__;
  wire __745__;
  wire __746__;
  wire __747__;
  wire __748__;
  wire __749__;
  wire __750__;
  wire __751__;
  wire __752__;
  wire __753__;
  wire __754__;
  wire __755__;
  wire __756__;
  wire __757__;
  wire __758__;
  wire __759__;
  wire __760__;
  wire __761__;
  wire __762__;
  wire __763__;
  wire __764__;
  wire __765__;
  wire __766__;
  wire __767__;
  wire __768__;
  wire __769__;
  wire __770__;
  wire __771__;
  wire __772__;
  wire __773__;
  wire __774__;
  wire __775__;
  wire __776__;
  wire __777__;
  wire __778__;
  wire __779__;
  wire __780__;
  wire __781__;
  wire __782__;
  wire __783__;
  wire __784__;
  wire __785__;
  wire __786__;
  wire __787__;
  wire __788__;
  wire __789__;
  wire __790__;
  wire __791__;
  wire __792__;
  wire __793__;
  wire __794__;
  wire __795__;
  wire __796__;
  wire __797__;
  wire __798__;
  wire __799__;
  wire __800__;
  wire __801__;
  wire __802__;
  wire __803__;
  wire __804__;
  wire __805__;
  wire __806__;
  wire __807__;
  wire __808__;
  wire __809__;
  wire __810__;
  wire __811__;
  wire __812__;
  wire __813__;
  wire __814__;
  wire __815__;
  wire __816__;
  wire __817__;
  wire __818__;
  wire __819__;
  wire __820__;
  wire __821__;
  wire __822__;
  wire __823__;
  wire __824__;
  wire __825__;
  wire __826__;
  wire __827__;
  wire __828__;
  wire __829__;
  wire __830__;
  wire __831__;
  wire __832__;
  wire __833__;
  wire __834__;
  wire __835__;
  wire __836__;
  wire __837__;
  wire __838__;
  wire __839__;
  wire __840__;
  wire __841__;
  wire __842__;
  wire __843__;
  wire __844__;
  wire __845__;
  wire __846__;
  wire __847__;
  wire __848__;
  wire __849__;
  wire __850__;
  wire __851__;
  wire __852__;
  wire __853__;
  wire __854__;
  wire __855__;
  wire __856__;
  wire __857__;
  wire __858__;
  wire __859__;
  wire __860__;
  wire __861__;
  wire __862__;
  wire __863__;
  wire __864__;
  wire __865__;
  wire __866__;
  wire __867__;
  wire __868__;
  wire __869__;
  wire __870__;
  wire __871__;
  wire __872__;
  wire __873__;
  wire __874__;
  wire __875__;
  wire __876__;
  wire __877__;
  wire __878__;
  wire __879__;
  wire __880__;
  wire __881__;
  wire __882__;
  wire __883__;
  wire __884__;
  wire __885__;
  wire __886__;
  wire __887__;
  wire __888__;
  wire __889__;
  wire __890__;
  wire __891__;
  wire __892__;
  wire __893__;
  wire __894__;
  wire __895__;
  wire __896__;
  wire __897__;
  wire __898__;
  wire __899__;
  wire __900__;
  wire __901__;
  wire __902__;
  wire __903__;
  wire __904__;
  wire __905__;
  wire __906__;
  wire __907__;
  wire __908__;
  wire __909__;
  wire __910__;
  wire __911__;
  wire __912__;
  wire __913__;
  wire __914__;
  wire __915__;
  wire __916__;
  wire __917__;
  wire __918__;
  wire __919__;
  wire __920__;
  wire __921__;
  wire __922__;
  wire __923__;
  wire __924__;
  wire __925__;
  wire __926__;
  wire __927__;
  wire __928__;
  wire __929__;
  wire __930__;
  wire __931__;
  wire __932__;
  wire __933__;
  wire __934__;
  wire __935__;
  wire __936__;
  wire __937__;
  wire __938__;
  wire __939__;
  wire __940__;
  wire __941__;
  wire __942__;
  wire __943__;
  wire __944__;
  wire __945__;
  wire __946__;
  wire __947__;
  wire __948__;
  wire __949__;
  wire __950__;
  wire __951__;
  wire __952__;
  wire __953__;
  wire __954__;
  wire __955__;
  wire __956__;
  wire __957__;
  wire __958__;
  wire __959__;
  wire __960__;
  wire __961__;
  wire __962__;
  wire __963__;
  wire __964__;
  wire __965__;
  wire __966__;
  wire __967__;
  wire __968__;
  wire __969__;
  wire __970__;
  wire __971__;
  wire __972__;
  wire __973__;
  wire __974__;
  wire __975__;
  wire __976__;
  wire __977__;
  wire __978__;
  wire __979__;
  wire __980__;
  wire __981__;
  wire __982__;
  wire __983__;
  wire __984__;
  wire __985__;
  wire __986__;
  wire __987__;
  wire __988__;
  wire __989__;
  wire __990__;
  wire __991__;
  wire __992__;
  wire __993__;
  wire __994__;
  wire __995__;
  wire __996__;
  wire __997__;
  wire __998__;
  wire __999__;
  wire __1000__;
  wire __1001__;
  wire __1002__;
  wire __1003__;
  wire __1004__;
  wire __1005__;
  wire __1006__;
  wire __1007__;
  wire __1008__;
  wire __1009__;
  wire __1010__;
  wire __1011__;
  wire __1012__;
  wire __1013__;
  wire __1014__;
  wire __1015__;
  wire __1016__;
  wire __1017__;
  wire __1018__;
  wire __1019__;
  wire __1020__;
  wire __1021__;
  wire __1022__;
  wire __1023__;
  wire __1024__;
  wire __1025__;
  wire __1026__;
  wire __1027__;
  wire __1028__;
  wire __1029__;
  wire __1030__;
  wire __1031__;
  wire __1032__;
  wire __1033__;
  wire __1034__;
  wire __1035__;
  wire __1036__;
  wire __1037__;
  wire __1038__;
  wire __1039__;
  wire __1040__;
  wire __1041__;
  wire __1042__;
  wire __1043__;
  wire __1044__;
  wire __1045__;
  wire __1046__;
  wire __1047__;
  wire __1048__;
  wire __1049__;
  wire __1050__;
  wire __1051__;
  wire __1052__;
  wire __1053__;
  wire __1054__;
  wire __1055__;
  wire __1056__;
  wire __1057__;
  wire __1058__;
  wire __1059__;
  wire __1060__;
  wire __1061__;
  wire __1062__;
  wire __1063__;
  wire __1064__;
  wire __1065__;
  wire __1066__;
  wire __1067__;
  wire __1068__;
  wire __1069__;
  wire __1070__;
  wire __1071__;
  wire __1072__;
  wire __1073__;
  wire __1074__;
  wire __1075__;
  wire __1076__;
  wire __1077__;
  wire __1078__;
  wire __1079__;
  wire __1080__;
  wire __1081__;
  wire __1082__;
  wire __1083__;
  wire __1084__;
  wire __1085__;
  wire __1086__;
  wire __1087__;
  wire __1088__;
  wire __1089__;
  wire __1090__;
  wire __1091__;
  wire __1092__;
  wire __1093__;
  wire __1094__;
  wire __1095__;
  wire __1096__;
  wire __1097__;
  wire __1098__;
  wire __1099__;
  wire __1100__;
  wire __1101__;
  wire __1102__;
  wire __1103__;
  wire __1104__;
  wire __1105__;
  wire __1106__;
  wire __1107__;
  wire __1108__;
  wire __1109__;
  wire __1110__;
  wire __1111__;
  wire __1112__;
  wire __1113__;
  wire __1114__;
  wire __1115__;
  wire __1116__;
  wire __1117__;
  wire __1118__;
  wire __1119__;
  wire __1120__;
  wire __1121__;
  wire __1122__;
  wire __1123__;
  wire __1124__;
  wire __1125__;
  wire __1126__;
  wire __1127__;
  wire __1128__;
  wire __1129__;
  wire __1130__;
  wire __1131__;
  wire __1132__;
  wire __1133__;
  wire __1134__;
  wire __1135__;
  wire __1136__;
  wire __1137__;
  wire __1138__;
  wire __1139__;
  wire __1140__;
  wire __1141__;
  wire __1142__;
  wire __1143__;
  wire __1144__;
  wire __1145__;
  wire __1146__;
  wire __1147__;
  wire __1148__;
  wire __1149__;
  wire __1150__;
  wire __1151__;
  wire __1152__;
  wire __1153__;
  wire __1154__;
  wire __1155__;
  wire __1156__;
  wire __1157__;
  wire __1158__;
  wire __1159__;
  wire __1160__;
  wire __1161__;
  wire __1162__;
  wire __1163__;
  wire __1164__;
  wire __1165__;
  wire __1166__;
  wire __1167__;
  wire __1168__;
  wire __1169__;
  wire __1170__;
  wire __1171__;
  wire __1172__;
  wire __1173__;
  wire __1174__;
  wire __1175__;
  wire __1176__;
  wire __1177__;
  wire __1178__;
  wire __1179__;
  wire __1180__;
  wire __1181__;
  wire __1182__;
  wire __1183__;
  wire __1184__;
  wire __1185__;
  wire __1186__;
  wire __1187__;
  wire __1188__;
  wire __1189__;
  wire __1190__;
  wire __1191__;
  wire __1192__;
  wire __1193__;
  wire __1194__;
  wire __1195__;
  wire __1196__;
  wire __1197__;
  wire __1198__;
  wire __1199__;
  wire __1200__;
  wire __1201__;
  wire __1202__;
  wire __1203__;
  wire __1204__;
  wire __1205__;
  wire __1206__;
  wire __1207__;
  wire __1208__;
  wire __1209__;
  wire __1210__;
  wire __1211__;
  wire __1212__;
  wire __1213__;
  wire __1214__;
  wire __1215__;
  wire __1216__;
  wire __1217__;
  wire __1218__;
  wire __1219__;
  wire __1220__;
  wire __1221__;
  wire __1222__;
  wire __1223__;
  wire __1224__;
  wire __1225__;
  wire __1226__;
  wire __1227__;
  wire __1228__;
  wire __1229__;
  wire __1230__;
  wire __1231__;
  wire __1232__;
  wire __1233__;
  wire __1234__;
  wire __1235__;
  wire __1236__;
  wire __1237__;
  wire __1238__;
  wire __1239__;
  wire __1240__;
  wire __1241__;
  wire __1242__;
  wire __1243__;
  wire __1244__;
  wire __1245__;
  wire __1246__;
  wire __1247__;
  wire __1248__;
  wire __1249__;
  wire __1250__;
  wire __1251__;
  wire __1252__;
  wire __1253__;
  wire __1254__;
  wire __1255__;
  wire __1256__;
  wire __1257__;
  wire __1258__;
  wire __1259__;
  wire __1260__;
  wire __1261__;
  wire __1262__;
  wire __1263__;
  wire __1264__;
  wire __1265__;
  wire __1266__;
  wire __1267__;
  wire __1268__;
  wire __1269__;
  wire __1270__;
  wire __1271__;
  wire __1272__;
  wire __1273__;
  wire __1274__;
  wire __1275__;
  wire __1276__;
  wire __1277__;
  wire __1278__;
  wire __1279__;
  wire __1280__;
  wire __1281__;
  wire __1282__;
  wire __1283__;
  wire __1284__;
  wire __1285__;
  wire __1286__;
  wire __1287__;
  wire __1288__;
  wire __1289__;
  wire __1290__;
  wire __1291__;
  wire __1292__;
  wire __1293__;
  wire __1294__;
  wire __1295__;
  wire __1296__;
  wire __1297__;
  wire __1298__;
  wire __1299__;
  wire __1300__;
  wire __1301__;
  wire __1302__;
  wire __1303__;
  wire __1304__;
  wire __1305__;
  wire __1306__;
  wire __1307__;
  wire __1308__;
  wire __1309__;
  wire __1310__;
  wire __1311__;
  wire __1312__;
  wire __1313__;
  wire __1314__;
  wire __1315__;
  wire __1316__;
  wire __1317__;
  wire __1318__;
  wire __1319__;
  wire __1320__;
  wire __1321__;
  wire __1322__;
  wire __1323__;
  wire __1324__;
  wire __1325__;
  wire __1326__;
  wire __1327__;
  wire __1328__;
  wire __1329__;
  wire __1330__;
  wire __1331__;
  wire __1332__;
  wire __1333__;
  wire __1334__;
  wire __1335__;
  wire __1336__;
  wire __1337__;
  wire __1338__;
  wire __1339__;
  wire __1340__;
  wire __1341__;
  wire __1342__;
  wire __1343__;
  wire __1344__;
  wire __1345__;
  wire __1346__;
  wire __1347__;
  wire __1348__;
  wire __1349__;
  wire __1350__;
  wire __1351__;
  wire __1352__;
  wire __1353__;
  wire __1354__;
  wire __1355__;
  wire __1356__;
  wire __1357__;
  wire __1358__;
  wire __1359__;
  wire __1360__;
  wire __1361__;
  wire __1362__;
  wire __1363__;
  wire __1364__;
  wire __1365__;
  wire __1366__;
  wire __1367__;
  wire __1368__;
  wire __1369__;
  wire __1370__;
  INV __1371__ (
    .I(g1700),
    .O(__0__)
  );
  INV __1372__ (
    .I(__119__),
    .O(__1__)
  );
  INV __1373__ (
    .I(g23),
    .O(__2__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1374__ (
    .D(__1244__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__3__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1375__ (
    .D(__1332__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__4__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1376__ (
    .D(__727__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__5__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1377__ (
    .D(__853__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__6__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1378__ (
    .D(__1133__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__7__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1379__ (
    .D(__1340__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__8__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1380__ (
    .D(__1160__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__9__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1381__ (
    .D(__951__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__10__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1382__ (
    .D(__1181__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__11__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1383__ (
    .D(__940__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__12__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1384__ (
    .D(__1360__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__13__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1385__ (
    .D(__1275__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__14__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1386__ (
    .D(__1346__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__15__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1387__ (
    .D(__943__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__16__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1388__ (
    .D(__1051__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__17__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1389__ (
    .D(__971__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__18__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1390__ (
    .D(__917__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__19__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1391__ (
    .D(__1154__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__20__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1392__ (
    .D(__500__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__21__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1393__ (
    .D(__924__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__22__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1394__ (
    .D(__1364__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__23__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1395__ (
    .D(__906__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__24__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1396__ (
    .D(__1159__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__25__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1397__ (
    .D(__1325__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__26__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1398__ (
    .D(__882__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__27__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1399__ (
    .D(__439__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__28__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1400__ (
    .D(__1169__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__29__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1401__ (
    .D(__1066__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__30__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1402__ (
    .D(__1186__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__31__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1403__ (
    .D(__1026__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__32__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1404__ (
    .D(__1063__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__33__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1405__ (
    .D(__1000__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__34__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1406__ (
    .D(__894__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__35__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1407__ (
    .D(__1249__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__36__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1408__ (
    .D(__1344__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__37__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1409__ (
    .D(__1239__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__38__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1410__ (
    .D(__987__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__39__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1411__ (
    .D(__1005__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__40__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1412__ (
    .D(__1079__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__41__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1413__ (
    .D(__899__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__42__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1414__ (
    .D(__1108__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__43__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1415__ (
    .D(__897__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__44__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1416__ (
    .D(__704__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__45__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1417__ (
    .D(__809__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__46__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1418__ (
    .D(__1151__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__47__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1419__ (
    .D(__993__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__48__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1420__ (
    .D(__1313__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__49__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1421__ (
    .D(__1033__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__50__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1422__ (
    .D(__1109__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__51__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1423__ (
    .D(__1197__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__52__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1424__ (
    .D(__931__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__53__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1425__ (
    .D(__1227__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__54__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1426__ (
    .D(__896__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__55__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1427__ (
    .D(__1028__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__56__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1428__ (
    .D(__1073__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__57__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1429__ (
    .D(__1359__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__58__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1430__ (
    .D(g83),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__59__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1431__ (
    .D(__1216__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__60__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1432__ (
    .D(__1193__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__61__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1433__ (
    .D(__838__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__62__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1434__ (
    .D(__779__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__63__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1435__ (
    .D(__1229__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__64__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1436__ (
    .D(__828__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__65__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1437__ (
    .D(__1157__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__66__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1438__ (
    .D(__1184__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__67__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1439__ (
    .D(__1047__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__68__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1440__ (
    .D(__1291__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__69__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1441__ (
    .D(__1046__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__70__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1442__ (
    .D(__744__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__71__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1443__ (
    .D(__925__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__72__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1444__ (
    .D(__1299__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__73__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1445__ (
    .D(__960__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__74__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1446__ (
    .D(__72__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__75__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1447__ (
    .D(__1087__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__76__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1448__ (
    .D(__1306__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__77__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1449__ (
    .D(__840__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__78__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1450__ (
    .D(__1363__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__79__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1451__ (
    .D(__839__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__80__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1452__ (
    .D(__1001__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__81__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1453__ (
    .D(__876__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__82__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1454__ (
    .D(__1254__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__83__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1455__ (
    .D(__1295__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__84__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1456__ (
    .D(__869__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__85__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1457__ (
    .D(__1037__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__86__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1458__ (
    .D(__1166__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__87__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1459__ (
    .D(__851__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__88__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1460__ (
    .D(__1240__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__89__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1461__ (
    .D(__743__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__90__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1462__ (
    .D(__877__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__91__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1463__ (
    .D(__1316__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__92__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1464__ (
    .D(__778__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__93__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1465__ (
    .D(__1158__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__94__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1466__ (
    .D(__738__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__95__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1467__ (
    .D(__1152__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__96__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1468__ (
    .D(__856__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__97__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1469__ (
    .D(__1202__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__98__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1470__ (
    .D(__946__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__99__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1471__ (
    .D(__1338__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__100__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1472__ (
    .D(__791__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__101__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1473__ (
    .D(__915__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__102__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1474__ (
    .D(__1149__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__103__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1475__ (
    .D(__997__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__104__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1476__ (
    .D(__852__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__105__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1477__ (
    .D(__1311__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__106__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1478__ (
    .D(__1237__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__107__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1479__ (
    .D(__1298__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__108__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1480__ (
    .D(__995__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__109__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1481__ (
    .D(__1256__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__110__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1482__ (
    .D(__1230__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__111__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1483__ (
    .D(__1103__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__112__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1484__ (
    .D(__1233__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__113__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1485__ (
    .D(__452__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__114__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1486__ (
    .D(__1080__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__115__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1487__ (
    .D(__830__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__116__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1488__ (
    .D(__964__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__117__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1489__ (
    .D(__949__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__118__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1490__ (
    .D(__29__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__119__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1491__ (
    .D(__726__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__120__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1492__ (
    .D(__1293__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__121__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1493__ (
    .D(__740__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__122__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1494__ (
    .D(__337__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__123__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1495__ (
    .D(__421__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__124__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1496__ (
    .D(__1125__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__125__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1497__ (
    .D(__1170__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__126__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1498__ (
    .D(__928__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__127__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1499__ (
    .D(__1176__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__128__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1500__ (
    .D(__1309__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__129__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1501__ (
    .D(__1145__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__130__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1502__ (
    .D(__945__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__131__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1503__ (
    .D(__1031__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__132__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1504__ (
    .D(__1164__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__133__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1505__ (
    .D(__1058__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__134__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1506__ (
    .D(__1141__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__135__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1507__ (
    .D(__1361__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__136__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1508__ (
    .D(__1196__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__137__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1509__ (
    .D(__246__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__138__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1510__ (
    .D(__837__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__139__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1511__ (
    .D(__773__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__140__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1512__ (
    .D(__1204__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__141__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1513__ (
    .D(__914__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__142__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1514__ (
    .D(__921__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__143__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1515__ (
    .D(__1334__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__144__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1516__ (
    .D(__682__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__145__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1517__ (
    .D(__1290__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__146__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1518__ (
    .D(__957__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__147__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1519__ (
    .D(__1140__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__148__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1520__ (
    .D(__1209__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__149__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1521__ (
    .D(__999__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__150__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1522__ (
    .D(__1323__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__151__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1523__ (
    .D(__825__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__152__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1524__ (
    .D(g103),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__153__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1525__ (
    .D(__991__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__154__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1526__ (
    .D(__911__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__155__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1527__ (
    .D(__1179__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__156__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1528__ (
    .D(__1232__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__157__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1529__ (
    .D(g28),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__158__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1530__ (
    .D(__975__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__159__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1531__ (
    .D(__1214__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__160__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1532__ (
    .D(__1162__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__161__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1533__ (
    .D(__1171__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__162__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1534__ (
    .D(__848__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__163__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1535__ (
    .D(__905__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__164__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1536__ (
    .D(__1297__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__165__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1537__ (
    .D(__998__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__166__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1538__ (
    .D(__1136__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__167__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1539__ (
    .D(__59__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__168__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1540__ (
    .D(__398__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__169__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1541__ (
    .D(__106__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__170__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1542__ (
    .D(__1182__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__171__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1543__ (
    .D(__1034__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__172__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1544__ (
    .D(__810__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__173__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1545__ (
    .D(__1187__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__174__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1546__ (
    .D(__1349__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__175__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1547__ (
    .D(__887__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__176__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1548__ (
    .D(__1024__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__177__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1549__ (
    .D(__855__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__178__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1550__ (
    .D(__1307__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__179__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1551__ (
    .D(g102),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__180__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1552__ (
    .D(__1175__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__181__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1553__ (
    .D(__763__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__182__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1554__ (
    .D(__36__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__183__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1555__ (
    .D(__1358__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__184__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1556__ (
    .D(__820__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__185__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1557__ (
    .D(__934__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__186__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1558__ (
    .D(__664__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__187__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1559__ (
    .D(__952__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__188__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1560__ (
    .D(__1320__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__189__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1561__ (
    .D(__1188__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__190__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1562__ (
    .D(__977__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__191__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1563__ (
    .D(__806__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__192__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1564__ (
    .D(__1343__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__193__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1565__ (
    .D(__1200__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__194__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1566__ (
    .D(__1135__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__195__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1567__ (
    .D(__168__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__196__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1568__ (
    .D(__1337__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__197__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1569__ (
    .D(__489__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__198__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1570__ (
    .D(__955__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__199__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1571__ (
    .D(__1177__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__200__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1572__ (
    .D(__1370__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__201__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1573__ (
    .D(__824__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__202__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1574__ (
    .D(__1210__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__203__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1575__ (
    .D(__844__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__204__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1576__ (
    .D(__1190__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__205__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1577__ (
    .D(__1246__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__206__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1578__ (
    .D(__1191__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__207__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1579__ (
    .D(__966__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__208__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1580__ (
    .D(__1173__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__209__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1581__ (
    .D(__1350__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__210__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1582__ (
    .D(__1096__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__211__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1583__ (
    .D(__1100__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__212__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1584__ (
    .D(__57__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__213__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1585__ (
    .D(__1035__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__214__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1586__ (
    .D(__1327__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__215__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1587__ (
    .D(__793__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__216__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1588__ (
    .D(__1105__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__217__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1589__ (
    .D(__1004__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__218__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1590__ (
    .D(__900__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__219__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1591__ (
    .D(__958__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__220__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1592__ (
    .D(__994__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__221__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1593__ (
    .D(__1228__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__222__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1594__ (
    .D(__706__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__223__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1595__ (
    .D(__967__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__224__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1596__ (
    .D(__1238__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__225__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1597__ (
    .D(__742__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__226__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1598__ (
    .D(__1331__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__227__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1599__ (
    .D(__739__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__228__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1600__ (
    .D(__27__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__229__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1601__ (
    .D(__1107__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__230__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1602__ (
    .D(__287__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__231__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1603__ (
    .D(__941__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__232__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1604__ (
    .D(g29),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__233__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1605__ (
    .D(__1139__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__234__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1606__ (
    .D(__1294__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__235__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1607__ (
    .D(__850__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__236__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1608__ (
    .D(__754__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__237__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1609__ (
    .D(__1120__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__238__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1610__ (
    .D(__1148__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__239__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1611__ (
    .D(__1044__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__240__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1612__ (
    .D(__1113__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__241__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1613__ (
    .D(__950__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__242__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1614__ (
    .D(__992__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__243__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1615__ (
    .D(__795__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__244__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1616__ (
    .D(__460__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__245__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1617__ (
    .D(__1278__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__246__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1618__ (
    .D(__1064__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__247__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1619__ (
    .D(__1088__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__248__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1620__ (
    .D(__338__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__249__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1621__ (
    .D(__705__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__250__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1622__ (
    .D(__1362__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__251__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1623__ (
    .D(__1213__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__252__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1624__ (
    .D(__776__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__253__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1625__ (
    .D(__1315__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__254__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1626__ (
    .D(__1212__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__255__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1627__ (
    .D(__1218__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__256__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1628__ (
    .D(__908__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__257__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1629__ (
    .D(__513__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__258__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1630__ (
    .D(__518__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__259__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1631__ (
    .D(__1195__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__260__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1632__ (
    .D(__1314__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__261__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1633__ (
    .D(__1077__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__262__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1634__ (
    .D(__821__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__263__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1635__ (
    .D(__919__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__264__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1636__ (
    .D(__1156__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__265__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1637__ (
    .D(__989__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__266__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1638__ (
    .D(__1057__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__267__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1639__ (
    .D(__1002__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__268__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1640__ (
    .D(__927__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__269__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1641__ (
    .D(__1303__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__270__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1642__ (
    .D(__854__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__271__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1643__ (
    .D(__932__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__272__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1644__ (
    .D(__956__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__273__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1645__ (
    .D(__774__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__274__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1646__ (
    .D(__983__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__275__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1647__ (
    .D(__953__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__276__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1648__ (
    .D(__751__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__277__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1649__ (
    .D(__196__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__278__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1650__ (
    .D(__1368__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__279__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1651__ (
    .D(__1091__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__280__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1652__ (
    .D(__974__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__281__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1653__ (
    .D(__807__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__282__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1654__ (
    .D(__768__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__283__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1655__ (
    .D(__823__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__284__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1656__ (
    .D(__1300__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__285__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1657__ (
    .D(__761__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__286__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1658__ (
    .D(__1348__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__287__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1659__ (
    .D(__1248__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__288__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1660__ (
    .D(__1095__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__289__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1661__ (
    .D(__205__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__290__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1662__ (
    .D(__980__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__291__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1663__ (
    .D(__1045__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__292__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1664__ (
    .D(__868__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__293__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1665__ (
    .D(__745__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__294__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1666__ (
    .D(__962__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__295__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1667__ (
    .D(__1357__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__296__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1668__ (
    .D(__1356__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__297__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1669__ (
    .D(__1207__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__298__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1670__ (
    .D(__182__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__299__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1671__ (
    .D(__1150__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__300__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1672__ (
    .D(__367__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__301__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1673__ (
    .D(__923__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__302__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1674__ (
    .D(g101),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__303__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1675__ (
    .D(__990__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__304__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1676__ (
    .D(__1211__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__305__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1677__ (
    .D(__1276__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__306__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1678__ (
    .D(__132__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__307__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1679__ (
    .D(__752__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__308__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1680__ (
    .D(__750__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__309__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1681__ (
    .D(__1043__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__310__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1682__ (
    .D(__1022__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__311__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1683__ (
    .D(__849__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__312__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1684__ (
    .D(__1285__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__313__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1685__ (
    .D(__1367__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__314__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1686__ (
    .D(__984__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__315__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1687__ (
    .D(__808__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__316__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1688__ (
    .D(__842__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__317__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1689__ (
    .D(__515__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__318__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1690__ (
    .D(__1163__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__319__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1691__ (
    .D(__701__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__320__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1692__ (
    .D(__891__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__321__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1693__ (
    .D(__1242__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__322__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1694__ (
    .D(__1180__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__323__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1695__ (
    .D(__969__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__324__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1696__ (
    .D(__947__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__325__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1697__ (
    .D(__910__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__326__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1698__ (
    .D(__973__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__327__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1699__ (
    .D(__788__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__328__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1700__ (
    .D(__1123__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__329__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1701__ (
    .D(__1292__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__330__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1702__ (
    .D(g104),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__331__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1703__ (
    .D(__1065__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__332__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1704__ (
    .D(__1236__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__333__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1705__ (
    .D(__1147__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__334__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1706__ (
    .D(__1250__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__335__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1707__ (
    .D(__1284__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__336__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1708__ (
    .D(__861__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__337__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1709__ (
    .D(__758__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__338__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1710__ (
    .D(__710__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__339__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1711__ (
    .D(__127__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__340__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1712__ (
    .D(__1347__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__341__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1713__ (
    .D(__922__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__342__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1714__ (
    .D(__1076__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__343__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1715__ (
    .D(__800__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__344__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1716__ (
    .D(__1161__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__345__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1717__ (
    .D(__858__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__346__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1718__ (
    .D(__1025__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__347__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1719__ (
    .D(__1324__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__348__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1720__ (
    .D(__1245__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__349__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1721__ (
    .D(__1174__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__350__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1722__ (
    .D(__1206__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__351__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1723__ (
    .D(__1116__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__352__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1724__ (
    .D(__1247__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__353__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1725__ (
    .D(__1266__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__354__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1726__ (
    .D(__1092__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__355__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1727__ (
    .D(__979__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__356__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1728__ (
    .D(__1132__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__357__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1729__ (
    .D(__1355__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__358__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1730__ (
    .D(__796__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__359__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1731__ (
    .D(__1234__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__360__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1732__ (
    .D(__753__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__361__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1733__ (
    .D(__1115__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__362__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1734__ (
    .D(__1283__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__363__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1735__ (
    .D(__948__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__364__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1736__ (
    .D(__832__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__365__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1737__ (
    .D(__1155__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__366__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1738__ (
    .D(__798__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__367__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1739__ (
    .D(__893__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__368__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1740__ (
    .D(__50__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__369__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1741__ (
    .D(__1366__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__370__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1742__ (
    .D(__1302__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__371__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1743__ (
    .D(__1351__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__372__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1744__ (
    .D(__978__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__373__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1745__ (
    .D(__959__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__374__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1746__ (
    .D(__907__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__375__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1747__ (
    .D(__1253__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__376__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1748__ (
    .D(__886__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__377__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1749__ (
    .D(__1322__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__378__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1750__ (
    .D(__1121__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__379__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1751__ (
    .D(__680__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__380__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1752__ (
    .D(__816__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__381__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1753__ (
    .D(__757__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__382__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1754__ (
    .D(__0__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__383__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1755__ (
    .D(__1329__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__384__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1756__ (
    .D(__909__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__385__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1757__ (
    .D(__827__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__386__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1758__ (
    .D(__826__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__387__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1759__ (
    .D(__885__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__388__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1760__ (
    .D(__1165__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__389__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1761__ (
    .D(__1106__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__390__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1762__ (
    .D(__845__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__391__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1763__ (
    .D(__741__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__392__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1764__ (
    .D(__87__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__393__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1765__ (
    .D(__200__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__394__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1766__ (
    .D(__1194__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__395__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1767__ (
    .D(__509__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__396__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1768__ (
    .D(__920__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__397__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1769__ (
    .D(__1118__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__398__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1770__ (
    .D(__1199__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__399__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1771__ (
    .D(__926__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__400__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1772__ (
    .D(__937__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__401__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1773__ (
    .D(__898__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__402__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1774__ (
    .D(__1049__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__403__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1775__ (
    .D(__1198__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__404__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1776__ (
    .D(__1138__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__405__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1777__ (
    .D(__883__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__406__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1778__ (
    .D(__154__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__407__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1779__ (
    .D(__1084__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__408__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1780__ (
    .D(__1352__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__409__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1781__ (
    .D(__1336__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__410__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1782__ (
    .D(__1260__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__411__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1783__ (
    .D(__1007__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__412__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1784__ (
    .D(__1262__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__413__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1785__ (
    .D(__1111__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__414__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1786__ (
    .D(__1006__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__415__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1787__ (
    .D(__1243__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__416__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1788__ (
    .D(__1078__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__417__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1789__ (
    .D(__430__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__418__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1790__ (
    .D(__769__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__419__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1791__ (
    .D(__1257__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__420__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1792__ (
    .D(__1119__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__421__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1793__ (
    .D(__1265__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__422__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1794__ (
    .D(__1143__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__423__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1795__ (
    .D(__976__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__424__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1796__ (
    .D(__772__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__425__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1797__ (
    .D(__737__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__426__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1798__ (
    .D(__703__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__427__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1799__ (
    .D(__675__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__428__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1800__ (
    .D(__1274__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__429__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1801__ (
    .D(__1030__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__430__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1802__ (
    .D(__1269__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__431__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1803__ (
    .D(__770__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__432__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1804__ (
    .D(__296__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__433__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1805__ (
    .D(__749__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__434__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1806__ (
    .D(__1231__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__435__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1807__ (
    .D(__1142__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__436__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1808__ (
    .D(__1124__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__437__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1809__ (
    .D(__970__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__438__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1810__ (
    .D(__1029__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__439__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1811__ (
    .D(__736__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__440__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1812__ (
    .D(__1131__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__441__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1813__ (
    .D(__930__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__442__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1814__ (
    .D(__836__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__443__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1815__ (
    .D(__1339__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__444__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1816__ (
    .D(__936__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__445__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1817__ (
    .D(__944__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__446__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1818__ (
    .D(__819__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__447__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1819__ (
    .D(__818__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__448__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1820__ (
    .D(__867__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__449__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1821__ (
    .D(__766__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__450__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1822__ (
    .D(__1146__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__451__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1823__ (
    .D(__1268__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__452__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1824__ (
    .D(__1094__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__453__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1825__ (
    .D(__822__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__454__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1826__ (
    .D(__1241__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__455__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1827__ (
    .D(__1153__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__456__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1828__ (
    .D(__1341__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__457__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1829__ (
    .D(__866__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__458__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1830__ (
    .D(__916__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__459__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1831__ (
    .D(__1205__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__460__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1832__ (
    .D(__782__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__461__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1833__ (
    .D(__1317__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__462__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1834__ (
    .D(__1185__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__463__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1835__ (
    .D(__986__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__464__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1836__ (
    .D(__765__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__465__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1837__ (
    .D(__1019__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__466__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1838__ (
    .D(__681__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__467__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1839__ (
    .D(__1277__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__468__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1840__ (
    .D(__1345__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__469__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1841__ (
    .D(__1093__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__470__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1842__ (
    .D(__1130__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__471__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1843__ (
    .D(__1075__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__472__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1844__ (
    .D(__1330__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__473__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1845__ (
    .D(__890__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__474__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1846__ (
    .D(__835__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__475__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1847__ (
    .D(__1134__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__476__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1848__ (
    .D(__1267__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__477__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1849__ (
    .D(__688__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__478__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1850__ (
    .D(__903__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__479__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1851__ (
    .D(__1252__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__480__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1852__ (
    .D(__1129__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__481__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1853__ (
    .D(__1203__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__482__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1854__ (
    .D(__1261__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__483__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1855__ (
    .D(__266__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__484__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1856__ (
    .D(__235__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__485__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1857__ (
    .D(__1235__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__486__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1858__ (
    .D(__1310__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__487__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1859__ (
    .D(__892__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__488__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1860__ (
    .D(__1089__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__489__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1861__ (
    .D(__1264__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__490__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1862__ (
    .D(__929__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__491__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1863__ (
    .D(__1128__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__492__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1864__ (
    .D(__735__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__493__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1865__ (
    .D(__1342__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__494__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1866__ (
    .D(__1042__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__495__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1867__ (
    .D(__111__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__496__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1868__ (
    .D(__684__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__497__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1869__ (
    .D(__470__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__498__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1870__ (
    .D(__1328__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__499__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1871__ (
    .D(__857__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__500__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1872__ (
    .D(__371__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__501__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1873__ (
    .D(__1012__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__502__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1874__ (
    .D(__865__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__503__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1875__ (
    .D(__1189__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__504__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1876__ (
    .D(__1112__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__505__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __1877__ (
    .D(__1099__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__506__)
  );
  LUT4 #(
    .INIT(16'h0010)
  ) __1879__ (
    .I3(__11__),
    .I2(__5__),
    .I1(g1696),
    .I0(__154__),
    .O(__508__)
  );
  LUT4 #(
    .INIT(16'hf088)
  ) __1880__ (
    .I3(__508__),
    .I2(__355__),
    .I1(g109),
    .I0(__396__),
    .O(__509__)
  );
  LUT4 #(
    .INIT(16'h0001)
  ) __1882__ (
    .I3(__295__),
    .I2(__414__),
    .I1(__112__),
    .I0(__273__),
    .O(__511__)
  );
  LUT5 #(
    .INIT(32'h00000004)
  ) __1883__ (
    .I4(__333__),
    .I3(__309__),
    .I2(__261__),
    .I1(__118__),
    .I0(__269__),
    .O(__512__)
  );
  LUT6 #(
    .INIT(64'h0caa0c0c0c0c0c0c)
  ) __1884__ (
    .I5(__56__),
    .I4(__512__),
    .I3(__295__),
    .I2(__511__),
    .I1(__258__),
    .I0(__416__),
    .O(__513__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __1885__ (
    .I2(__47__),
    .I1(__506__),
    .I0(__329__),
    .O(__514__)
  );
  LUT4 #(
    .INIT(16'hbf80)
  ) __1886__ (
    .I3(__318__),
    .I2(__38__),
    .I1(__150__),
    .I0(__116__),
    .O(__515__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __1887__ (
    .I1(__222__),
    .I0(__279__),
    .O(__516__)
  );
  LUT6 #(
    .INIT(64'h555555553000cfff)
  ) __1888__ (
    .I5(g18),
    .I4(__315__),
    .I3(__516__),
    .I2(__149__),
    .I1(__400__),
    .I0(__24__),
    .O(__517__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __1889__ (
    .I2(g109),
    .I1(__210__),
    .I0(__517__),
    .O(__518__)
  );
  LUT3 #(
    .INIT(8'h40)
  ) __1890__ (
    .I2(g109),
    .I1(__338__),
    .I0(__249__),
    .O(__519__)
  );
  LUT4 #(
    .INIT(16'h9009)
  ) __1891__ (
    .I3(__501__),
    .I2(__272__),
    .I1(__123__),
    .I0(__165__),
    .O(__520__)
  );
  LUT2 #(
    .INIT(4'h9)
  ) __1892__ (
    .I1(__75__),
    .I0(__410__),
    .O(__521__)
  );
  LUT6 #(
    .INIT(64'h9009000000000000)
  ) __1893__ (
    .I5(__521__),
    .I4(__520__),
    .I3(__498__),
    .I2(__88__),
    .I1(__496__),
    .I0(__208__),
    .O(__522__)
  );
  LUT6 #(
    .INIT(64'hb00b00000000b00b)
  ) __1894__ (
    .I5(__290__),
    .I4(__347__),
    .I3(__369__),
    .I2(__188__),
    .I1(__99__),
    .I0(__231__),
    .O(__523__)
  );
  LUT6 #(
    .INIT(64'hb00b000000000000)
  ) __1895__ (
    .I5(__523__),
    .I4(__522__),
    .I3(__307__),
    .I2(__162__),
    .I1(__231__),
    .I0(__99__),
    .O(__524__)
  );
  LUT6 #(
    .INIT(64'h0000000000000001)
  ) __1896__ (
    .I5(__162__),
    .I4(__188__),
    .I3(__208__),
    .I2(__272__),
    .I1(__499__),
    .I0(__7__),
    .O(__525__)
  );
  LUT3 #(
    .INIT(8'h01)
  ) __1897__ (
    .I2(__136__),
    .I1(__347__),
    .I0(__99__),
    .O(__526__)
  );
  LUT6 #(
    .INIT(64'h0000000000000040)
  ) __1898__ (
    .I5(__420__),
    .I4(__410__),
    .I3(__88__),
    .I2(__526__),
    .I1(__525__),
    .I0(__165__),
    .O(__527__)
  );
  LUT4 #(
    .INIT(16'h8000)
  ) __1899__ (
    .I3(__121__),
    .I2(__115__),
    .I1(__104__),
    .I0(__436__),
    .O(__528__)
  );
  LUT5 #(
    .INIT(32'hf0053333)
  ) __1900__ (
    .I4(__528__),
    .I3(__361__),
    .I2(__399__),
    .I1(__340__),
    .I0(__527__),
    .O(__529__)
  );
  LUT5 #(
    .INIT(32'h10000000)
  ) __1901__ (
    .I4(g48),
    .I3(g42),
    .I2(g43),
    .I1(g44),
    .I0(g45),
    .O(__530__)
  );
  LUT5 #(
    .INIT(32'h00000040)
  ) __1902__ (
    .I4(g42),
    .I3(g44),
    .I2(g48),
    .I1(g43),
    .I0(g45),
    .O(__531__)
  );
  LUT6 #(
    .INIT(64'h0000000500000003)
  ) __1903__ (
    .I5(g48),
    .I4(g41),
    .I3(g46),
    .I2(g47),
    .I1(g30),
    .I0(g31),
    .O(__532__)
  );
  LUT3 #(
    .INIT(8'h1f)
  ) __1904__ (
    .I2(__532__),
    .I1(__531__),
    .I0(__530__),
    .O(__533__)
  );
  LUT6 #(
    .INIT(64'h0000000010000000)
  ) __1905__ (
    .I5(g41),
    .I4(g48),
    .I3(g44),
    .I2(g43),
    .I1(g42),
    .I0(g45),
    .O(__534__)
  );
  LUT5 #(
    .INIT(32'h00008000)
  ) __1906__ (
    .I4(g45),
    .I3(g48),
    .I2(g42),
    .I1(g44),
    .I0(g43),
    .O(__535__)
  );
  LUT5 #(
    .INIT(32'h00000040)
  ) __1907__ (
    .I4(g42),
    .I3(g44),
    .I2(g48),
    .I1(g45),
    .I0(g43),
    .O(__536__)
  );
  LUT5 #(
    .INIT(32'h10000000)
  ) __1908__ (
    .I4(g48),
    .I3(g42),
    .I2(g45),
    .I1(g44),
    .I0(g43),
    .O(__537__)
  );
  LUT6 #(
    .INIT(64'h0005000300000000)
  ) __1909__ (
    .I5(g47),
    .I4(g48),
    .I3(g41),
    .I2(g46),
    .I1(g30),
    .I0(g31),
    .O(__538__)
  );
  LUT6 #(
    .INIT(64'h000100010001ffff)
  ) __1910__ (
    .I5(__532__),
    .I4(__538__),
    .I3(__537__),
    .I2(__536__),
    .I1(__535__),
    .I0(__534__),
    .O(__539__)
  );
  LUT6 #(
    .INIT(64'h0000efff00000000)
  ) __1911__ (
    .I5(g48),
    .I4(g31),
    .I3(__532__),
    .I2(g44),
    .I1(g45),
    .I0(g43),
    .O(__540__)
  );
  LUT6 #(
    .INIT(64'h0005000300000000)
  ) __1912__ (
    .I5(g46),
    .I4(g48),
    .I3(g41),
    .I2(g47),
    .I1(g30),
    .I0(g31),
    .O(__541__)
  );
  LUT6 #(
    .INIT(64'hd43fffffffffffff)
  ) __1913__ (
    .I5(g48),
    .I4(__541__),
    .I3(g45),
    .I2(g44),
    .I1(g43),
    .I0(g42),
    .O(__542__)
  );
  LUT5 #(
    .INIT(32'h00008000)
  ) __1914__ (
    .I4(g42),
    .I3(g48),
    .I2(g44),
    .I1(g45),
    .I0(g43),
    .O(__543__)
  );
  LUT5 #(
    .INIT(32'h80000000)
  ) __1915__ (
    .I4(g48),
    .I3(g42),
    .I2(g44),
    .I1(g45),
    .I0(g43),
    .O(__544__)
  );
  LUT4 #(
    .INIT(16'h01ff)
  ) __1916__ (
    .I3(__538__),
    .I2(__536__),
    .I1(__544__),
    .I0(__543__),
    .O(__545__)
  );
  LUT4 #(
    .INIT(16'h0080)
  ) __1917__ (
    .I3(g31),
    .I2(g46),
    .I1(g47),
    .I0(__534__),
    .O(__546__)
  );
  LUT6 #(
    .INIT(64'h0000000080000000)
  ) __1918__ (
    .I5(__546__),
    .I4(__545__),
    .I3(__542__),
    .I2(__540__),
    .I1(__539__),
    .I0(__533__),
    .O(__547__)
  );
  LUT6 #(
    .INIT(64'h007f7f7f7f7f7f7f)
  ) __1919__ (
    .I5(__532__),
    .I4(__530__),
    .I3(__408__),
    .I2(__537__),
    .I1(__541__),
    .I0(__458__),
    .O(__548__)
  );
  LUT5 #(
    .INIT(32'h0777ffff)
  ) __1920__ (
    .I4(__538__),
    .I3(__535__),
    .I2(g1173),
    .I1(__534__),
    .I0(g1197),
    .O(__549__)
  );
  LUT5 #(
    .INIT(32'h0777ffff)
  ) __1921__ (
    .I4(__538__),
    .I3(__537__),
    .I2(__469__),
    .I1(__536__),
    .I0(__426__),
    .O(__550__)
  );
  LUT3 #(
    .INIT(8'h35)
  ) __1922__ (
    .I2(g42),
    .I1(__342__),
    .I0(__65__),
    .O(__551__)
  );
  LUT4 #(
    .INIT(16'h0040)
  ) __1923__ (
    .I3(g45),
    .I2(g48),
    .I1(g44),
    .I0(g43),
    .O(__552__)
  );
  LUT6 #(
    .INIT(64'h00bfbfbfbfbfbfbf)
  ) __1924__ (
    .I5(__541__),
    .I4(__534__),
    .I3(g925),
    .I2(__532__),
    .I1(__552__),
    .I0(__551__),
    .O(__553__)
  );
  LUT5 #(
    .INIT(32'h00008000)
  ) __1925__ (
    .I4(g43),
    .I3(g48),
    .I2(g42),
    .I1(g44),
    .I0(g45),
    .O(__554__)
  );
  LUT6 #(
    .INIT(64'h007f7f7f7f7f7f7f)
  ) __1926__ (
    .I5(__532__),
    .I4(__531__),
    .I3(__15__),
    .I2(__541__),
    .I1(__268__),
    .I0(__554__),
    .O(__555__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __1927__ (
    .I2(g48),
    .I1(g42),
    .I0(g43),
    .O(__556__)
  );
  LUT3 #(
    .INIT(8'hb0)
  ) __1928__ (
    .I2(__294__),
    .I1(g48),
    .I0(g31),
    .O(__557__)
  );
  LUT6 #(
    .INIT(64'h00000000bfffffff)
  ) __1929__ (
    .I5(__557__),
    .I4(g45),
    .I3(__541__),
    .I2(g889),
    .I1(__556__),
    .I0(g44),
    .O(__558__)
  );
  LUT6 #(
    .INIT(64'h8000000000000000)
  ) __1930__ (
    .I5(__558__),
    .I4(__555__),
    .I3(__553__),
    .I2(__550__),
    .I1(__549__),
    .I0(__548__),
    .O(__559__)
  );
  LUT5 #(
    .INIT(32'hf0880000)
  ) __1931__ (
    .I4(__532__),
    .I3(__534__),
    .I2(__486__),
    .I1(__535__),
    .I0(__197__),
    .O(__560__)
  );
  LUT5 #(
    .INIT(32'h0777ffff)
  ) __1932__ (
    .I4(__538__),
    .I3(__544__),
    .I2(__441__),
    .I1(__543__),
    .I0(__318__),
    .O(__561__)
  );
  LUT5 #(
    .INIT(32'h0777ffff)
  ) __1933__ (
    .I4(__541__),
    .I3(__536__),
    .I2(__26__),
    .I1(__535__),
    .I0(g901),
    .O(__562__)
  );
  LUT5 #(
    .INIT(32'hf0880000)
  ) __1934__ (
    .I4(__532__),
    .I3(__536__),
    .I2(__133__),
    .I1(__537__),
    .I0(__191__),
    .O(__563__)
  );
  LUT4 #(
    .INIT(16'h0040)
  ) __1935__ (
    .I3(__563__),
    .I2(__562__),
    .I1(__561__),
    .I0(__560__),
    .O(__564__)
  );
  LUT4 #(
    .INIT(16'hbf00)
  ) __1936__ (
    .I3(g109),
    .I2(__564__),
    .I1(__559__),
    .I0(__547__),
    .O(__565__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __1937__ (
    .I2(__537__),
    .I1(__541__),
    .I0(__344__),
    .O(__566__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __1938__ (
    .I2(__541__),
    .I1(__536__),
    .I0(__298__),
    .O(__567__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __1939__ (
    .I2(__541__),
    .I1(__554__),
    .I0(__64__),
    .O(__568__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __1940__ (
    .I2(__541__),
    .I1(__535__),
    .I0(g904),
    .O(__569__)
  );
  LUT6 #(
    .INIT(64'h0000000080000000)
  ) __1941__ (
    .I5(g44),
    .I4(g48),
    .I3(g42),
    .I2(g45),
    .I1(g43),
    .I0(__541__),
    .O(__570__)
  );
  LUT6 #(
    .INIT(64'h0000000100000003)
  ) __1942__ (
    .I5(__570__),
    .I4(__569__),
    .I3(__568__),
    .I2(__567__),
    .I1(__566__),
    .I0(g892),
    .O(__571__)
  );
  LUT5 #(
    .INIT(32'hf0880000)
  ) __1943__ (
    .I4(__532__),
    .I3(__536__),
    .I2(__139__),
    .I1(__537__),
    .I0(__444__),
    .O(__572__)
  );
  LUT5 #(
    .INIT(32'h0777ffff)
  ) __1944__ (
    .I4(__538__),
    .I3(__537__),
    .I2(__427__),
    .I1(__536__),
    .I0(__397__),
    .O(__573__)
  );
  LUT5 #(
    .INIT(32'h0777ffff)
  ) __1945__ (
    .I4(__538__),
    .I3(__535__),
    .I2(g1176),
    .I1(__534__),
    .I0(g1200),
    .O(__574__)
  );
  LUT5 #(
    .INIT(32'hf0880000)
  ) __1946__ (
    .I4(__532__),
    .I3(__534__),
    .I2(__263__),
    .I1(__535__),
    .I0(__321__),
    .O(__575__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __1947__ (
    .I1(g44),
    .I0(g45),
    .O(__576__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __1948__ (
    .I1(g48),
    .I0(g43),
    .O(__577__)
  );
  LUT6 #(
    .INIT(64'hca00000000000000)
  ) __1949__ (
    .I5(__532__),
    .I4(__577__),
    .I3(__576__),
    .I2(g42),
    .I1(__312__),
    .I0(__323__),
    .O(__578__)
  );
  LUT5 #(
    .INIT(32'h00000040)
  ) __1950__ (
    .I4(__578__),
    .I3(__575__),
    .I2(__574__),
    .I1(__573__),
    .I0(__572__),
    .O(__579__)
  );
  LUT6 #(
    .INIT(64'h0000000010000000)
  ) __1951__ (
    .I5(g42),
    .I4(g48),
    .I3(__532__),
    .I2(g43),
    .I1(g44),
    .I0(g45),
    .O(__580__)
  );
  LUT6 #(
    .INIT(64'h0000000000008000)
  ) __1952__ (
    .I5(g44),
    .I4(g45),
    .I3(g48),
    .I2(__532__),
    .I1(g42),
    .I0(g43),
    .O(__581__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __1953__ (
    .I2(__538__),
    .I1(__544__),
    .I0(__454__),
    .O(__582__)
  );
  LUT5 #(
    .INIT(32'h335f3333)
  ) __1954__ (
    .I4(g48),
    .I3(g31),
    .I2(__543__),
    .I1(__274__),
    .I0(__304__),
    .O(__583__)
  );
  LUT6 #(
    .INIT(64'h0000153f00000000)
  ) __1955__ (
    .I5(__583__),
    .I4(__582__),
    .I3(__581__),
    .I2(__129__),
    .I1(__580__),
    .I0(__502__),
    .O(__584__)
  );
  LUT5 #(
    .INIT(32'hbfff0000)
  ) __1956__ (
    .I4(g109),
    .I3(__584__),
    .I2(__579__),
    .I1(__571__),
    .I0(__547__),
    .O(__585__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __1957__ (
    .I2(__538__),
    .I1(__544__),
    .I0(__431__),
    .O(__586__)
  );
  LUT5 #(
    .INIT(32'h335f3333)
  ) __1958__ (
    .I4(g48),
    .I3(g31),
    .I2(__543__),
    .I1(__425__),
    .I0(__108__),
    .O(__587__)
  );
  LUT6 #(
    .INIT(64'h0000153f00000000)
  ) __1959__ (
    .I5(__587__),
    .I4(__586__),
    .I3(__581__),
    .I2(__580__),
    .I1(__440__),
    .I0(__213__),
    .O(__588__)
  );
  LUT5 #(
    .INIT(32'hf0880000)
  ) __1960__ (
    .I4(__532__),
    .I3(__534__),
    .I2(__477__),
    .I1(__535__),
    .I0(__366__),
    .O(__589__)
  );
  LUT6 #(
    .INIT(64'h000f007700ff00ff)
  ) __1961__ (
    .I5(__532__),
    .I4(__536__),
    .I3(__589__),
    .I2(__97__),
    .I1(__537__),
    .I0(__447__),
    .O(__590__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __1962__ (
    .I2(__537__),
    .I1(__541__),
    .I0(__404__),
    .O(__591__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __1963__ (
    .I2(__541__),
    .I1(__536__),
    .I0(__223__),
    .O(__592__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __1964__ (
    .I2(__541__),
    .I1(__554__),
    .I0(__465__),
    .O(__593__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __1965__ (
    .I2(__541__),
    .I1(__535__),
    .I0(g907),
    .O(__594__)
  );
  LUT6 #(
    .INIT(64'h0000000100000003)
  ) __1966__ (
    .I5(__570__),
    .I4(__594__),
    .I3(__593__),
    .I2(__592__),
    .I1(__591__),
    .I0(g895),
    .O(__595__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __1967__ (
    .I2(__536__),
    .I1(__538__),
    .I0(__443__),
    .O(__596__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __1968__ (
    .I2(__537__),
    .I1(__538__),
    .I0(__90__),
    .O(__597__)
  );
  LUT5 #(
    .INIT(32'hca000000)
  ) __1969__ (
    .I4(__532__),
    .I3(__552__),
    .I2(g42),
    .I1(__84__),
    .I0(__46__),
    .O(__598__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __1970__ (
    .I2(__534__),
    .I1(__538__),
    .I0(g1203),
    .O(__599__)
  );
  LUT6 #(
    .INIT(64'h0000000080000000)
  ) __1971__ (
    .I5(g45),
    .I4(g48),
    .I3(g42),
    .I2(g44),
    .I1(g43),
    .I0(__538__),
    .O(__600__)
  );
  LUT6 #(
    .INIT(64'h0000000100000003)
  ) __1972__ (
    .I5(__600__),
    .I4(__599__),
    .I3(__598__),
    .I2(__597__),
    .I1(__596__),
    .I0(g1179),
    .O(__601__)
  );
  LUT6 #(
    .INIT(64'hbfffffff00000000)
  ) __1973__ (
    .I5(g109),
    .I4(__601__),
    .I3(__595__),
    .I2(__590__),
    .I1(__588__),
    .I0(__547__),
    .O(__602__)
  );
  LUT6 #(
    .INIT(64'hb0bb00000000b0bb)
  ) __1974__ (
    .I5(__299__),
    .I4(__602__),
    .I3(__28__),
    .I2(__585__),
    .I1(__21__),
    .I0(__565__),
    .O(__603__)
  );
  LUT6 #(
    .INIT(64'h00000000bfff0000)
  ) __1975__ (
    .I5(__28__),
    .I4(g109),
    .I3(__584__),
    .I2(__579__),
    .I1(__571__),
    .I0(__547__),
    .O(__604__)
  );
  LUT5 #(
    .INIT(32'h0001ffff)
  ) __1976__ (
    .I4(__532__),
    .I3(__537__),
    .I2(__536__),
    .I1(__535__),
    .I0(__534__),
    .O(__605__)
  );
  LUT5 #(
    .INIT(32'h0001ffff)
  ) __1977__ (
    .I4(__538__),
    .I3(__536__),
    .I2(__535__),
    .I1(__544__),
    .I0(__543__),
    .O(__606__)
  );
  LUT6 #(
    .INIT(64'h0000000080000000)
  ) __1978__ (
    .I5(__546__),
    .I4(__542__),
    .I3(__540__),
    .I2(__606__),
    .I1(__605__),
    .I0(__533__),
    .O(__607__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __1979__ (
    .I2(__536__),
    .I1(__538__),
    .I0(__109__),
    .O(__608__)
  );
  LUT5 #(
    .INIT(32'hf0880000)
  ) __1980__ (
    .I4(__532__),
    .I3(__536__),
    .I2(__271__),
    .I1(__537__),
    .I0(__435__),
    .O(__609__)
  );
  LUT5 #(
    .INIT(32'hf0880000)
  ) __1981__ (
    .I4(__532__),
    .I3(__534__),
    .I2(__131__),
    .I1(__535__),
    .I0(__66__),
    .O(__610__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __1982__ (
    .I2(__541__),
    .I1(__535__),
    .I0(g910),
    .O(__611__)
  );
  LUT6 #(
    .INIT(64'h0000000100000003)
  ) __1983__ (
    .I5(__581__),
    .I4(__611__),
    .I3(__610__),
    .I2(__609__),
    .I1(__608__),
    .I0(__229__),
    .O(__612__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __1984__ (
    .I2(__541__),
    .I1(__536__),
    .I0(__384__),
    .O(__613__)
  );
  LUT5 #(
    .INIT(32'h335f3333)
  ) __1985__ (
    .I4(g48),
    .I3(g31),
    .I2(__531__),
    .I1(__19__),
    .I0(__195__),
    .O(__614__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __1986__ (
    .I2(__538__),
    .I1(__543__),
    .I0(__190__),
    .O(__615__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __1987__ (
    .I2(__535__),
    .I1(__538__),
    .I0(g1182),
    .O(__616__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __1988__ (
    .I2(__538__),
    .I1(__544__),
    .I0(__209__),
    .O(__617__)
  );
  LUT6 #(
    .INIT(64'hca00000000000000)
  ) __1989__ (
    .I5(__532__),
    .I4(__577__),
    .I3(__576__),
    .I2(g42),
    .I1(__230__),
    .I0(__238__),
    .O(__618__)
  );
  LUT6 #(
    .INIT(64'h0000000000000004)
  ) __1990__ (
    .I5(__618__),
    .I4(__617__),
    .I3(__616__),
    .I2(__615__),
    .I1(__614__),
    .I0(__613__),
    .O(__619__)
  );
  LUT5 #(
    .INIT(32'h40ffbf00)
  ) __1991__ (
    .I4(__124__),
    .I3(g109),
    .I2(__619__),
    .I1(__612__),
    .I0(__607__),
    .O(__620__)
  );
  LUT5 #(
    .INIT(32'h0777ffff)
  ) __1992__ (
    .I4(__538__),
    .I3(__535__),
    .I2(g1170),
    .I1(__534__),
    .I0(g1194),
    .O(__621__)
  );
  LUT6 #(
    .INIT(64'h07770000ffff0000)
  ) __1993__ (
    .I5(__538__),
    .I4(__621__),
    .I3(__537__),
    .I2(__336__),
    .I1(__536__),
    .I0(__202__),
    .O(__622__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __1994__ (
    .I2(__532__),
    .I1(__535__),
    .I0(__80__),
    .O(__623__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __1995__ (
    .I2(__541__),
    .I1(__534__),
    .I0(g922),
    .O(__624__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __1996__ (
    .I2(__532__),
    .I1(__537__),
    .I0(__159__),
    .O(__625__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __1997__ (
    .I1(g48),
    .I0(g31),
    .O(__626__)
  );
  LUT6 #(
    .INIT(64'h0000000500000003)
  ) __1998__ (
    .I5(__626__),
    .I4(__625__),
    .I3(__624__),
    .I2(__623__),
    .I1(__140__),
    .I0(__546__),
    .O(__627__)
  );
  LUT3 #(
    .INIT(8'h35)
  ) __1999__ (
    .I2(g42),
    .I1(__442__),
    .I0(__93__),
    .O(__628__)
  );
  LUT6 #(
    .INIT(64'h00bfbfbfbfbfbfbf)
  ) __2000__ (
    .I5(__538__),
    .I4(__544__),
    .I3(__199__),
    .I2(__532__),
    .I1(__552__),
    .I0(__628__),
    .O(__629__)
  );
  LUT6 #(
    .INIT(64'h007f7f7f7f7f7f7f)
  ) __2001__ (
    .I5(__541__),
    .I4(__536__),
    .I3(__467__),
    .I2(__538__),
    .I1(__543__),
    .I0(__481__),
    .O(__630__)
  );
  LUT6 #(
    .INIT(64'h007f7f7f7f7f7f7f)
  ) __2002__ (
    .I5(__532__),
    .I4(__531__),
    .I3(__276__),
    .I2(__541__),
    .I1(__535__),
    .I0(g898),
    .O(__631__)
  );
  LUT6 #(
    .INIT(64'h007f7f7f7f7f7f7f)
  ) __2003__ (
    .I5(__532__),
    .I4(__536__),
    .I3(__100__),
    .I2(__537__),
    .I1(__541__),
    .I0(__39__),
    .O(__632__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __2004__ (
    .I1(g45),
    .I0(g44),
    .O(__633__)
  );
  LUT6 #(
    .INIT(64'h007f7f7fffffffff)
  ) __2005__ (
    .I5(__541__),
    .I4(__554__),
    .I3(__247__),
    .I2(__556__),
    .I1(__633__),
    .I0(g886),
    .O(__634__)
  );
  LUT5 #(
    .INIT(32'h0777ffff)
  ) __2006__ (
    .I4(__532__),
    .I3(__534__),
    .I2(__236__),
    .I1(__530__),
    .I0(__495__),
    .O(__635__)
  );
  LUT6 #(
    .INIT(64'h8000000000000000)
  ) __2007__ (
    .I5(__635__),
    .I4(__634__),
    .I3(__632__),
    .I2(__631__),
    .I1(__630__),
    .I0(__629__),
    .O(__636__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __2008__ (
    .I1(__394__),
    .I0(__301__),
    .O(__637__)
  );
  LUT6 #(
    .INIT(64'h00000000bfff0000)
  ) __2009__ (
    .I5(__637__),
    .I4(g109),
    .I3(__636__),
    .I2(__627__),
    .I1(__622__),
    .I0(__547__),
    .O(__638__)
  );
  LUT5 #(
    .INIT(32'h00008000)
  ) __2010__ (
    .I4(__546__),
    .I3(__542__),
    .I2(__540__),
    .I1(__606__),
    .I0(__605__),
    .O(__639__)
  );
  LUT6 #(
    .INIT(64'h0000000010000000)
  ) __2011__ (
    .I5(g42),
    .I4(g48),
    .I3(g45),
    .I2(__541__),
    .I1(g44),
    .I0(g43),
    .O(__640__)
  );
  LUT6 #(
    .INIT(64'h0000000010000000)
  ) __2012__ (
    .I5(g42),
    .I4(g48),
    .I3(g45),
    .I2(__538__),
    .I1(g44),
    .I0(g43),
    .O(__641__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __2013__ (
    .I5(__370__),
    .I4(__641__),
    .I3(__600__),
    .I2(g1185),
    .I1(__126__),
    .I0(__640__),
    .O(__642__)
  );
  LUT6 #(
    .INIT(64'h0000000080000000)
  ) __2014__ (
    .I5(g42),
    .I4(g48),
    .I3(g44),
    .I2(g45),
    .I1(g43),
    .I0(__538__),
    .O(__643__)
  );
  LUT6 #(
    .INIT(64'h0000000080000000)
  ) __2015__ (
    .I5(g45),
    .I4(g48),
    .I3(g42),
    .I2(g44),
    .I1(g43),
    .I0(__541__),
    .O(__644__)
  );
  LUT3 #(
    .INIT(8'hb0)
  ) __2016__ (
    .I2(__432__),
    .I1(g48),
    .I0(g31),
    .O(__645__)
  );
  LUT5 #(
    .INIT(32'hca000000)
  ) __2017__ (
    .I4(__532__),
    .I3(__552__),
    .I2(g42),
    .I1(__359__),
    .I0(__482__),
    .O(__646__)
  );
  LUT6 #(
    .INIT(64'h000000000000153f)
  ) __2018__ (
    .I5(__646__),
    .I4(__645__),
    .I3(__644__),
    .I2(__643__),
    .I1(__285__),
    .I0(g913),
    .O(__647__)
  );
  LUT5 #(
    .INIT(32'hf0880000)
  ) __2019__ (
    .I4(__532__),
    .I3(__536__),
    .I2(__78__),
    .I1(__537__),
    .I0(__62__),
    .O(__648__)
  );
  LUT6 #(
    .INIT(64'h000f007700ff00ff)
  ) __2020__ (
    .I5(__532__),
    .I4(__534__),
    .I3(__648__),
    .I2(__178__),
    .I1(__535__),
    .I0(__306__),
    .O(__649__)
  );
  LUT6 #(
    .INIT(64'h4000ffffbfff0000)
  ) __2021__ (
    .I5(__484__),
    .I4(g109),
    .I3(__649__),
    .I2(__647__),
    .I1(__642__),
    .I0(__639__),
    .O(__650__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __2022__ (
    .I1(__394__),
    .I0(__301__),
    .O(__651__)
  );
  LUT6 #(
    .INIT(64'h000000004000ffff)
  ) __2023__ (
    .I5(__651__),
    .I4(g109),
    .I3(__636__),
    .I2(__627__),
    .I1(__622__),
    .I0(__547__),
    .O(__652__)
  );
  LUT5 #(
    .INIT(32'h00f70000)
  ) __2024__ (
    .I4(g109),
    .I3(__21__),
    .I2(__547__),
    .I1(__564__),
    .I0(__559__),
    .O(__653__)
  );
  LUT6 #(
    .INIT(64'h0000000000000001)
  ) __2025__ (
    .I5(__653__),
    .I4(__652__),
    .I3(__650__),
    .I2(__638__),
    .I1(__620__),
    .I0(__604__),
    .O(__654__)
  );
  LUT6 #(
    .INIT(64'h8000000000000000)
  ) __2026__ (
    .I5(g48),
    .I4(g42),
    .I3(g44),
    .I2(g45),
    .I1(g43),
    .I0(__538__),
    .O(__655__)
  );
  LUT6 #(
    .INIT(64'h000f000f000f11ff)
  ) __2027__ (
    .I5(__537__),
    .I4(__535__),
    .I3(__532__),
    .I2(__538__),
    .I1(__536__),
    .I0(__534__),
    .O(__656__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __2028__ (
    .I2(__532__),
    .I1(__535__),
    .I0(__193__),
    .O(__657__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __2029__ (
    .I2(__532__),
    .I1(__537__),
    .I0(__167__),
    .O(__658__)
  );
  LUT6 #(
    .INIT(64'h007f7f7f7f7f7f7f)
  ) __2030__ (
    .I5(__537__),
    .I4(__541__),
    .I3(__401__),
    .I2(__535__),
    .I1(__538__),
    .I0(g1191),
    .O(__659__)
  );
  LUT6 #(
    .INIT(64'h007f7f7f7f7f7f7f)
  ) __2031__ (
    .I5(__537__),
    .I4(__538__),
    .I3(__122__),
    .I2(__541__),
    .I1(__535__),
    .I0(g919),
    .O(__660__)
  );
  LUT5 #(
    .INIT(32'h335f3333)
  ) __2032__ (
    .I4(g48),
    .I3(g31),
    .I2(__544__),
    .I1(__187__),
    .I0(__177__),
    .O(__661__)
  );
  LUT4 #(
    .INIT(16'h8000)
  ) __2033__ (
    .I3(__532__),
    .I2(g42),
    .I1(__552__),
    .I0(__310__),
    .O(__662__)
  );
  LUT6 #(
    .INIT(64'h0000000010000000)
  ) __2034__ (
    .I5(__662__),
    .I4(__661__),
    .I3(__660__),
    .I2(__659__),
    .I1(__658__),
    .I0(__657__),
    .O(__663__)
  );
  LUT6 #(
    .INIT(64'h10000000ffffffff)
  ) __2035__ (
    .I5(__663__),
    .I4(__656__),
    .I3(__542__),
    .I2(__540__),
    .I1(__655__),
    .I0(__546__),
    .O(__664__)
  );
  LUT4 #(
    .INIT(16'h8000)
  ) __2036__ (
    .I3(__656__),
    .I2(__545__),
    .I1(__542__),
    .I0(__540__),
    .O(__665__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __2037__ (
    .I1(g1188),
    .I0(__600__),
    .O(__666__)
  );
  LUT3 #(
    .INIT(8'h75)
  ) __2038__ (
    .I2(g48),
    .I1(g31),
    .I0(__428__),
    .O(__667__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __2039__ (
    .I2(__536__),
    .I1(__538__),
    .I0(__160__),
    .O(__668__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __2040__ (
    .I2(__537__),
    .I1(__417__),
    .I0(__538__),
    .O(__669__)
  );
  LUT6 #(
    .INIT(64'h000000000000153f)
  ) __2041__ (
    .I5(__669__),
    .I4(__668__),
    .I3(__409__),
    .I2(__147__),
    .I1(__655__),
    .I0(__643__),
    .O(__670__)
  );
  LUT3 #(
    .INIT(8'h1f)
  ) __2042__ (
    .I2(__532__),
    .I1(__535__),
    .I0(__534__),
    .O(__671__)
  );
  LUT5 #(
    .INIT(32'h0777ffff)
  ) __2043__ (
    .I4(__541__),
    .I3(__537__),
    .I2(__462__),
    .I1(__18__),
    .I0(__536__),
    .O(__672__)
  );
  LUT6 #(
    .INIT(64'h00efefef00000000)
  ) __2044__ (
    .I5(__672__),
    .I4(g916),
    .I3(__644__),
    .I2(__375__),
    .I1(__534__),
    .I0(__671__),
    .O(__673__)
  );
  LUT6 #(
    .INIT(64'h3b7f7f7f7f7f7f7f)
  ) __2045__ (
    .I5(g42),
    .I4(__577__),
    .I3(__172__),
    .I2(__4__),
    .I1(__532__),
    .I0(__537__),
    .O(__674__)
  );
  LUT6 #(
    .INIT(64'hefffffffffffffff)
  ) __2046__ (
    .I5(__674__),
    .I4(__673__),
    .I3(__670__),
    .I2(__667__),
    .I1(__666__),
    .I0(__665__),
    .O(__675__)
  );
  LUT5 #(
    .INIT(32'h8040201f)
  ) __2047__ (
    .I4(__169__),
    .I3(__485__),
    .I2(g109),
    .I1(__675__),
    .I0(__664__),
    .O(__676__)
  );
  LUT3 #(
    .INIT(8'h01)
  ) __2048__ (
    .I2(__484__),
    .I1(__169__),
    .I0(__28__),
    .O(__677__)
  );
  LUT6 #(
    .INIT(64'h0000000000000040)
  ) __2049__ (
    .I5(__485__),
    .I4(__299__),
    .I3(__21__),
    .I2(__677__),
    .I1(__651__),
    .I0(__124__),
    .O(__678__)
  );
  LUT4 #(
    .INIT(16'h7f00)
  ) __2050__ (
    .I3(__678__),
    .I2(__676__),
    .I1(__654__),
    .I0(__603__),
    .O(__679__)
  );
  LUT5 #(
    .INIT(32'h00d70000)
  ) __2051__ (
    .I4(__528__),
    .I3(__679__),
    .I2(__340__),
    .I1(__529__),
    .I0(__524__),
    .O(__680__)
  );
  LUT6 #(
    .INIT(64'hff00f870ff00ff00)
  ) __2052__ (
    .I5(__680__),
    .I4(__519__),
    .I3(__467__),
    .I2(__28__),
    .I1(g109),
    .I0(__380__),
    .O(__681__)
  );
  LUT6 #(
    .INIT(64'h0a0a0a0a060a0a0a)
  ) __2053__ (
    .I5(__11__),
    .I4(g1696),
    .I3(__53__),
    .I2(__154__),
    .I1(__226__),
    .I0(__145__),
    .O(__682__)
  );
  LUT6 #(
    .INIT(64'h8000000000000000)
  ) __2054__ (
    .I5(__405__),
    .I4(__445__),
    .I3(__456__),
    .I2(__237__),
    .I1(__453__),
    .I0(__214__),
    .O(__683__)
  );
  LUT4 #(
    .INIT(16'h0060)
  ) __2055__ (
    .I3(__407__),
    .I2(g109),
    .I1(__497__),
    .I0(__683__),
    .O(__684__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __2056__ (
    .I1(__32__),
    .I0(__12__),
    .O(__685__)
  );
  LUT4 #(
    .INIT(16'h0004)
  ) __2057__ (
    .I3(__166__),
    .I2(__437__),
    .I1(__357__),
    .I0(__216__),
    .O(__686__)
  );
  LUT6 #(
    .INIT(64'h0000ffffa0a03fff)
  ) __2058__ (
    .I5(__345__),
    .I4(__478__),
    .I3(__37__),
    .I2(__686__),
    .I1(__685__),
    .I0(__491__),
    .O(__687__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __2059__ (
    .I1(g18),
    .I0(__687__),
    .O(__688__)
  );
  LUT6 #(
    .INIT(64'hb00b00000000b00b)
  ) __2060__ (
    .I5(__365__),
    .I4(__23__),
    .I3(__255__),
    .I2(__293__),
    .I1(__334__),
    .I0(__186__),
    .O(__689__)
  );
  LUT4 #(
    .INIT(16'h9009)
  ) __2061__ (
    .I3(__355__),
    .I2(__250__),
    .I1(__326__),
    .I0(__206__),
    .O(__690__)
  );
  LUT2 #(
    .INIT(4'h9)
  ) __2062__ (
    .I1(__68__),
    .I0(__219__),
    .O(__691__)
  );
  LUT6 #(
    .INIT(64'h9009000000000000)
  ) __2063__ (
    .I5(__691__),
    .I4(__690__),
    .I3(__179__),
    .I2(__260__),
    .I1(__85__),
    .I0(__141__),
    .O(__692__)
  );
  LUT6 #(
    .INIT(64'hb00b000000000000)
  ) __2064__ (
    .I5(__692__),
    .I4(__689__),
    .I3(__95__),
    .I2(__251__),
    .I1(__186__),
    .I0(__334__),
    .O(__693__)
  );
  LUT6 #(
    .INIT(64'h0000000000000040)
  ) __2065__ (
    .I5(g48),
    .I4(g44),
    .I3(g45),
    .I2(__532__),
    .I1(g42),
    .I0(g43),
    .O(__694__)
  );
  LUT3 #(
    .INIT(8'he0)
  ) __2066__ (
    .I2(__463__),
    .I1(__694__),
    .I0(__675__),
    .O(__695__)
  );
  LUT6 #(
    .INIT(64'h0000000000000001)
  ) __2067__ (
    .I5(__95__),
    .I4(__317__),
    .I3(__326__),
    .I2(__365__),
    .I1(__334__),
    .I0(__179__),
    .O(__696__)
  );
  LUT3 #(
    .INIT(8'h01)
  ) __2068__ (
    .I2(__377__),
    .I1(__68__),
    .I0(__355__),
    .O(__697__)
  );
  LUT6 #(
    .INIT(64'h0000000000000040)
  ) __2069__ (
    .I5(__396__),
    .I4(__85__),
    .I3(__232__),
    .I2(__697__),
    .I1(__696__),
    .I0(__255__),
    .O(__698__)
  );
  LUT4 #(
    .INIT(16'h8000)
  ) __2070__ (
    .I3(__201__),
    .I2(__98__),
    .I1(__14__),
    .I0(__411__),
    .O(__699__)
  );
  LUT4 #(
    .INIT(16'h3e00)
  ) __2071__ (
    .I3(__699__),
    .I2(__406__),
    .I1(__71__),
    .I0(__698__),
    .O(__700__)
  );
  LUT6 #(
    .INIT(64'hd77d000000000000)
  ) __2072__ (
    .I5(__508__),
    .I4(__699__),
    .I3(__314__),
    .I2(__700__),
    .I1(__695__),
    .I0(__693__),
    .O(__701__)
  );
  LUT5 #(
    .INIT(32'hdfdd0000)
  ) __2073__ (
    .I4(g109),
    .I3(__106__),
    .I2(__170__),
    .I1(__320__),
    .I0(__433__),
    .O(__702__)
  );
  LUT5 #(
    .INIT(32'h7f800000)
  ) __2074__ (
    .I4(__702__),
    .I3(__427__),
    .I2(__701__),
    .I1(__469__),
    .I0(__336__),
    .O(__703__)
  );
  LUT6 #(
    .INIT(64'h0caa0c0c0c0c0c0c)
  ) __2075__ (
    .I5(__56__),
    .I4(__512__),
    .I3(__295__),
    .I2(__511__),
    .I1(__45__),
    .I0(__51__),
    .O(__704__)
  );
  LUT4 #(
    .INIT(16'hccca)
  ) __2076__ (
    .I3(__11__),
    .I2(g1696),
    .I1(__250__),
    .I0(__207__),
    .O(__705__)
  );
  LUT6 #(
    .INIT(64'hff00f870ff00ff00)
  ) __2077__ (
    .I5(__680__),
    .I4(__519__),
    .I3(__223__),
    .I2(__484__),
    .I1(g109),
    .I0(__380__),
    .O(__706__)
  );
  LUT6 #(
    .INIT(64'h0000000000000001)
  ) __2078__ (
    .I5(__6__),
    .I4(__91__),
    .I3(__267__),
    .I2(__346__),
    .I1(__423__),
    .I0(__102__),
    .O(__707__)
  );
  LUT3 #(
    .INIT(8'h01)
  ) __2079__ (
    .I2(__449__),
    .I1(__96__),
    .I0(__335__),
    .O(__708__)
  );
  LUT6 #(
    .INIT(64'h0000000000000040)
  ) __2080__ (
    .I5(__10__),
    .I4(__339__),
    .I3(__157__),
    .I2(__708__),
    .I1(__707__),
    .I0(__450__),
    .O(__709__)
  );
  LUT6 #(
    .INIT(64'hff003e3e00003e3e)
  ) __2081__ (
    .I5(g109),
    .I4(__679__),
    .I3(__339__),
    .I2(__55__),
    .I1(__341__),
    .I0(__709__),
    .O(__710__)
  );
  LUT6 #(
    .INIT(64'h0000008080808000)
  ) __2082__ (
    .I5(__414__),
    .I4(__112__),
    .I3(__273__),
    .I2(__362__),
    .I1(__176__),
    .I0(__67__),
    .O(__711__)
  );
  LUT6 #(
    .INIT(64'h8000000000000000)
  ) __2083__ (
    .I5(__120__),
    .I4(__472__),
    .I3(__77__),
    .I2(__328__),
    .I1(__490__),
    .I0(__711__),
    .O(__712__)
  );
  LUT6 #(
    .INIT(64'h00000000000000e1)
  ) __2084__ (
    .I5(__362__),
    .I4(__176__),
    .I3(__67__),
    .I2(__414__),
    .I1(__112__),
    .I0(__273__),
    .O(__713__)
  );
  LUT6 #(
    .INIT(64'h0000000000000004)
  ) __2085__ (
    .I5(__120__),
    .I4(__472__),
    .I3(__77__),
    .I2(__328__),
    .I1(__713__),
    .I0(__490__),
    .O(__714__)
  );
  LUT3 #(
    .INIT(8'h08)
  ) __2086__ (
    .I2(__56__),
    .I1(__295__),
    .I0(__273__),
    .O(__715__)
  );
  LUT4 #(
    .INIT(16'h0004)
  ) __2087__ (
    .I3(__333__),
    .I2(__309__),
    .I1(__118__),
    .I0(__261__),
    .O(__716__)
  );
  LUT6 #(
    .INIT(64'h00000000fef00000)
  ) __2088__ (
    .I5(__269__),
    .I4(__716__),
    .I3(__292__),
    .I2(__715__),
    .I1(__414__),
    .I0(__112__),
    .O(__717__)
  );
  LUT4 #(
    .INIT(16'hac00)
  ) __2089__ (
    .I3(__717__),
    .I2(__17__),
    .I1(__714__),
    .I0(__712__),
    .O(__718__)
  );
  LUT6 #(
    .INIT(64'h80c088ccc0c00c00)
  ) __2090__ (
    .I5(__273__),
    .I4(__414__),
    .I3(__295__),
    .I2(__112__),
    .I1(__718__),
    .I0(__56__),
    .O(__719__)
  );
  LUT3 #(
    .INIT(8'h01)
  ) __2091__ (
    .I2(__295__),
    .I1(__414__),
    .I0(__112__),
    .O(__720__)
  );
  LUT6 #(
    .INIT(64'h0000eeee0eeeeeee)
  ) __2092__ (
    .I5(__56__),
    .I4(__512__),
    .I3(__720__),
    .I2(__273__),
    .I1(__713__),
    .I0(__711__),
    .O(__721__)
  );
  LUT6 #(
    .INIT(64'h00000000aa008000)
  ) __2093__ (
    .I5(__269__),
    .I4(__56__),
    .I3(__716__),
    .I2(__720__),
    .I1(__273__),
    .I0(__51__),
    .O(__722__)
  );
  LUT6 #(
    .INIT(64'h0000fffffffdffff)
  ) __2094__ (
    .I5(__56__),
    .I4(__512__),
    .I3(__295__),
    .I2(__414__),
    .I1(__112__),
    .I0(__273__),
    .O(__723__)
  );
  LUT6 #(
    .INIT(64'h02020222aaaaaaaa)
  ) __2095__ (
    .I5(__512__),
    .I4(__414__),
    .I3(__112__),
    .I2(__292__),
    .I1(__715__),
    .I0(__723__),
    .O(__724__)
  );
  LUT5 #(
    .INIT(32'h000053ff)
  ) __2096__ (
    .I4(__511__),
    .I3(__717__),
    .I2(__17__),
    .I1(__714__),
    .I0(__712__),
    .O(__725__)
  );
  LUT6 #(
    .INIT(64'hffabaafeaaaaaaaa)
  ) __2097__ (
    .I5(__725__),
    .I4(__120__),
    .I3(__724__),
    .I2(__722__),
    .I1(__721__),
    .I0(__719__),
    .O(__726__)
  );
  LUT2 #(
    .INIT(4'he)
  ) __2098__ (
    .I1(__433__),
    .I0(__5__),
    .O(__727__)
  );
  LUT6 #(
    .INIT(64'h00000000000000e1)
  ) __2099__ (
    .I5(__60__),
    .I4(__110__),
    .I3(__503__),
    .I2(__32__),
    .I1(__37__),
    .I0(__12__),
    .O(__728__)
  );
  LUT6 #(
    .INIT(64'h0000000000000004)
  ) __2100__ (
    .I5(__479__),
    .I4(__327__),
    .I3(__363__),
    .I2(__189__),
    .I1(__728__),
    .I0(__33__),
    .O(__729__)
  );
  LUT6 #(
    .INIT(64'h0000008080808000)
  ) __2101__ (
    .I5(__32__),
    .I4(__37__),
    .I3(__12__),
    .I2(__60__),
    .I1(__110__),
    .I0(__503__),
    .O(__730__)
  );
  LUT6 #(
    .INIT(64'h8000000000000000)
  ) __2102__ (
    .I5(__479__),
    .I4(__327__),
    .I3(__363__),
    .I2(__189__),
    .I1(__33__),
    .I0(__730__),
    .O(__731__)
  );
  LUT6 #(
    .INIT(64'hbf0fbfbfbfbfbfbf)
  ) __2103__ (
    .I5(__37__),
    .I4(__345__),
    .I3(__478__),
    .I2(__686__),
    .I1(__429__),
    .I0(__685__),
    .O(__732__)
  );
  LUT4 #(
    .INIT(16'h00ca)
  ) __2104__ (
    .I3(__732__),
    .I2(__192__),
    .I1(__731__),
    .I0(__729__),
    .O(__733__)
  );
  LUT5 #(
    .INIT(32'h33ff337f)
  ) __2105__ (
    .I4(__733__),
    .I3(__478__),
    .I2(__37__),
    .I1(__686__),
    .I0(__345__),
    .O(__734__)
  );
  LUT6 #(
    .INIT(64'hf0f0e2e2f0f022e2)
  ) __2106__ (
    .I5(__37__),
    .I4(__345__),
    .I3(__685__),
    .I2(__493__),
    .I1(__734__),
    .I0(__125__),
    .O(__735__)
  );
  LUT4 #(
    .INIT(16'h00cd)
  ) __2107__ (
    .I3(__273__),
    .I2(__414__),
    .I1(__295__),
    .I0(__112__),
    .O(__736__)
  );
  LUT4 #(
    .INIT(16'hbf80)
  ) __2108__ (
    .I3(__426__),
    .I2(__393__),
    .I1(__701__),
    .I0(__116__),
    .O(__737__)
  );
  LUT4 #(
    .INIT(16'hf088)
  ) __2109__ (
    .I3(__508__),
    .I2(__179__),
    .I1(g109),
    .I0(__95__),
    .O(__738__)
  );
  LUT3 #(
    .INIT(8'hf4)
  ) __2110__ (
    .I2(__228__),
    .I1(g750),
    .I0(__438__),
    .O(__739__)
  );
  LUT4 #(
    .INIT(16'hbf80)
  ) __2111__ (
    .I3(__122__),
    .I2(__393__),
    .I1(__701__),
    .I0(__53__),
    .O(__740__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __2112__ (
    .I1(g109),
    .I0(__252__),
    .O(__741__)
  );
  LUT4 #(
    .INIT(16'hebee)
  ) __2113__ (
    .I3(g1696),
    .I2(__11__),
    .I1(__226__),
    .I0(__154__),
    .O(__742__)
  );
  LUT6 #(
    .INIT(64'h7fff800000000000)
  ) __2114__ (
    .I5(__702__),
    .I4(__90__),
    .I3(__701__),
    .I2(__469__),
    .I1(__336__),
    .I0(__427__),
    .O(__743__)
  );
  LUT4 #(
    .INIT(16'hf088)
  ) __2115__ (
    .I3(__508__),
    .I2(__377__),
    .I1(g109),
    .I0(__71__),
    .O(__744__)
  );
  LUT6 #(
    .INIT(64'hfffffffffdffffff)
  ) __2116__ (
    .I5(__547__),
    .I4(__562__),
    .I3(__561__),
    .I2(__563__),
    .I1(__560__),
    .I0(__559__),
    .O(__745__)
  );
  LUT3 #(
    .INIT(8'h35)
  ) __2117__ (
    .I2(g18),
    .I1(__494__),
    .I0(__283__),
    .O(__746__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __2118__ (
    .I1(__11__),
    .I0(g1696),
    .O(__747__)
  );
  LUT6 #(
    .INIT(64'hff00bb00ff000f00)
  ) __2119__ (
    .I5(__73__),
    .I4(__211__),
    .I3(__747__),
    .I2(__746__),
    .I1(g109),
    .I0(__745__),
    .O(__748__)
  );
  LUT4 #(
    .INIT(16'heeec)
  ) __2120__ (
    .I3(__11__),
    .I2(g1696),
    .I1(__748__),
    .I0(__434__),
    .O(__749__)
  );
  LUT6 #(
    .INIT(64'h5500005455005500)
  ) __2121__ (
    .I5(__118__),
    .I4(__333__),
    .I3(__309__),
    .I2(__261__),
    .I1(__269__),
    .I0(__511__),
    .O(__750__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __2122__ (
    .I1(g109),
    .I0(__128__),
    .O(__751__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __2123__ (
    .I1(g109),
    .I0(__308__),
    .O(__752__)
  );
  LUT4 #(
    .INIT(16'h88f0)
  ) __2124__ (
    .I3(__679__),
    .I2(__399__),
    .I1(g109),
    .I0(__361__),
    .O(__753__)
  );
  LUT5 #(
    .INIT(32'h00007800)
  ) __2125__ (
    .I4(__407__),
    .I3(g109),
    .I2(__237__),
    .I1(__453__),
    .I0(__214__),
    .O(__754__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __2126__ (
    .I1(__279__),
    .I0(__222__),
    .O(__755__)
  );
  LUT6 #(
    .INIT(64'h555555553000cfff)
  ) __2127__ (
    .I5(g18),
    .I4(__81__),
    .I3(__149__),
    .I2(__755__),
    .I1(__400__),
    .I0(__225__),
    .O(__756__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __2128__ (
    .I2(g109),
    .I1(__756__),
    .I0(__163__),
    .O(__757__)
  );
  LUT4 #(
    .INIT(16'h8000)
  ) __2129__ (
    .I3(__458__),
    .I2(__39__),
    .I1(__344__),
    .I0(__404__),
    .O(__758__)
  );
  LUT4 #(
    .INIT(16'h0080)
  ) __2130__ (
    .I3(__607__),
    .I2(g109),
    .I1(__619__),
    .I0(__612__),
    .O(__759__)
  );
  LUT3 #(
    .INIT(8'h35)
  ) __2131__ (
    .I2(g18),
    .I1(__174__),
    .I0(__374__),
    .O(__760__)
  );
  LUT6 #(
    .INIT(64'h0033000faaaaaaaa)
  ) __2132__ (
    .I5(__747__),
    .I4(__73__),
    .I3(__211__),
    .I2(__760__),
    .I1(__759__),
    .I0(__286__),
    .O(__761__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __2133__ (
    .I2(g109),
    .I1(__278__),
    .I0(__196__),
    .O(__762__)
  );
  LUT5 #(
    .INIT(32'h7f800000)
  ) __2134__ (
    .I4(__762__),
    .I3(__182__),
    .I2(__439__),
    .I1(__500__),
    .I0(__200__),
    .O(__763__)
  );
  LUT2 #(
    .INIT(4'he)
  ) __2135__ (
    .I1(g82),
    .I0(__353__),
    .O(__764__)
  );
  LUT6 #(
    .INIT(64'hfbfa000000000000)
  ) __2136__ (
    .I5(g109),
    .I4(__465__),
    .I3(__489__),
    .I2(g881),
    .I1(__198__),
    .I0(__245__),
    .O(__765__)
  );
  LUT4 #(
    .INIT(16'h88f0)
  ) __2137__ (
    .I3(__679__),
    .I2(__335__),
    .I1(g109),
    .I0(__450__),
    .O(__766__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __2138__ (
    .I1(__279__),
    .I0(__222__),
    .O(__767__)
  );
  LUT6 #(
    .INIT(64'hcfff3000aaaaaaaa)
  ) __2139__ (
    .I5(__747__),
    .I4(__308__),
    .I3(__400__),
    .I2(__767__),
    .I1(__149__),
    .I0(__283__),
    .O(__768__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __2140__ (
    .I1(g109),
    .I0(__217__),
    .O(__769__)
  );
  LUT4 #(
    .INIT(16'hbfff)
  ) __2141__ (
    .I3(__649__),
    .I2(__647__),
    .I1(__642__),
    .I0(__639__),
    .O(__770__)
  );
  LUT6 #(
    .INIT(64'h40bfbf40bf4040bf)
  ) __2142__ (
    .I5(__675__),
    .I4(__770__),
    .I3(__664__),
    .I2(__619__),
    .I1(__612__),
    .I0(__607__),
    .O(__771__)
  );
  LUT5 #(
    .INIT(32'hbfffffff)
  ) __2143__ (
    .I4(__601__),
    .I3(__595__),
    .I2(__590__),
    .I1(__588__),
    .I0(__547__),
    .O(__772__)
  );
  LUT4 #(
    .INIT(16'hbfff)
  ) __2144__ (
    .I3(__636__),
    .I2(__627__),
    .I1(__622__),
    .I0(__547__),
    .O(__773__)
  );
  LUT4 #(
    .INIT(16'hbfff)
  ) __2145__ (
    .I3(__584__),
    .I2(__579__),
    .I1(__571__),
    .I0(__547__),
    .O(__774__)
  );
  LUT3 #(
    .INIT(8'h0d)
  ) __2146__ (
    .I2(__253__),
    .I1(g31),
    .I0(g48),
    .O(__775__)
  );
  LUT6 #(
    .INIT(64'h9669699669969669)
  ) __2147__ (
    .I5(__745__),
    .I4(__775__),
    .I3(__774__),
    .I2(__773__),
    .I1(__772__),
    .I0(__771__),
    .O(__776__)
  );
  LUT5 #(
    .INIT(32'hfffeffff)
  ) __2148__ (
    .I4(g48),
    .I3(g41),
    .I2(g30),
    .I1(g31),
    .I0(__776__),
    .O(__777__)
  );
  LUT6 #(
    .INIT(64'hff00bf80aaaaaaaa)
  ) __2149__ (
    .I5(g109),
    .I4(__276__),
    .I3(__93__),
    .I2(g18),
    .I1(__212__),
    .I0(__34__),
    .O(__778__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __2150__ (
    .I1(g109),
    .I0(__63__),
    .O(__779__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __2151__ (
    .I1(__468__),
    .I0(__297__),
    .O(__780__)
  );
  LUT6 #(
    .INIT(64'h555555553000cfff)
  ) __2152__ (
    .I5(__679__),
    .I4(__6__),
    .I3(__156__),
    .I2(__780__),
    .I1(__61__),
    .I0(__501__),
    .O(__781__)
  );
  LUT4 #(
    .INIT(16'ha3aa)
  ) __2153__ (
    .I3(g750),
    .I2(__438__),
    .I1(__781__),
    .I0(__461__),
    .O(__782__)
  );
  LUT2 #(
    .INIT(4'he)
  ) __2154__ (
    .I1(g82),
    .I0(__254__),
    .O(__783__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __2155__ (
    .I1(__120__),
    .I0(__711__),
    .O(__784__)
  );
  LUT3 #(
    .INIT(8'he1)
  ) __2156__ (
    .I2(__414__),
    .I1(__112__),
    .I0(__273__),
    .O(__785__)
  );
  LUT5 #(
    .INIT(32'h00000004)
  ) __2157__ (
    .I4(__362__),
    .I3(__176__),
    .I2(__67__),
    .I1(__785__),
    .I0(__120__),
    .O(__786__)
  );
  LUT6 #(
    .INIT(64'haacc0000f0f0f0f0)
  ) __2158__ (
    .I5(__723__),
    .I4(__717__),
    .I3(__472__),
    .I2(__457__),
    .I1(__786__),
    .I0(__784__),
    .O(__787__)
  );
  LUT4 #(
    .INIT(16'hbeaa)
  ) __2159__ (
    .I3(__725__),
    .I2(__328__),
    .I1(__787__),
    .I0(__719__),
    .O(__788__)
  );
  LUT3 #(
    .INIT(8'h35)
  ) __2160__ (
    .I2(g18),
    .I1(__424__),
    .I0(__389__),
    .O(__789__)
  );
  LUT5 #(
    .INIT(32'h000044f0)
  ) __2161__ (
    .I4(__211__),
    .I3(__73__),
    .I2(__789__),
    .I1(g109),
    .I0(__773__),
    .O(__790__)
  );
  LUT4 #(
    .INIT(16'haaa3)
  ) __2162__ (
    .I3(__11__),
    .I2(g1696),
    .I1(__790__),
    .I0(__101__),
    .O(__791__)
  );
  LUT3 #(
    .INIT(8'h04)
  ) __2163__ (
    .I2(__166__),
    .I1(__357__),
    .I0(__437__),
    .O(__792__)
  );
  LUT6 #(
    .INIT(64'h0001ffffffff0001)
  ) __2164__ (
    .I5(__792__),
    .I4(__216__),
    .I3(__37__),
    .I2(__32__),
    .I1(__345__),
    .I0(__12__),
    .O(__793__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __2165__ (
    .I2(__47__),
    .I1(__413__),
    .I0(__270__),
    .O(__794__)
  );
  LUT5 #(
    .INIT(32'h53ac0000)
  ) __2166__ (
    .I4(g109),
    .I3(__376__),
    .I2(g18),
    .I1(__16__),
    .I0(__185__),
    .O(__795__)
  );
  LUT6 #(
    .INIT(64'hff00bf80aaaaaaaa)
  ) __2167__ (
    .I5(g109),
    .I4(__276__),
    .I3(__359__),
    .I2(g18),
    .I1(__212__),
    .I0(__466__),
    .O(__796__)
  );
  LUT5 #(
    .INIT(32'h80000000)
  ) __2168__ (
    .I4(__421__),
    .I3(__182__),
    .I2(__439__),
    .I1(__500__),
    .I0(__200__),
    .O(__797__)
  );
  LUT6 #(
    .INIT(64'h7fff800000000000)
  ) __2169__ (
    .I5(__762__),
    .I4(__367__),
    .I3(__235__),
    .I2(__398__),
    .I1(__266__),
    .I0(__797__),
    .O(__798__)
  );
  LUT5 #(
    .INIT(32'hdfdd0000)
  ) __2170__ (
    .I4(g109),
    .I3(__338__),
    .I2(__249__),
    .I1(__380__),
    .I0(__114__),
    .O(__799__)
  );
  LUT5 #(
    .INIT(32'h7f800000)
  ) __2171__ (
    .I4(__799__),
    .I3(__344__),
    .I2(__458__),
    .I1(__39__),
    .I0(__680__),
    .O(__800__)
  );
  LUT6 #(
    .INIT(64'h8088808888880000)
  ) __2172__ (
    .I5(__37__),
    .I4(__32__),
    .I3(__345__),
    .I2(__478__),
    .I1(__12__),
    .I0(__733__),
    .O(__801__)
  );
  LUT6 #(
    .INIT(64'h0000fffffffdffff)
  ) __2173__ (
    .I5(__478__),
    .I4(__686__),
    .I3(__32__),
    .I2(__345__),
    .I1(__12__),
    .I0(__37__),
    .O(__802__)
  );
  LUT5 #(
    .INIT(32'h00eef0f0)
  ) __2174__ (
    .I4(__802__),
    .I3(__732__),
    .I2(__491__),
    .I1(__729__),
    .I0(__731__),
    .O(__803__)
  );
  LUT4 #(
    .INIT(16'h0001)
  ) __2175__ (
    .I3(__37__),
    .I2(__32__),
    .I1(__345__),
    .I0(__12__),
    .O(__804__)
  );
  LUT5 #(
    .INIT(32'h0000f3f5)
  ) __2176__ (
    .I4(__804__),
    .I3(__192__),
    .I2(__732__),
    .I1(__731__),
    .I0(__729__),
    .O(__805__)
  );
  LUT4 #(
    .INIT(16'hbeaa)
  ) __2177__ (
    .I3(__805__),
    .I2(__192__),
    .I1(__803__),
    .I0(__801__),
    .O(__806__)
  );
  LUT6 #(
    .INIT(64'hcfff3000aaaaaaaa)
  ) __2178__ (
    .I5(__747__),
    .I4(__152__),
    .I3(__400__),
    .I2(__755__),
    .I1(__149__),
    .I0(__282__),
    .O(__807__)
  );
  LUT5 #(
    .INIT(32'h53ac0000)
  ) __2179__ (
    .I4(g109),
    .I3(__476__),
    .I2(g18),
    .I1(__142__),
    .I0(__392__),
    .O(__808__)
  );
  LUT6 #(
    .INIT(64'hff00bf80aaaaaaaa)
  ) __2180__ (
    .I5(g109),
    .I4(__276__),
    .I3(__46__),
    .I2(g18),
    .I1(__212__),
    .I0(__387__),
    .O(__809__)
  );
  LUT6 #(
    .INIT(64'hfafcfafafafafafa)
  ) __2181__ (
    .I5(__56__),
    .I4(__512__),
    .I3(__295__),
    .I2(__511__),
    .I1(__258__),
    .I0(__173__),
    .O(__810__)
  );
  LUT6 #(
    .INIT(64'h0000000000000001)
  ) __2182__ (
    .I5(__24__),
    .I4(__175__),
    .I3(__256__),
    .I2(__480__),
    .I1(__113__),
    .I0(__194__),
    .O(__811__)
  );
  LUT6 #(
    .INIT(64'h0000000000000001)
  ) __2183__ (
    .I5(__185__),
    .I4(__225__),
    .I3(__504__),
    .I2(__392__),
    .I1(__224__),
    .I0(__379__),
    .O(__812__)
  );
  LUT6 #(
    .INIT(64'h0000000000000040)
  ) __2184__ (
    .I5(__494__),
    .I4(__174__),
    .I3(__289__),
    .I2(__812__),
    .I1(__811__),
    .I0(__325__),
    .O(__813__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __2185__ (
    .I1(__302__),
    .I0(__415__),
    .O(__814__)
  );
  LUT6 #(
    .INIT(64'h0000000000000004)
  ) __2186__ (
    .I5(__44__),
    .I4(__424__),
    .I3(__288__),
    .I2(__155__),
    .I1(__814__),
    .I0(__252__),
    .O(__815__)
  );
  LUT4 #(
    .INIT(16'h8000)
  ) __2187__ (
    .I3(g109),
    .I2(__49__),
    .I1(__815__),
    .I0(__813__),
    .O(__816__)
  );
  LUT6 #(
    .INIT(64'h555555550300fcff)
  ) __2188__ (
    .I5(g18),
    .I4(__243__),
    .I3(__755__),
    .I2(__400__),
    .I1(__149__),
    .I0(__504__),
    .O(__817__)
  );
  LUT4 #(
    .INIT(16'haaa3)
  ) __2189__ (
    .I3(__11__),
    .I2(g1696),
    .I1(__817__),
    .I0(__448__),
    .O(__818__)
  );
  LUT6 #(
    .INIT(64'hff00bf80aaaaaaaa)
  ) __2190__ (
    .I5(g109),
    .I4(__15__),
    .I3(__447__),
    .I2(g18),
    .I1(__212__),
    .I0(__483__),
    .O(__819__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __2191__ (
    .I1(g109),
    .I0(__379__),
    .O(__820__)
  );
  LUT6 #(
    .INIT(64'hff00bf80aaaaaaaa)
  ) __2192__ (
    .I5(g109),
    .I4(__15__),
    .I3(__263__),
    .I2(g18),
    .I1(__212__),
    .I0(__171__),
    .O(__821__)
  );
  LUT4 #(
    .INIT(16'hbf80)
  ) __2193__ (
    .I3(__454__),
    .I2(__11__),
    .I1(g1696),
    .I0(__585__),
    .O(__822__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __2194__ (
    .I1(g1700),
    .I0(__284__),
    .O(__823__)
  );
  LUT4 #(
    .INIT(16'hbf80)
  ) __2195__ (
    .I3(__202__),
    .I2(__393__),
    .I1(__701__),
    .I0(__145__),
    .O(__824__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __2196__ (
    .I1(g109),
    .I0(__152__),
    .O(__825__)
  );
  LUT5 #(
    .INIT(32'h53ac0000)
  ) __2197__ (
    .I4(g109),
    .I3(__94__),
    .I2(g18),
    .I1(__204__),
    .I0(__44__),
    .O(__826__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __2198__ (
    .I1(g109),
    .I0(__386__),
    .O(__827__)
  );
  LUT6 #(
    .INIT(64'hff00bf80aaaaaaaa)
  ) __2199__ (
    .I5(g109),
    .I4(__276__),
    .I3(__65__),
    .I2(g18),
    .I1(__212__),
    .I0(__316__),
    .O(__828__)
  );
  LUT2 #(
    .INIT(4'h2)
  ) __2200__ (
    .I1(__11__),
    .I0(g1696),
    .O(__829__)
  );
  LUT6 #(
    .INIT(64'h00007fff00008000)
  ) __2201__ (
    .I5(__116__),
    .I4(__154__),
    .I3(__145__),
    .I2(__829__),
    .I1(__53__),
    .I0(__226__),
    .O(__830__)
  );
  LUT4 #(
    .INIT(16'h1fe0)
  ) __2202__ (
    .I3(__314__),
    .I2(__463__),
    .I1(__694__),
    .I0(__675__),
    .O(__831__)
  );
  LUT6 #(
    .INIT(64'hffff00f088888888)
  ) __2203__ (
    .I5(__508__),
    .I4(__700__),
    .I3(__699__),
    .I2(__831__),
    .I1(g109),
    .I0(__365__),
    .O(__832__)
  );
  LUT5 #(
    .INIT(32'h55595555)
  ) __2204__ (
    .I4(__468__),
    .I3(__297__),
    .I2(__156__),
    .I1(__61__),
    .I0(__91__),
    .O(__833__)
  );
  LUT6 #(
    .INIT(64'h8000bfffaaaaaaaa)
  ) __2205__ (
    .I5(__678__),
    .I4(__307__),
    .I3(__676__),
    .I2(__654__),
    .I1(__603__),
    .I0(__833__),
    .O(__834__)
  );
  LUT4 #(
    .INIT(16'ha3aa)
  ) __2206__ (
    .I3(g750),
    .I2(__438__),
    .I1(__834__),
    .I0(__475__),
    .O(__835__)
  );
  LUT4 #(
    .INIT(16'hbf80)
  ) __2207__ (
    .I3(__443__),
    .I2(__393__),
    .I1(__701__),
    .I0(__280__),
    .O(__836__)
  );
  LUT6 #(
    .INIT(64'hff00bf80aaaaaaaa)
  ) __2208__ (
    .I5(g109),
    .I4(__15__),
    .I3(__139__),
    .I2(g18),
    .I1(__212__),
    .I0(__356__),
    .O(__837__)
  );
  LUT6 #(
    .INIT(64'hff00bf80aaaaaaaa)
  ) __2209__ (
    .I5(g109),
    .I4(__15__),
    .I3(__62__),
    .I2(g18),
    .I1(__212__),
    .I0(__419__),
    .O(__838__)
  );
  LUT6 #(
    .INIT(64'hff00bf80aaaaaaaa)
  ) __2210__ (
    .I5(g109),
    .I4(__15__),
    .I3(__80__),
    .I2(g18),
    .I1(__212__),
    .I0(__107__),
    .O(__839__)
  );
  LUT6 #(
    .INIT(64'hff00bf80aaaaaaaa)
  ) __2211__ (
    .I5(g109),
    .I4(__15__),
    .I3(__78__),
    .I2(g18),
    .I1(__212__),
    .I0(__163__),
    .O(__840__)
  );
  LUT2 #(
    .INIT(4'he)
  ) __2212__ (
    .I1(g82),
    .I0(__30__),
    .O(__841__)
  );
  LUT4 #(
    .INIT(16'hf088)
  ) __2213__ (
    .I3(__508__),
    .I2(__232__),
    .I1(g109),
    .I0(__317__),
    .O(__842__)
  );
  LUT6 #(
    .INIT(64'hfffff0f0ffffccaa)
  ) __2214__ (
    .I5(__73__),
    .I4(__211__),
    .I3(g18),
    .I2(__565__),
    .I1(__44__),
    .I0(__282__),
    .O(__843__)
  );
  LUT4 #(
    .INIT(16'hccca)
  ) __2215__ (
    .I3(__11__),
    .I2(g1696),
    .I1(__204__),
    .I0(__843__),
    .O(__844__)
  );
  LUT6 #(
    .INIT(64'hf0f0e2e2f0f022e2)
  ) __2216__ (
    .I5(__37__),
    .I4(__345__),
    .I3(__685__),
    .I2(__391__),
    .I1(__734__),
    .I0(__291__),
    .O(__845__)
  );
  LUT4 #(
    .INIT(16'h0001)
  ) __2217__ (
    .I3(__422__),
    .I2(__265__),
    .I1(__373__),
    .I0(__242__),
    .O(__846__)
  );
  LUT6 #(
    .INIT(64'h00ff00fff0f01111)
  ) __2218__ (
    .I5(g18),
    .I4(__846__),
    .I3(__49__),
    .I2(__264__),
    .I1(__694__),
    .I0(__770__),
    .O(__847__)
  );
  LUT6 #(
    .INIT(64'h6996966900000000)
  ) __2219__ (
    .I5(g109),
    .I4(__128__),
    .I3(__483__),
    .I2(__163__),
    .I1(__203__),
    .I0(__847__),
    .O(__848__)
  );
  LUT6 #(
    .INIT(64'hff00bf80aaaaaaaa)
  ) __2220__ (
    .I5(g109),
    .I4(__276__),
    .I3(__312__),
    .I2(g18),
    .I1(__212__),
    .I0(__22__),
    .O(__849__)
  );
  LUT6 #(
    .INIT(64'hff00bf80aaaaaaaa)
  ) __2221__ (
    .I5(g109),
    .I4(__15__),
    .I3(__236__),
    .I2(g18),
    .I1(__212__),
    .I0(__135__),
    .O(__850__)
  );
  LUT4 #(
    .INIT(16'h88f0)
  ) __2222__ (
    .I3(__679__),
    .I2(__99__),
    .I1(g109),
    .I0(__88__),
    .O(__851__)
  );
  LUT5 #(
    .INIT(32'h53ac0000)
  ) __2223__ (
    .I4(g109),
    .I3(__34__),
    .I2(g18),
    .I1(__305__),
    .I0(__504__),
    .O(__852__)
  );
  LUT4 #(
    .INIT(16'h88f0)
  ) __2224__ (
    .I3(__679__),
    .I2(__267__),
    .I1(g109),
    .I0(__6__),
    .O(__853__)
  );
  LUT6 #(
    .INIT(64'hff00bf80aaaaaaaa)
  ) __2225__ (
    .I5(g109),
    .I4(__15__),
    .I3(__271__),
    .I2(g18),
    .I1(__212__),
    .I0(__382__),
    .O(__854__)
  );
  LUT6 #(
    .INIT(64'hff00bf80aaaaaaaa)
  ) __2226__ (
    .I5(g109),
    .I4(__15__),
    .I3(__178__),
    .I2(g18),
    .I1(__212__),
    .I0(__79__),
    .O(__855__)
  );
  LUT6 #(
    .INIT(64'hff00bf80aaaaaaaa)
  ) __2227__ (
    .I5(g109),
    .I4(__15__),
    .I3(__97__),
    .I2(g18),
    .I1(__212__),
    .I0(__69__),
    .O(__856__)
  );
  LUT5 #(
    .INIT(32'h6fffffff)
  ) __2228__ (
    .I4(g109),
    .I3(__278__),
    .I2(__196__),
    .I1(__500__),
    .I0(__200__),
    .O(__857__)
  );
  LUT4 #(
    .INIT(16'h88f0)
  ) __2229__ (
    .I3(__679__),
    .I2(__96__),
    .I1(g109),
    .I0(__346__),
    .O(__858__)
  );
  LUT4 #(
    .INIT(16'h0004)
  ) __2230__ (
    .I3(g41),
    .I2(g30),
    .I1(g48),
    .I0(g31),
    .O(__859__)
  );
  LUT4 #(
    .INIT(16'hbfff)
  ) __2231__ (
    .I3(__859__),
    .I2(__619__),
    .I1(__612__),
    .I0(__607__),
    .O(__860__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __2232__ (
    .I2(g18),
    .I1(__424__),
    .I0(__101__),
    .O(__861__)
  );
  LUT2 #(
    .INIT(4'he)
  ) __2233__ (
    .I1(g82),
    .I0(__41__),
    .O(__862__)
  );
  LUT4 #(
    .INIT(16'ha596)
  ) __2234__ (
    .I3(__37__),
    .I2(__32__),
    .I1(__12__),
    .I0(__60__),
    .O(__863__)
  );
  LUT6 #(
    .INIT(64'hfc0355aa00000000)
  ) __2235__ (
    .I5(__805__),
    .I4(__802__),
    .I3(__503__),
    .I2(__732__),
    .I1(__863__),
    .I0(__493__),
    .O(__864__)
  );
  LUT2 #(
    .INIT(4'he)
  ) __2236__ (
    .I1(__801__),
    .I0(__864__),
    .O(__865__)
  );
  LUT4 #(
    .INIT(16'h7800)
  ) __2237__ (
    .I3(__799__),
    .I2(__458__),
    .I1(__39__),
    .I0(__680__),
    .O(__866__)
  );
  LUT4 #(
    .INIT(16'h88f0)
  ) __2238__ (
    .I3(__679__),
    .I2(__10__),
    .I1(g109),
    .I0(__449__),
    .O(__867__)
  );
  LUT4 #(
    .INIT(16'hccca)
  ) __2239__ (
    .I3(__11__),
    .I2(g1696),
    .I1(__293__),
    .I0(__473__),
    .O(__868__)
  );
  LUT4 #(
    .INIT(16'hf088)
  ) __2240__ (
    .I3(__508__),
    .I2(__95__),
    .I1(g109),
    .I0(__85__),
    .O(__869__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __2241__ (
    .I2(__47__),
    .I1(__286__),
    .I0(__181__),
    .O(__870__)
  );
  LUT6 #(
    .INIT(64'h0000000000000001)
  ) __2242__ (
    .I5(__161__),
    .I4(__81__),
    .I3(__20__),
    .I2(__315__),
    .I1(__74__),
    .I0(__459__),
    .O(__871__)
  );
  LUT3 #(
    .INIT(8'h01)
  ) __2243__ (
    .I2(__243__),
    .I1(__83__),
    .I0(__152__),
    .O(__872__)
  );
  LUT6 #(
    .INIT(64'h0000000000000040)
  ) __2244__ (
    .I5(__354__),
    .I4(__386__),
    .I3(__63__),
    .I2(__872__),
    .I1(__871__),
    .I0(__308__),
    .O(__873__)
  );
  LUT2 #(
    .INIT(4'h2)
  ) __2245__ (
    .I1(__400__),
    .I0(__149__),
    .O(__874__)
  );
  LUT6 #(
    .INIT(64'hc03f3f6a3fc0c095)
  ) __2246__ (
    .I5(__150__),
    .I4(__92__),
    .I3(__487__),
    .I2(__767__),
    .I1(__874__),
    .I0(__873__),
    .O(__875__)
  );
  LUT5 #(
    .INIT(32'hf0f0f066)
  ) __2247__ (
    .I4(__11__),
    .I3(g1696),
    .I2(__82__),
    .I1(__875__),
    .I0(__847__),
    .O(__876__)
  );
  LUT4 #(
    .INIT(16'h88f0)
  ) __2248__ (
    .I3(__679__),
    .I2(__346__),
    .I1(g109),
    .I0(__91__),
    .O(__877__)
  );
  LUT6 #(
    .INIT(64'hffff555500330fff)
  ) __2249__ (
    .I5(__429__),
    .I4(__37__),
    .I3(__345__),
    .I2(__478__),
    .I1(__12__),
    .I0(__32__),
    .O(__878__)
  );
  LUT6 #(
    .INIT(64'hfffb00aa00000000)
  ) __2250__ (
    .I5(__368__),
    .I4(__37__),
    .I3(__345__),
    .I2(__12__),
    .I1(__478__),
    .I0(__32__),
    .O(__879__)
  );
  LUT3 #(
    .INIT(8'h04)
  ) __2251__ (
    .I2(__37__),
    .I1(__12__),
    .I0(__32__),
    .O(__880__)
  );
  LUT5 #(
    .INIT(32'h00007d55)
  ) __2252__ (
    .I4(__880__),
    .I3(__879__),
    .I2(__759__),
    .I1(__878__),
    .I0(__27__),
    .O(__881__)
  );
  LUT5 #(
    .INIT(32'h202a757f)
  ) __2253__ (
    .I4(__881__),
    .I3(__144__),
    .I2(__47__),
    .I1(__773__),
    .I0(__804__),
    .O(__882__)
  );
  LUT4 #(
    .INIT(16'hf088)
  ) __2254__ (
    .I3(__508__),
    .I2(__71__),
    .I1(g109),
    .I0(__406__),
    .O(__883__)
  );
  LUT5 #(
    .INIT(32'h55595555)
  ) __2255__ (
    .I4(__297__),
    .I3(__468__),
    .I2(__156__),
    .I1(__61__),
    .I0(__346__),
    .O(__884__)
  );
  LUT6 #(
    .INIT(64'haaccaaaaaa0faaaa)
  ) __2256__ (
    .I5(__679__),
    .I4(g750),
    .I3(__438__),
    .I2(__884__),
    .I1(__496__),
    .I0(__388__),
    .O(__885__)
  );
  LUT4 #(
    .INIT(16'hf088)
  ) __2257__ (
    .I3(__508__),
    .I2(__317__),
    .I1(g109),
    .I0(__377__),
    .O(__886__)
  );
  LUT6 #(
    .INIT(64'hcdccfeccfdcccecc)
  ) __2258__ (
    .I5(__717__),
    .I4(__176__),
    .I3(__725__),
    .I2(__723__),
    .I1(__719__),
    .I0(__173__),
    .O(__887__)
  );
  LUT5 #(
    .INIT(32'h55555559)
  ) __2259__ (
    .I4(__297__),
    .I3(__468__),
    .I2(__156__),
    .I1(__61__),
    .I0(__96__),
    .O(__888__)
  );
  LUT6 #(
    .INIT(64'h8000bfffaaaaaaaa)
  ) __2260__ (
    .I5(__678__),
    .I4(__498__),
    .I3(__676__),
    .I2(__654__),
    .I1(__603__),
    .I0(__888__),
    .O(__889__)
  );
  LUT4 #(
    .INIT(16'ha3aa)
  ) __2261__ (
    .I3(g750),
    .I2(__438__),
    .I1(__889__),
    .I0(__474__),
    .O(__890__)
  );
  LUT6 #(
    .INIT(64'hff00bf80aaaaaaaa)
  ) __2262__ (
    .I5(g109),
    .I4(__15__),
    .I3(__321__),
    .I2(g18),
    .I1(__212__),
    .I0(__390__),
    .O(__891__)
  );
  LUT5 #(
    .INIT(32'hccccfcfd)
  ) __2263__ (
    .I4(__37__),
    .I3(__32__),
    .I2(__345__),
    .I1(__357__),
    .I0(__12__),
    .O(__892__)
  );
  LUT5 #(
    .INIT(32'haaaa0a08)
  ) __2264__ (
    .I4(__37__),
    .I3(__32__),
    .I2(__345__),
    .I1(__12__),
    .I0(__130__),
    .O(__893__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __2265__ (
    .I3(__11__),
    .I2(g1696),
    .I1(__35__),
    .I0(__275__),
    .O(__894__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __2266__ (
    .I2(g109),
    .I1(g743),
    .I0(g744),
    .O(__895__)
  );
  LUT4 #(
    .INIT(16'h88f0)
  ) __2267__ (
    .I3(__679__),
    .I2(__341__),
    .I1(g109),
    .I0(__55__),
    .O(__896__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __2268__ (
    .I1(g109),
    .I0(__302__),
    .O(__897__)
  );
  LUT5 #(
    .INIT(32'h53ac0000)
  ) __2269__ (
    .I4(g109),
    .I3(__244__),
    .I2(g18),
    .I1(__451__),
    .I0(__24__),
    .O(__898__)
  );
  LUT6 #(
    .INIT(64'h000000007f800000)
  ) __2270__ (
    .I5(__407__),
    .I4(g109),
    .I3(__42__),
    .I2(__378__),
    .I1(__497__),
    .I0(__683__),
    .O(__899__)
  );
  LUT4 #(
    .INIT(16'hccca)
  ) __2271__ (
    .I3(__11__),
    .I2(g1696),
    .I1(__219__),
    .I0(__332__),
    .O(__900__)
  );
  LUT6 #(
    .INIT(64'hfefe7f7ffe7f7ffe)
  ) __2272__ (
    .I5(__37__),
    .I4(__32__),
    .I3(__12__),
    .I2(__60__),
    .I1(__110__),
    .I0(__503__),
    .O(__901__)
  );
  LUT6 #(
    .INIT(64'hfc0355aa00000000)
  ) __2273__ (
    .I5(__805__),
    .I4(__802__),
    .I3(__479__),
    .I2(__732__),
    .I1(__901__),
    .I0(__241__),
    .O(__902__)
  );
  LUT2 #(
    .INIT(4'he)
  ) __2274__ (
    .I1(__801__),
    .I0(__902__),
    .O(__903__)
  );
  LUT6 #(
    .INIT(64'h55555555c0003fff)
  ) __2275__ (
    .I5(g18),
    .I4(__20__),
    .I3(__400__),
    .I2(__516__),
    .I1(__149__),
    .I0(__174__),
    .O(__904__)
  );
  LUT4 #(
    .INIT(16'haaa3)
  ) __2276__ (
    .I3(__11__),
    .I2(g1696),
    .I1(__904__),
    .I0(__164__),
    .O(__905__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __2277__ (
    .I1(g109),
    .I0(__480__),
    .O(__906__)
  );
  LUT6 #(
    .INIT(64'hff00bf80aaaaaaaa)
  ) __2278__ (
    .I5(g109),
    .I4(__15__),
    .I3(__375__),
    .I2(g18),
    .I1(__212__),
    .I0(__376__),
    .O(__907__)
  );
  LUT5 #(
    .INIT(32'haaaa0a08)
  ) __2279__ (
    .I4(__273__),
    .I3(__414__),
    .I2(__295__),
    .I1(__112__),
    .I0(__364__),
    .O(__908__)
  );
  LUT2 #(
    .INIT(4'hd)
  ) __2280__ (
    .I1(__383__),
    .I0(g1700),
    .O(__909__)
  );
  LUT4 #(
    .INIT(16'hf088)
  ) __2281__ (
    .I3(__508__),
    .I2(__255__),
    .I1(g109),
    .I0(__326__),
    .O(__910__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __2282__ (
    .I1(g109),
    .I0(__44__),
    .O(__911__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __2283__ (
    .I1(g109),
    .I0(__664__),
    .O(__912__)
  );
  LUT6 #(
    .INIT(64'hfffff0f0ffffccaa)
  ) __2284__ (
    .I5(__73__),
    .I4(__211__),
    .I3(g18),
    .I2(__912__),
    .I1(__392__),
    .I0(__448__),
    .O(__913__)
  );
  LUT4 #(
    .INIT(16'hccca)
  ) __2285__ (
    .I3(__11__),
    .I2(g1696),
    .I1(__142__),
    .I0(__913__),
    .O(__914__)
  );
  LUT4 #(
    .INIT(16'h88f0)
  ) __2286__ (
    .I3(__679__),
    .I2(__423__),
    .I1(g109),
    .I0(__102__),
    .O(__915__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __2287__ (
    .I1(g109),
    .I0(__459__),
    .O(__916__)
  );
  LUT3 #(
    .INIT(8'hbf)
  ) __2288__ (
    .I2(__619__),
    .I1(__612__),
    .I0(__607__),
    .O(__917__)
  );
  LUT6 #(
    .INIT(64'h0000000000000040)
  ) __2289__ (
    .I5(__694__),
    .I4(__585__),
    .I3(__745__),
    .I2(__602__),
    .I1(__759__),
    .I0(__773__),
    .O(__918__)
  );
  LUT4 #(
    .INIT(16'ha3aa)
  ) __2290__ (
    .I3(g1696),
    .I2(__11__),
    .I1(__918__),
    .I0(__264__),
    .O(__919__)
  );
  LUT4 #(
    .INIT(16'hbf80)
  ) __2291__ (
    .I3(__397__),
    .I2(__393__),
    .I1(__701__),
    .I0(__324__),
    .O(__920__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __2292__ (
    .I1(g109),
    .I0(__79__),
    .O(__921__)
  );
  LUT6 #(
    .INIT(64'hff00bf80aaaaaaaa)
  ) __2293__ (
    .I5(g109),
    .I4(__276__),
    .I3(__342__),
    .I2(g18),
    .I1(__212__),
    .I0(__31__),
    .O(__922__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __2294__ (
    .I1(g109),
    .I0(__415__),
    .O(__923__)
  );
  LUT5 #(
    .INIT(32'h53ac0000)
  ) __2295__ (
    .I4(g109),
    .I3(__372__),
    .I2(g18),
    .I1(__403__),
    .I0(__224__),
    .O(__924__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __2296__ (
    .I2(g18),
    .I1(__225__),
    .I0(__492__),
    .O(__925__)
  );
  LUT3 #(
    .INIT(8'h40)
  ) __2297__ (
    .I2(g109),
    .I1(__400__),
    .I0(__183__),
    .O(__926__)
  );
  LUT6 #(
    .INIT(64'h0001ffffffff0001)
  ) __2298__ (
    .I5(__716__),
    .I4(__269__),
    .I3(__295__),
    .I2(__414__),
    .I1(__112__),
    .I0(__273__),
    .O(__927__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __2299__ (
    .I2(g18),
    .I1(__224__),
    .I0(__403__),
    .O(__928__)
  );
  LUT6 #(
    .INIT(64'hf0f0e2e2f0f022e2)
  ) __2300__ (
    .I5(__37__),
    .I4(__345__),
    .I3(__685__),
    .I2(__491__),
    .I1(__734__),
    .I0(__446__),
    .O(__929__)
  );
  LUT6 #(
    .INIT(64'hff00bf80aaaaaaaa)
  ) __2301__ (
    .I5(g109),
    .I4(__276__),
    .I3(__442__),
    .I2(g18),
    .I1(__212__),
    .I0(__13__),
    .O(__930__)
  );
  LUT5 #(
    .INIT(32'h0c0c060c)
  ) __2302__ (
    .I4(__11__),
    .I3(g1696),
    .I2(__154__),
    .I1(__53__),
    .I0(__226__),
    .O(__931__)
  );
  LUT4 #(
    .INIT(16'h88f0)
  ) __2303__ (
    .I3(__679__),
    .I2(__165__),
    .I1(g109),
    .I0(__272__),
    .O(__932__)
  );
  LUT2 #(
    .INIT(4'he)
  ) __2304__ (
    .I1(g82),
    .I0(__184__),
    .O(__933__)
  );
  LUT4 #(
    .INIT(16'hccca)
  ) __2305__ (
    .I3(__11__),
    .I2(g1696),
    .I1(__186__),
    .I0(__35__),
    .O(__934__)
  );
  LUT5 #(
    .INIT(32'h80000000)
  ) __2306__ (
    .I4(__405__),
    .I3(__456__),
    .I2(__237__),
    .I1(__453__),
    .I0(__214__),
    .O(__935__)
  );
  LUT4 #(
    .INIT(16'h0060)
  ) __2307__ (
    .I3(__407__),
    .I2(g109),
    .I1(__445__),
    .I0(__935__),
    .O(__936__)
  );
  LUT6 #(
    .INIT(64'hff00f870ff00ff00)
  ) __2308__ (
    .I5(__680__),
    .I4(__519__),
    .I3(__401__),
    .I2(__21__),
    .I1(g109),
    .I0(__380__),
    .O(__937__)
  );
  LUT3 #(
    .INIT(8'hfe)
  ) __2309__ (
    .I2(g41),
    .I1(g30),
    .I0(g31),
    .O(__938__)
  );
  LUT6 #(
    .INIT(64'hefffffffffffffff)
  ) __2310__ (
    .I5(g48),
    .I4(__584__),
    .I3(__579__),
    .I2(__571__),
    .I1(__938__),
    .I0(__547__),
    .O(__939__)
  );
  LUT6 #(
    .INIT(64'h3f00f3c500000000)
  ) __2311__ (
    .I5(g18),
    .I4(__37__),
    .I3(__12__),
    .I2(__32__),
    .I1(__733__),
    .I0(__345__),
    .O(__940__)
  );
  LUT4 #(
    .INIT(16'hf088)
  ) __2312__ (
    .I3(__508__),
    .I2(__396__),
    .I1(g109),
    .I0(__232__),
    .O(__941__)
  );
  LUT6 #(
    .INIT(64'h555555550300fcff)
  ) __2313__ (
    .I5(g18),
    .I4(__63__),
    .I3(__516__),
    .I2(__400__),
    .I1(__149__),
    .I0(__494__),
    .O(__942__)
  );
  LUT4 #(
    .INIT(16'haaa3)
  ) __2314__ (
    .I3(__11__),
    .I2(g1696),
    .I1(__942__),
    .I0(__16__),
    .O(__943__)
  );
  LUT6 #(
    .INIT(64'hf0f0e2e2f0f022e2)
  ) __2315__ (
    .I5(__37__),
    .I4(__345__),
    .I3(__685__),
    .I2(__446__),
    .I1(__734__),
    .I0(__391__),
    .O(__944__)
  );
  LUT6 #(
    .INIT(64'hff00bf80aaaaaaaa)
  ) __2316__ (
    .I5(g109),
    .I4(__15__),
    .I3(__131__),
    .I2(g18),
    .I1(__212__),
    .I0(__143__),
    .O(__945__)
  );
  LUT4 #(
    .INIT(16'h88f0)
  ) __2317__ (
    .I3(__679__),
    .I2(__188__),
    .I1(g109),
    .I0(__99__),
    .O(__946__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __2318__ (
    .I1(g109),
    .I0(__504__),
    .O(__947__)
  );
  LUT5 #(
    .INIT(32'hffff5501)
  ) __2319__ (
    .I4(__118__),
    .I3(__295__),
    .I2(__414__),
    .I1(__112__),
    .I0(__273__),
    .O(__948__)
  );
  LUT5 #(
    .INIT(32'haaaa0a08)
  ) __2320__ (
    .I4(__273__),
    .I3(__414__),
    .I2(__295__),
    .I1(__112__),
    .I0(__151__),
    .O(__949__)
  );
  LUT3 #(
    .INIT(8'hb0)
  ) __2321__ (
    .I2(__242__),
    .I1(g1696),
    .I0(__11__),
    .O(__950__)
  );
  LUT4 #(
    .INIT(16'h88f0)
  ) __2322__ (
    .I3(__679__),
    .I2(__91__),
    .I1(g109),
    .I0(__10__),
    .O(__951__)
  );
  LUT4 #(
    .INIT(16'h880f)
  ) __2323__ (
    .I3(__679__),
    .I2(__529__),
    .I1(g109),
    .I0(__188__),
    .O(__952__)
  );
  LUT4 #(
    .INIT(16'hf800)
  ) __2324__ (
    .I3(g109),
    .I2(__276__),
    .I1(g18),
    .I0(__212__),
    .O(__953__)
  );
  LUT5 #(
    .INIT(32'hbfff0000)
  ) __2325__ (
    .I4(g109),
    .I3(__636__),
    .I2(__627__),
    .I1(__622__),
    .I0(__547__),
    .O(__954__)
  );
  LUT4 #(
    .INIT(16'hbf80)
  ) __2326__ (
    .I3(__199__),
    .I2(__11__),
    .I1(g1696),
    .I0(__954__),
    .O(__955__)
  );
  LUT6 #(
    .INIT(64'he4e464e400000000)
  ) __2327__ (
    .I5(g18),
    .I4(__56__),
    .I3(__295__),
    .I2(__414__),
    .I1(__273__),
    .I0(__718__),
    .O(__956__)
  );
  LUT4 #(
    .INIT(16'hbf80)
  ) __2328__ (
    .I3(__147__),
    .I2(__38__),
    .I1(__150__),
    .I0(__226__),
    .O(__957__)
  );
  LUT5 #(
    .INIT(32'h53ac0000)
  ) __2329__ (
    .I4(g109),
    .I3(__466__),
    .I2(g18),
    .I1(__117__),
    .I0(__24__),
    .O(__958__)
  );
  LUT4 #(
    .INIT(16'haaa3)
  ) __2330__ (
    .I3(__11__),
    .I2(g1696),
    .I1(__517__),
    .I0(__374__),
    .O(__959__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __2331__ (
    .I1(g109),
    .I0(__74__),
    .O(__960__)
  );
  LUT6 #(
    .INIT(64'h0000ffff8fffffff)
  ) __2332__ (
    .I5(__56__),
    .I4(__512__),
    .I3(__295__),
    .I2(__273__),
    .I1(__718__),
    .I0(__471__),
    .O(__961__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __2333__ (
    .I2(g18),
    .I1(__295__),
    .I0(__961__),
    .O(__962__)
  );
  LUT6 #(
    .INIT(64'hffff0f0fffff3355)
  ) __2334__ (
    .I5(__73__),
    .I4(__211__),
    .I3(g18),
    .I2(__585__),
    .I1(__24__),
    .I0(__451__),
    .O(__963__)
  );
  LUT4 #(
    .INIT(16'haaa3)
  ) __2335__ (
    .I3(__11__),
    .I2(g1696),
    .I1(__963__),
    .I0(__117__),
    .O(__964__)
  );
  LUT6 #(
    .INIT(64'hffff7fffffffffff)
  ) __2336__ (
    .I5(__859__),
    .I4(__547__),
    .I3(__601__),
    .I2(__595__),
    .I1(__590__),
    .I0(__588__),
    .O(__965__)
  );
  LUT4 #(
    .INIT(16'h88f0)
  ) __2337__ (
    .I3(__679__),
    .I2(__88__),
    .I1(g109),
    .I0(__208__),
    .O(__966__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __2338__ (
    .I1(g109),
    .I0(__113__),
    .O(__967__)
  );
  LUT6 #(
    .INIT(64'h0000000080000000)
  ) __2339__ (
    .I5(__11__),
    .I4(g1696),
    .I3(__116__),
    .I2(__145__),
    .I1(__53__),
    .I0(__226__),
    .O(__968__)
  );
  LUT3 #(
    .INIT(8'h06)
  ) __2340__ (
    .I2(__154__),
    .I1(__324__),
    .I0(__968__),
    .O(__969__)
  );
  LUT3 #(
    .INIT(8'h60)
  ) __2341__ (
    .I2(__196__),
    .I1(g750),
    .I0(__438__),
    .O(__970__)
  );
  LUT6 #(
    .INIT(64'hff00f870ff00ff00)
  ) __2342__ (
    .I5(__680__),
    .I4(__519__),
    .I3(__18__),
    .I2(__301__),
    .I1(g109),
    .I0(__380__),
    .O(__971__)
  );
  LUT6 #(
    .INIT(64'h00aa00ccf0f0f0f0)
  ) __2343__ (
    .I5(__802__),
    .I4(__479__),
    .I3(__732__),
    .I2(__281__),
    .I1(__728__),
    .I0(__730__),
    .O(__972__)
  );
  LUT4 #(
    .INIT(16'hbeaa)
  ) __2344__ (
    .I3(__805__),
    .I2(__327__),
    .I1(__972__),
    .I0(__801__),
    .O(__973__)
  );
  LUT6 #(
    .INIT(64'hf0f0e2e2f0f022e2)
  ) __2345__ (
    .I5(__37__),
    .I4(__345__),
    .I3(__685__),
    .I2(__281__),
    .I1(__734__),
    .I0(__241__),
    .O(__974__)
  );
  LUT6 #(
    .INIT(64'hff00bf80aaaaaaaa)
  ) __2346__ (
    .I5(g109),
    .I4(__15__),
    .I3(__159__),
    .I2(g18),
    .I1(__212__),
    .I0(__203__),
    .O(__975__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __2347__ (
    .I1(g109),
    .I0(__155__),
    .O(__976__)
  );
  LUT6 #(
    .INIT(64'hff00bf80aaaaaaaa)
  ) __2348__ (
    .I5(g109),
    .I4(__15__),
    .I3(__191__),
    .I2(g18),
    .I1(__212__),
    .I0(__277__),
    .O(__977__)
  );
  LUT3 #(
    .INIT(8'hb0)
  ) __2349__ (
    .I2(__373__),
    .I1(g1696),
    .I0(__11__),
    .O(__978__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __2350__ (
    .I2(g109),
    .I1(__69__),
    .I0(__904__),
    .O(__979__)
  );
  LUT6 #(
    .INIT(64'hf0f0e2e2f0f022e2)
  ) __2351__ (
    .I5(__37__),
    .I4(__345__),
    .I3(__685__),
    .I2(__291__),
    .I1(__734__),
    .I0(__281__),
    .O(__980__)
  );
  LUT5 #(
    .INIT(32'h55595555)
  ) __2352__ (
    .I4(__297__),
    .I3(__61__),
    .I2(__156__),
    .I1(__468__),
    .I0(__157__),
    .O(__981__)
  );
  LUT6 #(
    .INIT(64'h8000bfffaaaaaaaa)
  ) __2353__ (
    .I5(__678__),
    .I4(__231__),
    .I3(__676__),
    .I2(__654__),
    .I1(__603__),
    .I0(__981__),
    .O(__982__)
  );
  LUT4 #(
    .INIT(16'ha3aa)
  ) __2354__ (
    .I3(g750),
    .I2(__438__),
    .I1(__982__),
    .I0(__275__),
    .O(__983__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __2355__ (
    .I1(g109),
    .I0(__315__),
    .O(__984__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __2356__ (
    .I1(__196__),
    .I0(g750),
    .O(__985__)
  );
  LUT6 #(
    .INIT(64'h0caa0c0c0c0c0c0c)
  ) __2357__ (
    .I5(__56__),
    .I4(__512__),
    .I3(__295__),
    .I2(__511__),
    .I1(__464__),
    .I0(__173__),
    .O(__986__)
  );
  LUT3 #(
    .INIT(8'h60)
  ) __2358__ (
    .I2(__799__),
    .I1(__39__),
    .I0(__680__),
    .O(__987__)
  );
  LUT4 #(
    .INIT(16'h8000)
  ) __2359__ (
    .I3(__182__),
    .I2(__439__),
    .I1(__500__),
    .I0(__200__),
    .O(__988__)
  );
  LUT6 #(
    .INIT(64'h7800000000000000)
  ) __2360__ (
    .I5(g109),
    .I4(__278__),
    .I3(__196__),
    .I2(__266__),
    .I1(__421__),
    .I0(__988__),
    .O(__989__)
  );
  LUT4 #(
    .INIT(16'hbf80)
  ) __2361__ (
    .I3(__304__),
    .I2(__38__),
    .I1(__150__),
    .I0(__324__),
    .O(__990__)
  );
  LUT4 #(
    .INIT(16'hccca)
  ) __2362__ (
    .I3(__11__),
    .I2(g1696),
    .I1(__154__),
    .I0(__385__),
    .O(__991__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __2363__ (
    .I1(g109),
    .I0(__243__),
    .O(__992__)
  );
  LUT5 #(
    .INIT(32'h53ac0000)
  ) __2364__ (
    .I4(g109),
    .I3(__135__),
    .I2(g18),
    .I1(__215__),
    .I0(__504__),
    .O(__993__)
  );
  LUT5 #(
    .INIT(32'h53ac0000)
  ) __2365__ (
    .I4(g109),
    .I3(__143__),
    .I2(g18),
    .I1(__282__),
    .I0(__44__),
    .O(__994__)
  );
  LUT4 #(
    .INIT(16'hbf80)
  ) __2366__ (
    .I3(__109__),
    .I2(__393__),
    .I1(__701__),
    .I0(__25__),
    .O(__995__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __2367__ (
    .I1(g109),
    .I0(__114__),
    .O(__996__)
  );
  LUT6 #(
    .INIT(64'hf8ff0f0000000000)
  ) __2368__ (
    .I5(__996__),
    .I4(__104__),
    .I3(__436__),
    .I2(__679__),
    .I1(__121__),
    .I0(__115__),
    .O(__997__)
  );
  LUT5 #(
    .INIT(32'h00545500)
  ) __2369__ (
    .I4(__357__),
    .I3(__166__),
    .I2(__437__),
    .I1(__216__),
    .I0(__804__),
    .O(__998__)
  );
  LUT3 #(
    .INIT(8'hb0)
  ) __2370__ (
    .I2(__150__),
    .I1(g1696),
    .I0(__11__),
    .O(__999__)
  );
  LUT5 #(
    .INIT(32'h53ac0000)
  ) __2371__ (
    .I4(g109),
    .I3(__316__),
    .I2(g18),
    .I1(__492__),
    .I0(__225__),
    .O(__1000__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __2372__ (
    .I1(g109),
    .I0(__81__),
    .O(__1001__)
  );
  LUT6 #(
    .INIT(64'hfbfa000000000000)
  ) __2373__ (
    .I5(g109),
    .I4(__268__),
    .I3(__489__),
    .I2(g881),
    .I1(__198__),
    .I0(__245__),
    .O(__1002__)
  );
  LUT3 #(
    .INIT(8'h35)
  ) __2374__ (
    .I2(g18),
    .I1(__185__),
    .I0(__16__),
    .O(__1003__)
  );
  LUT6 #(
    .INIT(64'h0f030003aaaaaaaa)
  ) __2375__ (
    .I5(__747__),
    .I4(__602__),
    .I3(__73__),
    .I2(__211__),
    .I1(__1003__),
    .I0(__218__),
    .O(__1004__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __2376__ (
    .I3(__11__),
    .I2(g1696),
    .I1(__40__),
    .I0(__388__),
    .O(__1005__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __2377__ (
    .I1(g109),
    .I0(__288__),
    .O(__1006__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __2378__ (
    .I3(__11__),
    .I2(g1696),
    .I1(__412__),
    .I0(__54__),
    .O(__1007__)
  );
  LUT3 #(
    .INIT(8'h40)
  ) __2379__ (
    .I2(g18),
    .I1(__212__),
    .I0(__15__),
    .O(__1008__)
  );
  LUT6 #(
    .INIT(64'h0000000080000000)
  ) __2380__ (
    .I5(__203__),
    .I4(__356__),
    .I3(__1008__),
    .I2(__128__),
    .I1(__483__),
    .I0(__69__),
    .O(__1009__)
  );
  LUT5 #(
    .INIT(32'h00000040)
  ) __2381__ (
    .I4(__259__),
    .I3(__217__),
    .I2(__277__),
    .I1(__163__),
    .I0(__148__),
    .O(__1010__)
  );
  LUT6 #(
    .INIT(64'h8000000000000000)
  ) __2382__ (
    .I5(__382__),
    .I4(__210__),
    .I3(__419__),
    .I2(__240__),
    .I1(__1010__),
    .I0(__1009__),
    .O(__1011__)
  );
  LUT3 #(
    .INIT(8'he0)
  ) __2383__ (
    .I2(g109),
    .I1(__502__),
    .I0(__1011__),
    .O(__1012__)
  );
  LUT6 #(
    .INIT(64'h000000008aaa0000)
  ) __2384__ (
    .I5(__170__),
    .I4(g109),
    .I3(__619__),
    .I2(__612__),
    .I1(__607__),
    .I0(__106__),
    .O(__1013__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __2385__ (
    .I2(g109),
    .I1(__664__),
    .I0(__52__),
    .O(__1014__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __2386__ (
    .I2(g109),
    .I1(__320__),
    .I0(__772__),
    .O(__1015__)
  );
  LUT6 #(
    .INIT(64'h00000000bfff0000)
  ) __2387__ (
    .I5(__146__),
    .I4(g109),
    .I3(__649__),
    .I2(__647__),
    .I1(__642__),
    .I0(__639__),
    .O(__1016__)
  );
  LUT4 #(
    .INIT(16'h8000)
  ) __2388__ (
    .I3(g109),
    .I2(__675__),
    .I1(__38__),
    .I0(__150__),
    .O(__1017__)
  );
  LUT6 #(
    .INIT(64'hfffffffe00000001)
  ) __2389__ (
    .I5(__776__),
    .I4(__1017__),
    .I3(__1016__),
    .I2(__1015__),
    .I1(__1014__),
    .I0(__1013__),
    .O(__1018__)
  );
  LUT5 #(
    .INIT(32'h53ac0000)
  ) __2390__ (
    .I4(g109),
    .I3(__227__),
    .I2(g18),
    .I1(__58__),
    .I0(__185__),
    .O(__1019__)
  );
  LUT5 #(
    .INIT(32'h55555559)
  ) __2391__ (
    .I4(__297__),
    .I3(__468__),
    .I2(__61__),
    .I1(__156__),
    .I0(__449__),
    .O(__1020__)
  );
  LUT6 #(
    .INIT(64'h8000bfffaaaaaaaa)
  ) __2392__ (
    .I5(__678__),
    .I4(__290__),
    .I3(__676__),
    .I2(__654__),
    .I1(__603__),
    .I0(__1020__),
    .O(__1021__)
  );
  LUT4 #(
    .INIT(16'ha3aa)
  ) __2393__ (
    .I3(g750),
    .I2(__438__),
    .I1(__1021__),
    .I0(__311__),
    .O(__1022__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __2394__ (
    .I2(g109),
    .I1(g741),
    .I0(g742),
    .O(__1023__)
  );
  LUT4 #(
    .INIT(16'hbf80)
  ) __2395__ (
    .I3(__177__),
    .I2(__38__),
    .I1(__150__),
    .I0(__53__),
    .O(__1024__)
  );
  LUT4 #(
    .INIT(16'h88f0)
  ) __2396__ (
    .I3(__679__),
    .I2(__410__),
    .I1(g109),
    .I0(__347__),
    .O(__1025__)
  );
  LUT4 #(
    .INIT(16'hac00)
  ) __2397__ (
    .I3(g18),
    .I2(__733__),
    .I1(__32__),
    .I0(__12__),
    .O(__1026__)
  );
  LUT5 #(
    .INIT(32'h00000010)
  ) __2398__ (
    .I4(__56__),
    .I3(__295__),
    .I2(__273__),
    .I1(__414__),
    .I0(__112__),
    .O(__1027__)
  );
  LUT6 #(
    .INIT(64'hfdffcc0000000000)
  ) __2399__ (
    .I5(g18),
    .I4(__56__),
    .I3(__512__),
    .I2(__295__),
    .I1(__1027__),
    .I0(__258__),
    .O(__1028__)
  );
  LUT6 #(
    .INIT(64'h7800000000000000)
  ) __2400__ (
    .I5(g109),
    .I4(__278__),
    .I3(__196__),
    .I2(__439__),
    .I1(__500__),
    .I0(__200__),
    .O(__1029__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __2401__ (
    .I2(g109),
    .I1(__38__),
    .I0(__150__),
    .O(__1030__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __2402__ (
    .I2(g18),
    .I1(__504__),
    .I0(__305__),
    .O(__1031__)
  );
  LUT2 #(
    .INIT(4'he)
  ) __2403__ (
    .I1(g82),
    .I0(__3__),
    .O(__1032__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __2404__ (
    .I2(g18),
    .I1(__494__),
    .I0(__348__),
    .O(__1033__)
  );
  LUT6 #(
    .INIT(64'hff00bf80aaaaaaaa)
  ) __2405__ (
    .I5(g109),
    .I4(__276__),
    .I3(__172__),
    .I2(g18),
    .I1(__212__),
    .I0(__227__),
    .O(__1034__)
  );
  LUT3 #(
    .INIT(8'h04)
  ) __2406__ (
    .I2(__407__),
    .I1(g109),
    .I0(__214__),
    .O(__1035__)
  );
  LUT5 #(
    .INIT(32'h55595555)
  ) __2407__ (
    .I4(__297__),
    .I3(__468__),
    .I2(__61__),
    .I1(__156__),
    .I0(__267__),
    .O(__1036__)
  );
  LUT6 #(
    .INIT(64'haaccaaaaaa0faaaa)
  ) __2408__ (
    .I5(__679__),
    .I4(g750),
    .I3(__438__),
    .I2(__1036__),
    .I1(__123__),
    .I0(__86__),
    .O(__1037__)
  );
  LUT3 #(
    .INIT(8'h40)
  ) __2409__ (
    .I2(g18),
    .I1(__212__),
    .I0(__276__),
    .O(__1038__)
  );
  LUT6 #(
    .INIT(64'h0000000000000040)
  ) __2410__ (
    .I5(__372__),
    .I4(__70__),
    .I3(__22__),
    .I2(__31__),
    .I1(__1038__),
    .I0(__34__),
    .O(__1039__)
  );
  LUT5 #(
    .INIT(32'h00008000)
  ) __2411__ (
    .I4(__387__),
    .I3(__105__),
    .I2(__94__),
    .I1(__13__),
    .I0(__227__),
    .O(__1040__)
  );
  LUT6 #(
    .INIT(64'h0000000000000040)
  ) __2412__ (
    .I5(__220__),
    .I4(__476__),
    .I3(__466__),
    .I2(__1040__),
    .I1(__1039__),
    .I0(__316__),
    .O(__1041__)
  );
  LUT3 #(
    .INIT(8'he0)
  ) __2413__ (
    .I2(g109),
    .I1(__495__),
    .I0(__1041__),
    .O(__1042__)
  );
  LUT6 #(
    .INIT(64'hff00bf80aaaaaaaa)
  ) __2414__ (
    .I5(g109),
    .I4(__276__),
    .I3(__310__),
    .I2(g18),
    .I1(__212__),
    .I0(__105__),
    .O(__1043__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __2415__ (
    .I2(g109),
    .I1(__259__),
    .I0(__942__),
    .O(__1044__)
  );
  LUT6 #(
    .INIT(64'h55505553aaaaaaab)
  ) __2416__ (
    .I5(__512__),
    .I4(__295__),
    .I3(__414__),
    .I2(__112__),
    .I1(__273__),
    .I0(__292__),
    .O(__1045__)
  );
  LUT5 #(
    .INIT(32'h69960000)
  ) __2417__ (
    .I4(g109),
    .I3(__372__),
    .I2(__70__),
    .I1(__22__),
    .I0(__13__),
    .O(__1046__)
  );
  LUT4 #(
    .INIT(16'hf088)
  ) __2418__ (
    .I3(__508__),
    .I2(__85__),
    .I1(g109),
    .I0(__68__),
    .O(__1047__)
  );
  LUT3 #(
    .INIT(8'h35)
  ) __2419__ (
    .I2(g18),
    .I1(__224__),
    .I0(__82__),
    .O(__1048__)
  );
  LUT6 #(
    .INIT(64'h0f030003aaaaaaaa)
  ) __2420__ (
    .I5(__747__),
    .I4(__954__),
    .I3(__73__),
    .I2(__211__),
    .I1(__1048__),
    .I0(__403__),
    .O(__1049__)
  );
  LUT5 #(
    .INIT(32'hee00f0f0)
  ) __2421__ (
    .I4(__723__),
    .I3(__717__),
    .I2(__258__),
    .I1(__714__),
    .I0(__712__),
    .O(__1050__)
  );
  LUT4 #(
    .INIT(16'hbeaa)
  ) __2422__ (
    .I3(__725__),
    .I2(__17__),
    .I1(__1050__),
    .I0(__719__),
    .O(__1051__)
  );
  LUT3 #(
    .INIT(8'h40)
  ) __2423__ (
    .I2(g109),
    .I1(__489__),
    .I0(__198__),
    .O(__1052__)
  );
  LUT4 #(
    .INIT(16'hbf00)
  ) __2424__ (
    .I3(g109),
    .I2(__619__),
    .I1(__612__),
    .I0(__607__),
    .O(__1053__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __2425__ (
    .I2(g109),
    .I1(__380__),
    .I0(__772__),
    .O(__1054__)
  );
  LUT5 #(
    .INIT(32'h0777ffff)
  ) __2426__ (
    .I4(g109),
    .I3(__745__),
    .I2(g881),
    .I1(__773__),
    .I0(g877),
    .O(__1055__)
  );
  LUT6 #(
    .INIT(64'h0000153f00000000)
  ) __2427__ (
    .I5(__1055__),
    .I4(__1054__),
    .I3(__585__),
    .I2(__519__),
    .I1(__1053__),
    .I0(__1052__),
    .O(__1056__)
  );
  LUT4 #(
    .INIT(16'h88f0)
  ) __2428__ (
    .I3(__679__),
    .I2(__449__),
    .I1(g109),
    .I0(__267__),
    .O(__1057__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __2429__ (
    .I3(__11__),
    .I2(g1696),
    .I1(__134__),
    .I0(__330__),
    .O(__1058__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __2430__ (
    .I1(__479__),
    .I0(__730__),
    .O(__1059__)
  );
  LUT3 #(
    .INIT(8'he1)
  ) __2431__ (
    .I2(__32__),
    .I1(__37__),
    .I0(__12__),
    .O(__1060__)
  );
  LUT5 #(
    .INIT(32'h00000004)
  ) __2432__ (
    .I4(__60__),
    .I3(__110__),
    .I2(__503__),
    .I1(__1060__),
    .I0(__479__),
    .O(__1061__)
  );
  LUT6 #(
    .INIT(64'h00aa00ccf0f0f0f0)
  ) __2433__ (
    .I5(__802__),
    .I4(__327__),
    .I3(__732__),
    .I2(__291__),
    .I1(__1061__),
    .I0(__1059__),
    .O(__1062__)
  );
  LUT4 #(
    .INIT(16'hbeaa)
  ) __2434__ (
    .I3(__805__),
    .I2(__33__),
    .I1(__1062__),
    .I0(__801__),
    .O(__1063__)
  );
  LUT6 #(
    .INIT(64'hfbfa000000000000)
  ) __2435__ (
    .I5(g109),
    .I4(__247__),
    .I3(__489__),
    .I2(g881),
    .I1(__198__),
    .I0(__245__),
    .O(__1064__)
  );
  LUT4 #(
    .INIT(16'hccac)
  ) __2436__ (
    .I3(g1696),
    .I2(__11__),
    .I1(__332__),
    .I0(__76__),
    .O(__1065__)
  );
  LUT3 #(
    .INIT(8'hb0)
  ) __2437__ (
    .I2(__30__),
    .I1(g750),
    .I0(__438__),
    .O(__1066__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __2438__ (
    .I1(__500__),
    .I0(__200__),
    .O(__1067__)
  );
  LUT3 #(
    .INIT(8'h10)
  ) __2439__ (
    .I2(__112__),
    .I1(__414__),
    .I0(__273__),
    .O(__1068__)
  );
  LUT4 #(
    .INIT(16'hf013)
  ) __2440__ (
    .I3(__292__),
    .I2(__273__),
    .I1(__295__),
    .I0(__112__),
    .O(__1069__)
  );
  LUT6 #(
    .INIT(64'hfffb00aa00000000)
  ) __2441__ (
    .I5(__234__),
    .I4(__273__),
    .I3(__295__),
    .I2(__112__),
    .I1(__56__),
    .I0(__414__),
    .O(__1070__)
  );
  LUT6 #(
    .INIT(64'hf55f555511331111)
  ) __2442__ (
    .I5(__471__),
    .I4(__1070__),
    .I3(__1069__),
    .I2(__371__),
    .I1(__1068__),
    .I0(__57__),
    .O(__1071__)
  );
  LUT5 #(
    .INIT(32'hf8880000)
  ) __2443__ (
    .I4(__367__),
    .I3(__235__),
    .I2(__398__),
    .I1(__266__),
    .I0(__421__),
    .O(__1072__)
  );
  LUT6 #(
    .INIT(64'h0707ffff00ff00ff)
  ) __2444__ (
    .I5(__511__),
    .I4(__1072__),
    .I3(__1071__),
    .I2(__1067__),
    .I1(__182__),
    .I0(__439__),
    .O(__1073__)
  );
  LUT5 #(
    .INIT(32'h202a757f)
  ) __2445__ (
    .I4(__45__),
    .I3(__713__),
    .I2(__120__),
    .I1(__711__),
    .I0(__723__),
    .O(__1074__)
  );
  LUT5 #(
    .INIT(32'hfeabaaaa)
  ) __2446__ (
    .I4(__725__),
    .I3(__472__),
    .I2(__724__),
    .I1(__1074__),
    .I0(__719__),
    .O(__1075__)
  );
  LUT3 #(
    .INIT(8'hf4)
  ) __2447__ (
    .I2(__343__),
    .I1(g750),
    .I0(__438__),
    .O(__1076__)
  );
  LUT6 #(
    .INIT(64'hf0f0e2e2f0f022e2)
  ) __2448__ (
    .I5(__37__),
    .I4(__345__),
    .I3(__685__),
    .I2(__262__),
    .I1(__734__),
    .I0(__493__),
    .O(__1077__)
  );
  LUT4 #(
    .INIT(16'hbf80)
  ) __2449__ (
    .I3(__417__),
    .I2(__393__),
    .I1(__701__),
    .I0(__226__),
    .O(__1078__)
  );
  LUT3 #(
    .INIT(8'hf4)
  ) __2450__ (
    .I2(__41__),
    .I1(g750),
    .I0(__438__),
    .O(__1079__)
  );
  LUT6 #(
    .INIT(64'hefff300000000000)
  ) __2451__ (
    .I5(__996__),
    .I4(__115__),
    .I3(__104__),
    .I2(__436__),
    .I1(__679__),
    .I0(__121__),
    .O(__1080__)
  );
  LUT6 #(
    .INIT(64'h0000000080000000)
  ) __2452__ (
    .I5(__376__),
    .I4(__107__),
    .I3(__1008__),
    .I2(__48__),
    .I1(__221__),
    .I0(__239__),
    .O(__1081__)
  );
  LUT5 #(
    .INIT(32'h00000080)
  ) __2453__ (
    .I4(__244__),
    .I3(__171__),
    .I2(__322__),
    .I1(__402__),
    .I0(__135__),
    .O(__1082__)
  );
  LUT6 #(
    .INIT(64'h0000000000008000)
  ) __2454__ (
    .I5(__390__),
    .I4(__143__),
    .I3(__79__),
    .I2(__350__),
    .I1(__1082__),
    .I0(__1081__),
    .O(__1083__)
  );
  LUT3 #(
    .INIT(8'he0)
  ) __2455__ (
    .I2(g109),
    .I1(__408__),
    .I0(__1083__),
    .O(__1084__)
  );
  LUT5 #(
    .INIT(32'h65555555)
  ) __2456__ (
    .I4(__297__),
    .I3(__468__),
    .I2(__61__),
    .I1(__156__),
    .I0(__10__),
    .O(__1085__)
  );
  LUT6 #(
    .INIT(64'h8000bfffaaaaaaaa)
  ) __2457__ (
    .I5(__678__),
    .I4(__75__),
    .I3(__676__),
    .I2(__654__),
    .I1(__603__),
    .I0(__1085__),
    .O(__1086__)
  );
  LUT4 #(
    .INIT(16'ha3aa)
  ) __2458__ (
    .I3(g750),
    .I2(__438__),
    .I1(__1086__),
    .I0(__76__),
    .O(__1087__)
  );
  LUT4 #(
    .INIT(16'hb8aa)
  ) __2459__ (
    .I3(__11__),
    .I2(__474__),
    .I1(g1696),
    .I0(__248__),
    .O(__1088__)
  );
  LUT4 #(
    .INIT(16'h8000)
  ) __2460__ (
    .I3(__268__),
    .I2(__247__),
    .I1(__64__),
    .I0(__465__),
    .O(__1089__)
  );
  LUT4 #(
    .INIT(16'h0080)
  ) __2461__ (
    .I3(__11__),
    .I2(g1696),
    .I1(__53__),
    .I0(__226__),
    .O(__1090__)
  );
  LUT6 #(
    .INIT(64'h00007fff00008000)
  ) __2462__ (
    .I5(__280__),
    .I4(__154__),
    .I3(__324__),
    .I2(__116__),
    .I1(__145__),
    .I0(__1090__),
    .O(__1091__)
  );
  LUT4 #(
    .INIT(16'hf088)
  ) __2463__ (
    .I3(__508__),
    .I2(__326__),
    .I1(g109),
    .I0(__355__),
    .O(__1092__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __2464__ (
    .I2(g18),
    .I1(__185__),
    .I0(__58__),
    .O(__1093__)
  );
  LUT4 #(
    .INIT(16'h0060)
  ) __2465__ (
    .I3(__407__),
    .I2(g109),
    .I1(__453__),
    .I0(__214__),
    .O(__1094__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __2466__ (
    .I1(g109),
    .I0(__224__),
    .O(__1095__)
  );
  LUT4 #(
    .INIT(16'haab8)
  ) __2467__ (
    .I3(__11__),
    .I2(__154__),
    .I1(g1696),
    .I0(__211__),
    .O(__1096__)
  );
  LUT3 #(
    .INIT(8'h35)
  ) __2468__ (
    .I2(g18),
    .I1(__504__),
    .I0(__215__),
    .O(__1097__)
  );
  LUT6 #(
    .INIT(64'h00f5003300000000)
  ) __2469__ (
    .I5(__747__),
    .I4(__73__),
    .I3(__211__),
    .I2(__770__),
    .I1(__1097__),
    .I0(g109),
    .O(__1098__)
  );
  LUT4 #(
    .INIT(16'heeec)
  ) __2470__ (
    .I3(__11__),
    .I2(g1696),
    .I1(__1098__),
    .I0(__506__),
    .O(__1099__)
  );
  LUT5 #(
    .INIT(32'h80000000)
  ) __2471__ (
    .I4(g109),
    .I3(__49__),
    .I2(__815__),
    .I1(__813__),
    .I0(__89__),
    .O(__1100__)
  );
  LUT3 #(
    .INIT(8'h6b)
  ) __2472__ (
    .I2(__414__),
    .I1(__112__),
    .I0(__273__),
    .O(__1101__)
  );
  LUT5 #(
    .INIT(32'h8b00cfcf)
  ) __2473__ (
    .I4(__718__),
    .I3(__1101__),
    .I2(__511__),
    .I1(__715__),
    .I0(__471__),
    .O(__1102__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __2474__ (
    .I2(g18),
    .I1(__112__),
    .I0(__1102__),
    .O(__1103__)
  );
  LUT6 #(
    .INIT(64'h55555555c0003fff)
  ) __2475__ (
    .I5(g18),
    .I4(__386__),
    .I3(__400__),
    .I2(__149__),
    .I1(__767__),
    .I0(__224__),
    .O(__1104__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __2476__ (
    .I2(g109),
    .I1(__1104__),
    .I0(__240__),
    .O(__1105__)
  );
  LUT5 #(
    .INIT(32'h53ac0000)
  ) __2477__ (
    .I4(g109),
    .I3(__322__),
    .I2(g18),
    .I1(__82__),
    .I0(__224__),
    .O(__1106__)
  );
  LUT6 #(
    .INIT(64'hff00bf80aaaaaaaa)
  ) __2478__ (
    .I5(g109),
    .I4(__276__),
    .I3(__230__),
    .I2(g18),
    .I1(__212__),
    .I0(__220__),
    .O(__1107__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __2479__ (
    .I3(__11__),
    .I2(g1696),
    .I1(__43__),
    .I0(__913__),
    .O(__1108__)
  );
  LUT6 #(
    .INIT(64'h0caa0c0c0c0c0c0c)
  ) __2480__ (
    .I5(__56__),
    .I4(__512__),
    .I3(__295__),
    .I2(__511__),
    .I1(__51__),
    .I0(__319__),
    .O(__1109__)
  );
  LUT2 #(
    .INIT(4'he)
  ) __2481__ (
    .I1(g82),
    .I0(__228__),
    .O(__1110__)
  );
  LUT4 #(
    .INIT(16'hac00)
  ) __2482__ (
    .I3(g18),
    .I2(__718__),
    .I1(__414__),
    .I0(__112__),
    .O(__1111__)
  );
  LUT6 #(
    .INIT(64'h00007fff00008000)
  ) __2483__ (
    .I5(__505__),
    .I4(__154__),
    .I3(__25__),
    .I2(__280__),
    .I1(__324__),
    .I0(__968__),
    .O(__1112__)
  );
  LUT6 #(
    .INIT(64'hf0f0e2e2f0f022e2)
  ) __2484__ (
    .I5(__37__),
    .I4(__345__),
    .I3(__685__),
    .I2(__241__),
    .I1(__734__),
    .I0(__262__),
    .O(__1113__)
  );
  LUT6 #(
    .INIT(64'h300c0000aaaaaaaa)
  ) __2485__ (
    .I5(__723__),
    .I4(__717__),
    .I3(__176__),
    .I2(__67__),
    .I1(__785__),
    .I0(__319__),
    .O(__1114__)
  );
  LUT4 #(
    .INIT(16'hbeaa)
  ) __2486__ (
    .I3(__725__),
    .I2(__362__),
    .I1(__1114__),
    .I0(__719__),
    .O(__1115__)
  );
  LUT6 #(
    .INIT(64'h0caa0c0c0c0c0c0c)
  ) __2487__ (
    .I5(__56__),
    .I4(__512__),
    .I3(__295__),
    .I2(__511__),
    .I1(__352__),
    .I0(__457__),
    .O(__1116__)
  );
  LUT6 #(
    .INIT(64'h8000000000000000)
  ) __2488__ (
    .I5(__266__),
    .I4(__421__),
    .I3(__182__),
    .I2(__439__),
    .I1(__500__),
    .I0(__200__),
    .O(__1117__)
  );
  LUT5 #(
    .INIT(32'h60000000)
  ) __2489__ (
    .I4(g109),
    .I3(__278__),
    .I2(__196__),
    .I1(__398__),
    .I0(__1117__),
    .O(__1118__)
  );
  LUT6 #(
    .INIT(64'h7fff800000000000)
  ) __2490__ (
    .I5(__762__),
    .I4(__421__),
    .I3(__182__),
    .I2(__439__),
    .I1(__500__),
    .I0(__200__),
    .O(__1119__)
  );
  LUT6 #(
    .INIT(64'hff00bf80aaaaaaaa)
  ) __2491__ (
    .I5(g109),
    .I4(__276__),
    .I3(__238__),
    .I2(g18),
    .I1(__212__),
    .I0(__94__),
    .O(__1120__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __2492__ (
    .I1(g109),
    .I0(__174__),
    .O(__1121__)
  );
  LUT2 #(
    .INIT(4'h2)
  ) __2493__ (
    .I1(g1696),
    .I0(__11__),
    .O(__1122__)
  );
  LUT6 #(
    .INIT(64'h00dd0000f0f0f0f0)
  ) __2494__ (
    .I5(__1122__),
    .I4(__73__),
    .I3(__211__),
    .I2(__329__),
    .I1(__772__),
    .I0(g109),
    .O(__1123__)
  );
  LUT5 #(
    .INIT(32'h50045050)
  ) __2495__ (
    .I4(__357__),
    .I3(__166__),
    .I2(__437__),
    .I1(__216__),
    .I0(__804__),
    .O(__1124__)
  );
  LUT6 #(
    .INIT(64'hf0f0e2e2f0f0ffe2)
  ) __2496__ (
    .I5(__37__),
    .I4(__345__),
    .I3(__685__),
    .I2(__125__),
    .I1(__734__),
    .I0(__491__),
    .O(__1125__)
  );
  LUT3 #(
    .INIT(8'h35)
  ) __2497__ (
    .I2(g18),
    .I1(__225__),
    .I0(__164__),
    .O(__1126__)
  );
  LUT5 #(
    .INIT(32'hff44fff0)
  ) __2498__ (
    .I4(__73__),
    .I3(__211__),
    .I2(__1126__),
    .I1(g109),
    .I0(__675__),
    .O(__1127__)
  );
  LUT4 #(
    .INIT(16'haaa3)
  ) __2499__ (
    .I3(__11__),
    .I2(g1696),
    .I1(__1127__),
    .I0(__492__),
    .O(__1128__)
  );
  LUT4 #(
    .INIT(16'hbf80)
  ) __2500__ (
    .I3(__481__),
    .I2(__38__),
    .I1(__150__),
    .I0(__145__),
    .O(__1129__)
  );
  LUT6 #(
    .INIT(64'ha0aaa0aa606aa0aa)
  ) __2501__ (
    .I5(__56__),
    .I4(__295__),
    .I3(__720__),
    .I2(__273__),
    .I1(__718__),
    .I0(__471__),
    .O(__1130__)
  );
  LUT4 #(
    .INIT(16'hbf80)
  ) __2502__ (
    .I3(__441__),
    .I2(__11__),
    .I1(g1696),
    .I0(__565__),
    .O(__1131__)
  );
  LUT5 #(
    .INIT(32'haaaa0a08)
  ) __2503__ (
    .I4(__37__),
    .I3(__32__),
    .I2(__345__),
    .I1(__12__),
    .I0(__8__),
    .O(__1132__)
  );
  LUT4 #(
    .INIT(16'h88f0)
  ) __2504__ (
    .I3(__679__),
    .I2(__136__),
    .I1(g109),
    .I0(__7__),
    .O(__1133__)
  );
  LUT5 #(
    .INIT(32'h53ac0000)
  ) __2505__ (
    .I4(g109),
    .I3(__387__),
    .I2(g18),
    .I1(__101__),
    .I0(__424__),
    .O(__1134__)
  );
  LUT4 #(
    .INIT(16'h00cd)
  ) __2506__ (
    .I3(__37__),
    .I2(__32__),
    .I1(__345__),
    .I0(__12__),
    .O(__1135__)
  );
  LUT6 #(
    .INIT(64'hff00bf80aaaaaaaa)
  ) __2507__ (
    .I5(g109),
    .I4(__15__),
    .I3(__167__),
    .I2(g18),
    .I1(__212__),
    .I0(__240__),
    .O(__1136__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __2508__ (
    .I2(__237__),
    .I1(__453__),
    .I0(__214__),
    .O(__1137__)
  );
  LUT5 #(
    .INIT(32'h00007800)
  ) __2509__ (
    .I4(__407__),
    .I3(g109),
    .I2(__405__),
    .I1(__456__),
    .I0(__1137__),
    .O(__1138__)
  );
  LUT5 #(
    .INIT(32'haaaa0a08)
  ) __2510__ (
    .I4(__273__),
    .I3(__414__),
    .I2(__295__),
    .I1(__112__),
    .I0(__257__),
    .O(__1139__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __2511__ (
    .I1(g109),
    .I0(__419__),
    .O(__1140__)
  );
  LUT5 #(
    .INIT(32'h53ac0000)
  ) __2512__ (
    .I4(g109),
    .I3(__239__),
    .I2(g18),
    .I1(__164__),
    .I0(__225__),
    .O(__1141__)
  );
  LUT6 #(
    .INIT(64'hff8000ff00000000)
  ) __2513__ (
    .I5(__996__),
    .I4(__436__),
    .I3(__679__),
    .I2(__121__),
    .I1(__115__),
    .I0(__104__),
    .O(__1142__)
  );
  LUT4 #(
    .INIT(16'h88f0)
  ) __2514__ (
    .I3(__679__),
    .I2(__450__),
    .I1(g109),
    .I0(__423__),
    .O(__1143__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __2515__ (
    .I2(__47__),
    .I1(__395__),
    .I0(__360__),
    .O(__1144__)
  );
  LUT5 #(
    .INIT(32'haaaa0a08)
  ) __2516__ (
    .I4(__37__),
    .I3(__32__),
    .I2(__345__),
    .I1(__12__),
    .I0(__488__),
    .O(__1145__)
  );
  LUT4 #(
    .INIT(16'haaa3)
  ) __2517__ (
    .I3(__11__),
    .I2(g1696),
    .I1(__1104__),
    .I0(__451__),
    .O(__1146__)
  );
  LUT4 #(
    .INIT(16'hf088)
  ) __2518__ (
    .I3(__508__),
    .I2(__365__),
    .I1(g109),
    .I0(__334__),
    .O(__1147__)
  );
  LUT5 #(
    .INIT(32'h53ac0000)
  ) __2519__ (
    .I4(g109),
    .I3(__171__),
    .I2(g18),
    .I1(__448__),
    .I0(__392__),
    .O(__1148__)
  );
  LUT6 #(
    .INIT(64'h0033000faaaaaaaa)
  ) __2520__ (
    .I5(__747__),
    .I4(__73__),
    .I3(__211__),
    .I2(__760__),
    .I1(__759__),
    .I0(__103__),
    .O(__1149__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __2521__ (
    .I3(__11__),
    .I2(g1696),
    .I1(__300__),
    .I0(__843__),
    .O(__1150__)
  );
  LUT3 #(
    .INIT(8'h60)
  ) __2522__ (
    .I2(g1700),
    .I1(__47__),
    .I0(__284__),
    .O(__1151__)
  );
  LUT4 #(
    .INIT(16'h88f0)
  ) __2523__ (
    .I3(__679__),
    .I2(__157__),
    .I1(g109),
    .I0(__96__),
    .O(__1152__)
  );
  LUT6 #(
    .INIT(64'h000000007f800000)
  ) __2524__ (
    .I5(__407__),
    .I4(g109),
    .I3(__456__),
    .I2(__237__),
    .I1(__453__),
    .I0(__214__),
    .O(__1153__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __2525__ (
    .I1(g109),
    .I0(__20__),
    .O(__1154__)
  );
  LUT6 #(
    .INIT(64'hff00bf80aaaaaaaa)
  ) __2526__ (
    .I5(g109),
    .I4(__15__),
    .I3(__366__),
    .I2(g18),
    .I1(__212__),
    .I0(__322__),
    .O(__1155__)
  );
  LUT3 #(
    .INIT(8'hb0)
  ) __2527__ (
    .I2(__265__),
    .I1(g1696),
    .I0(__11__),
    .O(__1156__)
  );
  LUT6 #(
    .INIT(64'hff00bf80aaaaaaaa)
  ) __2528__ (
    .I5(g109),
    .I4(__15__),
    .I3(__66__),
    .I2(g18),
    .I1(__212__),
    .I0(__402__),
    .O(__1157__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __2529__ (
    .I1(g109),
    .I0(__70__),
    .O(__1158__)
  );
  LUT5 #(
    .INIT(32'h007f0080)
  ) __2530__ (
    .I4(__25__),
    .I3(__154__),
    .I2(__280__),
    .I1(__324__),
    .I0(__968__),
    .O(__1159__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __2531__ (
    .I3(__11__),
    .I2(g1696),
    .I1(__9__),
    .I0(__358__),
    .O(__1160__)
  );
  LUT6 #(
    .INIT(64'h33bfcc0000000000)
  ) __2532__ (
    .I5(g18),
    .I4(__345__),
    .I3(__478__),
    .I2(__37__),
    .I1(__686__),
    .I0(__733__),
    .O(__1161__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __2533__ (
    .I1(g109),
    .I0(__161__),
    .O(__1162__)
  );
  LUT6 #(
    .INIT(64'h0caa0c0c0c0c0c0c)
  ) __2534__ (
    .I5(__56__),
    .I4(__512__),
    .I3(__295__),
    .I2(__511__),
    .I1(__319__),
    .I0(__464__),
    .O(__1163__)
  );
  LUT6 #(
    .INIT(64'hff00bf80aaaaaaaa)
  ) __2535__ (
    .I5(g109),
    .I4(__15__),
    .I3(__133__),
    .I2(g18),
    .I1(__212__),
    .I0(__210__),
    .O(__1164__)
  );
  LUT4 #(
    .INIT(16'haaa3)
  ) __2536__ (
    .I3(__11__),
    .I2(g1696),
    .I1(__756__),
    .I0(__389__),
    .O(__1165__)
  );
  LUT4 #(
    .INIT(16'h0bff)
  ) __2537__ (
    .I3(g109),
    .I2(__320__),
    .I1(__106__),
    .I0(__170__),
    .O(__1166__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __2538__ (
    .I2(__505__),
    .I1(__144__),
    .I0(__145__),
    .O(__1167__)
  );
  LUT4 #(
    .INIT(16'h8000)
  ) __2539__ (
    .I3(__53__),
    .I2(__226__),
    .I1(__47__),
    .I0(__284__),
    .O(__1168__)
  );
  LUT6 #(
    .INIT(64'h0000000080000000)
  ) __2540__ (
    .I5(__116__),
    .I4(__25__),
    .I3(__280__),
    .I2(__324__),
    .I1(__1168__),
    .I0(__1167__),
    .O(__1169__)
  );
  LUT6 #(
    .INIT(64'hff00f870ff00ff00)
  ) __2541__ (
    .I5(__680__),
    .I4(__519__),
    .I3(__126__),
    .I2(__485__),
    .I1(g109),
    .I0(__380__),
    .O(__1170__)
  );
  LUT4 #(
    .INIT(16'h88f0)
  ) __2542__ (
    .I3(__679__),
    .I2(__208__),
    .I1(g109),
    .I0(__162__),
    .O(__1171__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __2543__ (
    .I1(__11__),
    .I0(g1696),
    .O(__1172__)
  );
  LUT6 #(
    .INIT(64'hdfff8aaaffffaaaa)
  ) __2544__ (
    .I5(g109),
    .I4(__209__),
    .I3(__619__),
    .I2(__612__),
    .I1(__607__),
    .I0(__1172__),
    .O(__1173__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __2545__ (
    .I1(g109),
    .I0(__390__),
    .O(__1174__)
  );
  LUT6 #(
    .INIT(64'haaaafcccaaaaaaaa)
  ) __2546__ (
    .I5(__11__),
    .I4(g1696),
    .I3(__585__),
    .I2(__73__),
    .I1(__211__),
    .I0(__181__),
    .O(__1175__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __2547__ (
    .I1(g109),
    .I0(__483__),
    .O(__1176__)
  );
  LUT4 #(
    .INIT(16'h7fff)
  ) __2548__ (
    .I3(g109),
    .I2(__278__),
    .I1(__196__),
    .I0(__200__),
    .O(__1177__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __2549__ (
    .I1(g109),
    .I0(__138__),
    .O(__1178__)
  );
  LUT6 #(
    .INIT(64'hffff400000000000)
  ) __2550__ (
    .I5(__1178__),
    .I4(__156__),
    .I3(__297__),
    .I2(__468__),
    .I1(__61__),
    .I0(__679__),
    .O(__1179__)
  );
  LUT6 #(
    .INIT(64'hff00bf80aaaaaaaa)
  ) __2551__ (
    .I5(g109),
    .I4(__276__),
    .I3(__323__),
    .I2(g18),
    .I1(__212__),
    .I0(__476__),
    .O(__1180__)
  );
  LUT4 #(
    .INIT(16'h0060)
  ) __2552__ (
    .I3(__383__),
    .I2(g1700),
    .I1(__11__),
    .I0(g1696),
    .O(__1181__)
  );
  LUT5 #(
    .INIT(32'h53ac0000)
  ) __2553__ (
    .I4(g109),
    .I3(__221__),
    .I2(g18),
    .I1(__389__),
    .I0(__424__),
    .O(__1182__)
  );
  LUT6 #(
    .INIT(64'hd1d1d11d1d1d1dd1)
  ) __2554__ (
    .I5(__414__),
    .I4(__112__),
    .I3(__273__),
    .I2(__176__),
    .I1(__723__),
    .I0(__464__),
    .O(__1183__)
  );
  LUT5 #(
    .INIT(32'hfeabaaaa)
  ) __2555__ (
    .I4(__725__),
    .I3(__67__),
    .I2(__724__),
    .I1(__1183__),
    .I0(__719__),
    .O(__1184__)
  );
  LUT4 #(
    .INIT(16'hccca)
  ) __2556__ (
    .I3(__11__),
    .I2(g1696),
    .I1(__463__),
    .I0(__412__),
    .O(__1185__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __2557__ (
    .I1(g109),
    .I0(__22__),
    .O(__1186__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __2558__ (
    .I1(g109),
    .I0(__325__),
    .O(__1187__)
  );
  LUT4 #(
    .INIT(16'hbf80)
  ) __2559__ (
    .I3(__190__),
    .I2(__38__),
    .I1(__150__),
    .I0(__25__),
    .O(__1188__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __2560__ (
    .I1(g109),
    .I0(__194__),
    .O(__1189__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __2561__ (
    .I2(g18),
    .I1(__392__),
    .I0(__142__),
    .O(__1190__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __2562__ (
    .I3(__11__),
    .I2(g1696),
    .I1(__207__),
    .I0(__461__),
    .O(__1191__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __2563__ (
    .I1(__297__),
    .I0(__468__),
    .O(__1192__)
  );
  LUT6 #(
    .INIT(64'h00000000ef300000)
  ) __2564__ (
    .I5(__138__),
    .I4(g109),
    .I3(__61__),
    .I2(__1192__),
    .I1(__679__),
    .I0(__156__),
    .O(__1193__)
  );
  LUT4 #(
    .INIT(16'haaa3)
  ) __2565__ (
    .I3(__11__),
    .I2(g1696),
    .I1(__963__),
    .I0(__395__),
    .O(__1194__)
  );
  LUT4 #(
    .INIT(16'hccca)
  ) __2566__ (
    .I3(__11__),
    .I2(g1696),
    .I1(__260__),
    .I0(__248__),
    .O(__1195__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __2567__ (
    .I3(__11__),
    .I2(g1696),
    .I1(__137__),
    .I0(__86__),
    .O(__1196__)
  );
  LUT5 #(
    .INIT(32'h7fff8000)
  ) __2568__ (
    .I4(__407__),
    .I3(__378__),
    .I2(__497__),
    .I1(__683__),
    .I0(__42__),
    .O(__1197__)
  );
  LUT6 #(
    .INIT(64'h7fff800000000000)
  ) __2569__ (
    .I5(__799__),
    .I4(__404__),
    .I3(__458__),
    .I2(__39__),
    .I1(__344__),
    .I0(__680__),
    .O(__1198__)
  );
  LUT4 #(
    .INIT(16'h88f0)
  ) __2570__ (
    .I3(__679__),
    .I2(__7__),
    .I1(g109),
    .I0(__399__),
    .O(__1199__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __2571__ (
    .I1(g109),
    .I0(__225__),
    .O(__1200__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __2572__ (
    .I1(g109),
    .I0(__433__),
    .O(__1201__)
  );
  LUT6 #(
    .INIT(64'hbfc03fc000000000)
  ) __2573__ (
    .I5(__1201__),
    .I4(__201__),
    .I3(__98__),
    .I2(__14__),
    .I1(__508__),
    .I0(__411__),
    .O(__1202__)
  );
  LUT6 #(
    .INIT(64'hff00bf80aaaaaaaa)
  ) __2574__ (
    .I5(g109),
    .I4(__276__),
    .I3(__482__),
    .I2(g18),
    .I1(__212__),
    .I0(__70__),
    .O(__1203__)
  );
  LUT4 #(
    .INIT(16'hccca)
  ) __2575__ (
    .I3(__11__),
    .I2(g1696),
    .I1(__141__),
    .I0(__455__),
    .O(__1204__)
  );
  LUT4 #(
    .INIT(16'h0bff)
  ) __2576__ (
    .I3(g109),
    .I2(g881),
    .I1(__489__),
    .I0(__198__),
    .O(__1205__)
  );
  LUT3 #(
    .INIT(8'hf4)
  ) __2577__ (
    .I2(__351__),
    .I1(g750),
    .I0(__438__),
    .O(__1206__)
  );
  LUT6 #(
    .INIT(64'hff00f870ff00ff00)
  ) __2578__ (
    .I5(__680__),
    .I4(__519__),
    .I3(__298__),
    .I2(__124__),
    .I1(g109),
    .I0(__380__),
    .O(__1207__)
  );
  LUT5 #(
    .INIT(32'hfffeffff)
  ) __2579__ (
    .I4(g48),
    .I3(g41),
    .I2(g30),
    .I1(g31),
    .I0(__664__),
    .O(__1208__)
  );
  LUT3 #(
    .INIT(8'h40)
  ) __2580__ (
    .I2(g109),
    .I1(__149__),
    .I0(__183__),
    .O(__1209__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __2581__ (
    .I1(g109),
    .I0(__277__),
    .O(__1210__)
  );
  LUT4 #(
    .INIT(16'heeec)
  ) __2582__ (
    .I3(__11__),
    .I2(g1696),
    .I1(__1098__),
    .I0(__305__),
    .O(__1211__)
  );
  LUT4 #(
    .INIT(16'hf088)
  ) __2583__ (
    .I3(__508__),
    .I2(__68__),
    .I1(g109),
    .I0(__255__),
    .O(__1212__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __2584__ (
    .I1(g109),
    .I0(__424__),
    .O(__1213__)
  );
  LUT4 #(
    .INIT(16'hbf80)
  ) __2585__ (
    .I3(__160__),
    .I2(__393__),
    .I1(__701__),
    .I0(__144__),
    .O(__1214__)
  );
  LUT3 #(
    .INIT(8'h04)
  ) __2586__ (
    .I2(g1696),
    .I1(g1700),
    .I0(__383__),
    .O(__1215__)
  );
  LUT6 #(
    .INIT(64'hffd0ff20ff10ffe0)
  ) __2587__ (
    .I5(__732__),
    .I4(__60__),
    .I3(__801__),
    .I2(__805__),
    .I1(__802__),
    .I0(__125__),
    .O(__1216__)
  );
  LUT2 #(
    .INIT(4'he)
  ) __2588__ (
    .I1(g82),
    .I0(__351__),
    .O(__1217__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __2589__ (
    .I1(g109),
    .I0(__392__),
    .O(__1218__)
  );
  LUT3 #(
    .INIT(8'hc1)
  ) __2590__ (
    .I2(__55__),
    .I1(__341__),
    .I0(__709__),
    .O(__1219__)
  );
  LUT5 #(
    .INIT(32'h55555559)
  ) __2591__ (
    .I4(__468__),
    .I3(__61__),
    .I2(__156__),
    .I1(__297__),
    .I0(__1219__),
    .O(__1220__)
  );
  LUT6 #(
    .INIT(64'h5333333355555555)
  ) __2592__ (
    .I5(__678__),
    .I4(__676__),
    .I3(__654__),
    .I2(__603__),
    .I1(__340__),
    .I0(__1220__),
    .O(__1221__)
  );
  LUT5 #(
    .INIT(32'h55555559)
  ) __2593__ (
    .I4(__297__),
    .I3(__61__),
    .I2(__156__),
    .I1(__468__),
    .I0(__339__),
    .O(__1222__)
  );
  LUT6 #(
    .INIT(64'h8000bfffaaaaaaaa)
  ) __2594__ (
    .I5(__678__),
    .I4(__369__),
    .I3(__676__),
    .I2(__654__),
    .I1(__603__),
    .I0(__1222__),
    .O(__1223__)
  );
  LUT6 #(
    .INIT(64'ha35c5ca35ca3a35c)
  ) __2595__ (
    .I5(__1223__),
    .I4(__982__),
    .I3(__889__),
    .I2(__679__),
    .I1(__884__),
    .I0(__496__),
    .O(__1224__)
  );
  LUT6 #(
    .INIT(64'h5ca3a35ca35c5ca3)
  ) __2596__ (
    .I5(__834__),
    .I4(__1086__),
    .I3(__1021__),
    .I2(__679__),
    .I1(__1036__),
    .I0(__123__),
    .O(__1225__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __2597__ (
    .I1(g750),
    .I0(__438__),
    .O(__1226__)
  );
  LUT6 #(
    .INIT(64'h3cc3c33caaaaaaaa)
  ) __2598__ (
    .I5(__1226__),
    .I4(__781__),
    .I3(__1225__),
    .I2(__1224__),
    .I1(__1221__),
    .I0(__54__),
    .O(__1227__)
  );
  LUT3 #(
    .INIT(8'h40)
  ) __2599__ (
    .I2(g109),
    .I1(__222__),
    .I0(__183__),
    .O(__1228__)
  );
  LUT6 #(
    .INIT(64'hfbfa000000000000)
  ) __2600__ (
    .I5(g109),
    .I4(__64__),
    .I3(__489__),
    .I2(g881),
    .I1(__198__),
    .I0(__245__),
    .O(__1229__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __2601__ (
    .I2(g18),
    .I1(__174__),
    .I0(__103__),
    .O(__1230__)
  );
  LUT6 #(
    .INIT(64'hff00bf80aaaaaaaa)
  ) __2602__ (
    .I5(g109),
    .I4(__15__),
    .I3(__435__),
    .I2(g18),
    .I1(__212__),
    .I0(__148__),
    .O(__1231__)
  );
  LUT4 #(
    .INIT(16'h88f0)
  ) __2603__ (
    .I3(__679__),
    .I2(__339__),
    .I1(g109),
    .I0(__157__),
    .O(__1232__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __2604__ (
    .I1(g109),
    .I0(__494__),
    .O(__1233__)
  );
  LUT4 #(
    .INIT(16'ha3aa)
  ) __2605__ (
    .I3(__11__),
    .I2(g1696),
    .I1(__790__),
    .I0(__360__),
    .O(__1234__)
  );
  LUT6 #(
    .INIT(64'hff00bf80aaaaaaaa)
  ) __2606__ (
    .I5(g109),
    .I4(__15__),
    .I3(__486__),
    .I2(g18),
    .I1(__212__),
    .I0(__239__),
    .O(__1235__)
  );
  LUT6 #(
    .INIT(64'haaaaffffffffaaaa)
  ) __2607__ (
    .I5(__118__),
    .I4(__333__),
    .I3(__309__),
    .I2(__261__),
    .I1(__269__),
    .I0(__511__),
    .O(__1236__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __2608__ (
    .I1(g109),
    .I0(__350__),
    .O(__1237__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __2609__ (
    .I1(g109),
    .I0(__256__),
    .O(__1238__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __2610__ (
    .I1(__150__),
    .I0(__418__),
    .O(__1239__)
  );
  LUT4 #(
    .INIT(16'h00e0)
  ) __2611__ (
    .I3(__212__),
    .I2(g109),
    .I1(__89__),
    .I0(__381__),
    .O(__1240__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __2612__ (
    .I3(__11__),
    .I2(g1696),
    .I1(__455__),
    .I0(__475__),
    .O(__1241__)
  );
  LUT5 #(
    .INIT(32'h53ac0000)
  ) __2613__ (
    .I4(g109),
    .I3(__402__),
    .I2(g18),
    .I1(__283__),
    .I0(__494__),
    .O(__1242__)
  );
  LUT6 #(
    .INIT(64'h0caa0c0c0c0c0c0c)
  ) __2614__ (
    .I5(__56__),
    .I4(__512__),
    .I3(__295__),
    .I2(__511__),
    .I1(__416__),
    .I0(__352__),
    .O(__1243__)
  );
  LUT3 #(
    .INIT(8'hf4)
  ) __2615__ (
    .I2(__3__),
    .I1(g750),
    .I0(__438__),
    .O(__1244__)
  );
  LUT3 #(
    .INIT(8'hb0)
  ) __2616__ (
    .I2(__349__),
    .I1(g750),
    .I0(__438__),
    .O(__1245__)
  );
  LUT4 #(
    .INIT(16'hccca)
  ) __2617__ (
    .I3(__11__),
    .I2(g1696),
    .I1(__206__),
    .I0(__137__),
    .O(__1246__)
  );
  LUT3 #(
    .INIT(8'hb0)
  ) __2618__ (
    .I2(__353__),
    .I1(g750),
    .I0(__438__),
    .O(__1247__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __2619__ (
    .I1(g109),
    .I0(__49__),
    .O(__1248__)
  );
  LUT6 #(
    .INIT(64'hfffffffffffffffd)
  ) __2620__ (
    .I5(g48),
    .I4(g42),
    .I3(g44),
    .I2(g45),
    .I1(g43),
    .I0(__538__),
    .O(__1249__)
  );
  LUT4 #(
    .INIT(16'h88f0)
  ) __2621__ (
    .I3(__679__),
    .I2(__6__),
    .I1(g109),
    .I0(__335__),
    .O(__1250__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __2622__ (
    .I2(__47__),
    .I1(__218__),
    .I0(__300__),
    .O(__1251__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __2623__ (
    .I1(g109),
    .I0(__185__),
    .O(__1252__)
  );
  LUT5 #(
    .INIT(32'h53ac0000)
  ) __2624__ (
    .I4(g109),
    .I3(__48__),
    .I2(g18),
    .I1(__374__),
    .I0(__174__),
    .O(__1253__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __2625__ (
    .I1(g109),
    .I0(__83__),
    .O(__1254__)
  );
  LUT6 #(
    .INIT(64'h03000030aaaaaaaa)
  ) __2626__ (
    .I5(__802__),
    .I4(__60__),
    .I3(__503__),
    .I2(__1060__),
    .I1(__732__),
    .I0(__262__),
    .O(__1255__)
  );
  LUT4 #(
    .INIT(16'hbeaa)
  ) __2627__ (
    .I3(__805__),
    .I2(__110__),
    .I1(__1255__),
    .I0(__801__),
    .O(__1256__)
  );
  LUT4 #(
    .INIT(16'h88f0)
  ) __2628__ (
    .I3(__679__),
    .I2(__499__),
    .I1(g109),
    .I0(__420__),
    .O(__1257__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __2629__ (
    .I2(__47__),
    .I1(__434__),
    .I0(__43__),
    .O(__1258__)
  );
  LUT2 #(
    .INIT(4'he)
  ) __2630__ (
    .I1(g82),
    .I0(__313__),
    .O(__1259__)
  );
  LUT6 #(
    .INIT(64'hffff800000000000)
  ) __2631__ (
    .I5(__1201__),
    .I4(__411__),
    .I3(__201__),
    .I2(__98__),
    .I1(__14__),
    .I0(__508__),
    .O(__1260__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __2632__ (
    .I1(g109),
    .I0(__148__),
    .O(__1261__)
  );
  LUT6 #(
    .INIT(64'h0f030003aaaaaaaa)
  ) __2633__ (
    .I5(__747__),
    .I4(__954__),
    .I3(__73__),
    .I2(__211__),
    .I1(__1048__),
    .I0(__413__),
    .O(__1262__)
  );
  LUT6 #(
    .INIT(64'h55ffff330f0f0f0f)
  ) __2634__ (
    .I5(__723__),
    .I4(__472__),
    .I3(__328__),
    .I2(__352__),
    .I1(__786__),
    .I0(__784__),
    .O(__1263__)
  );
  LUT5 #(
    .INIT(32'hfeabaaaa)
  ) __2635__ (
    .I4(__725__),
    .I3(__490__),
    .I2(__1263__),
    .I1(__724__),
    .I0(__719__),
    .O(__1264__)
  );
  LUT3 #(
    .INIT(8'hb0)
  ) __2636__ (
    .I2(__422__),
    .I1(g1696),
    .I0(__11__),
    .O(__1265__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __2637__ (
    .I1(g109),
    .I0(__354__),
    .O(__1266__)
  );
  LUT6 #(
    .INIT(64'hff00bf80aaaaaaaa)
  ) __2638__ (
    .I5(g109),
    .I4(__15__),
    .I3(__477__),
    .I2(g18),
    .I1(__212__),
    .I0(__221__),
    .O(__1267__)
  );
  LUT6 #(
    .INIT(64'hfffffffffffdffff)
  ) __2639__ (
    .I5(g48),
    .I4(g42),
    .I3(g44),
    .I2(g45),
    .I1(g43),
    .I0(__541__),
    .O(__1268__)
  );
  LUT4 #(
    .INIT(16'hbf80)
  ) __2640__ (
    .I3(__431__),
    .I2(__11__),
    .I1(g1696),
    .I0(__602__),
    .O(__1269__)
  );
  LUT5 #(
    .INIT(32'hf0008888)
  ) __2641__ (
    .I4(__47__),
    .I3(__770__),
    .I2(__917__),
    .I1(__280__),
    .I0(__324__),
    .O(__1270__)
  );
  LUT6 #(
    .INIT(64'h00000fff00007777)
  ) __2642__ (
    .I5(__47__),
    .I4(__1270__),
    .I3(__675__),
    .I2(__664__),
    .I1(__505__),
    .I0(__25__),
    .O(__1271__)
  );
  LUT5 #(
    .INIT(32'hf0008888)
  ) __2643__ (
    .I4(__47__),
    .I3(__774__),
    .I2(__772__),
    .I1(__116__),
    .I0(__145__),
    .O(__1272__)
  );
  LUT6 #(
    .INIT(64'h00000fff00007777)
  ) __2644__ (
    .I5(__47__),
    .I4(__1272__),
    .I3(__745__),
    .I2(__773__),
    .I1(__53__),
    .I0(__226__),
    .O(__1273__)
  );
  LUT6 #(
    .INIT(64'hfcfcfcfc0055ff00)
  ) __2645__ (
    .I5(__804__),
    .I4(__686__),
    .I3(__429__),
    .I2(__1273__),
    .I1(__1271__),
    .I0(__685__),
    .O(__1274__)
  );
  LUT6 #(
    .INIT(64'hbc3c3c3c00000000)
  ) __2646__ (
    .I5(__1201__),
    .I4(__201__),
    .I3(__98__),
    .I2(__14__),
    .I1(__508__),
    .I0(__411__),
    .O(__1275__)
  );
  LUT6 #(
    .INIT(64'hff00bf80aaaaaaaa)
  ) __2647__ (
    .I5(g109),
    .I4(__15__),
    .I3(__306__),
    .I2(g18),
    .I1(__212__),
    .I0(__244__),
    .O(__1276__)
  );
  LUT6 #(
    .INIT(64'hf8ff0f0000000000)
  ) __2648__ (
    .I5(__1178__),
    .I4(__468__),
    .I3(__297__),
    .I2(__679__),
    .I1(__61__),
    .I0(__156__),
    .O(__1277__)
  );
  LUT6 #(
    .INIT(64'hfffffffffffffffd)
  ) __2649__ (
    .I5(g48),
    .I4(g42),
    .I3(g44),
    .I2(g45),
    .I1(g43),
    .I0(__541__),
    .O(__1278__)
  );
  LUT5 #(
    .INIT(32'h00000004)
  ) __2650__ (
    .I4(__32__),
    .I3(__345__),
    .I2(__478__),
    .I1(__37__),
    .I0(__12__),
    .O(__1279__)
  );
  LUT3 #(
    .INIT(8'h40)
  ) __2651__ (
    .I2(__37__),
    .I1(__345__),
    .I0(__478__),
    .O(__1280__)
  );
  LUT6 #(
    .INIT(64'h00ff00ff00ff45ff)
  ) __2652__ (
    .I5(__478__),
    .I4(__1280__),
    .I3(__686__),
    .I2(__429__),
    .I1(__685__),
    .I0(__1279__),
    .O(__1281__)
  );
  LUT6 #(
    .INIT(64'h55ffff330f0f0f0f)
  ) __2653__ (
    .I5(__802__),
    .I4(__327__),
    .I3(__33__),
    .I2(__391__),
    .I1(__1061__),
    .I0(__1059__),
    .O(__1282__)
  );
  LUT5 #(
    .INIT(32'hfeabaaaa)
  ) __2654__ (
    .I4(__805__),
    .I3(__363__),
    .I2(__1282__),
    .I1(__1281__),
    .I0(__801__),
    .O(__1283__)
  );
  LUT3 #(
    .INIT(8'h60)
  ) __2655__ (
    .I2(__702__),
    .I1(__701__),
    .I0(__336__),
    .O(__1284__)
  );
  LUT3 #(
    .INIT(8'hb0)
  ) __2656__ (
    .I2(__313__),
    .I1(g750),
    .I0(__438__),
    .O(__1285__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __2657__ (
    .I1(__694__),
    .I0(__675__),
    .O(__1286__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __2658__ (
    .I1(__23__),
    .I0(__186__),
    .O(__1287__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __2659__ (
    .I1(__260__),
    .I0(__251__),
    .O(__1288__)
  );
  LUT6 #(
    .INIT(64'h9669699669969669)
  ) __2660__ (
    .I5(__219__),
    .I4(__206__),
    .I3(__141__),
    .I2(__293__),
    .I1(__1288__),
    .I0(__1287__),
    .O(__1289__)
  );
  LUT6 #(
    .INIT(64'hcffcfccfaaaaaaaa)
  ) __2661__ (
    .I5(__747__),
    .I4(__314__),
    .I3(__250__),
    .I2(__1289__),
    .I1(__1286__),
    .I0(__146__),
    .O(__1290__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __2662__ (
    .I2(g109),
    .I1(__382__),
    .I0(__817__),
    .O(__1291__)
  );
  LUT4 #(
    .INIT(16'ha3aa)
  ) __2663__ (
    .I3(g750),
    .I2(__438__),
    .I1(__1223__),
    .I0(__330__),
    .O(__1292__)
  );
  LUT6 #(
    .INIT(64'hffff400000000000)
  ) __2664__ (
    .I5(__996__),
    .I4(__121__),
    .I3(__115__),
    .I2(__104__),
    .I1(__436__),
    .I0(__679__),
    .O(__1293__)
  );
  LUT6 #(
    .INIT(64'h7800000000000000)
  ) __2665__ (
    .I5(g109),
    .I4(__278__),
    .I3(__196__),
    .I2(__235__),
    .I1(__398__),
    .I0(__1117__),
    .O(__1294__)
  );
  LUT6 #(
    .INIT(64'hff00bf80aaaaaaaa)
  ) __2666__ (
    .I5(g109),
    .I4(__276__),
    .I3(__84__),
    .I2(g18),
    .I1(__212__),
    .I0(__372__),
    .O(__1295__)
  );
  LUT6 #(
    .INIT(64'hefffffffffffffff)
  ) __2667__ (
    .I5(g48),
    .I4(__636__),
    .I3(__627__),
    .I2(__622__),
    .I1(__938__),
    .I0(__547__),
    .O(__1296__)
  );
  LUT4 #(
    .INIT(16'h88f0)
  ) __2668__ (
    .I3(__679__),
    .I2(__347__),
    .I1(g109),
    .I0(__165__),
    .O(__1297__)
  );
  LUT4 #(
    .INIT(16'hbf80)
  ) __2669__ (
    .I3(__108__),
    .I2(__38__),
    .I1(__150__),
    .I0(__280__),
    .O(__1298__)
  );
  LUT3 #(
    .INIT(8'he0)
  ) __2670__ (
    .I2(__73__),
    .I1(__11__),
    .I0(g1696),
    .O(__1299__)
  );
  LUT4 #(
    .INIT(16'hbf80)
  ) __2671__ (
    .I3(__285__),
    .I2(__38__),
    .I1(__150__),
    .I0(__505__),
    .O(__1300__)
  );
  LUT6 #(
    .INIT(64'h0000000000000004)
  ) __2672__ (
    .I5(__1017__),
    .I4(__1016__),
    .I3(__1015__),
    .I2(__1014__),
    .I1(__1056__),
    .I0(__1013__),
    .O(__1301__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __2673__ (
    .I2(g18),
    .I1(__44__),
    .I0(__204__),
    .O(__1302__)
  );
  LUT4 #(
    .INIT(16'ha3aa)
  ) __2674__ (
    .I3(__11__),
    .I2(g1696),
    .I1(__1127__),
    .I0(__270__),
    .O(__1303__)
  );
  LUT6 #(
    .INIT(64'h7ffffffc7fffffff)
  ) __2675__ (
    .I5(__713__),
    .I4(__120__),
    .I3(__472__),
    .I2(__328__),
    .I1(__490__),
    .I0(__711__),
    .O(__1304__)
  );
  LUT4 #(
    .INIT(16'h44f0)
  ) __2676__ (
    .I3(__723__),
    .I2(__416__),
    .I1(__717__),
    .I0(__1304__),
    .O(__1305__)
  );
  LUT4 #(
    .INIT(16'hbeaa)
  ) __2677__ (
    .I3(__725__),
    .I2(__77__),
    .I1(__1305__),
    .I0(__719__),
    .O(__1306__)
  );
  LUT4 #(
    .INIT(16'hf088)
  ) __2678__ (
    .I3(__508__),
    .I2(__334__),
    .I1(g109),
    .I0(__179__),
    .O(__1307__)
  );
  LUT2 #(
    .INIT(4'he)
  ) __2679__ (
    .I1(g82),
    .I0(__349__),
    .O(__1308__)
  );
  LUT4 #(
    .INIT(16'hf800)
  ) __2680__ (
    .I3(g109),
    .I2(__129__),
    .I1(g18),
    .I0(__212__),
    .O(__1309__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __2681__ (
    .I1(g109),
    .I0(__487__),
    .O(__1310__)
  );
  LUT4 #(
    .INIT(16'h8000)
  ) __2682__ (
    .I3(__469__),
    .I2(__336__),
    .I1(__427__),
    .I0(__90__),
    .O(__1311__)
  );
  LUT6 #(
    .INIT(64'hf00707f007f0f007)
  ) __2683__ (
    .I5(__302__),
    .I4(__415__),
    .I3(__289__),
    .I2(__49__),
    .I1(__815__),
    .I0(__813__),
    .O(__1312__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __2684__ (
    .I1(g109),
    .I0(__1312__),
    .O(__1313__)
  );
  LUT6 #(
    .INIT(64'h5050500450505050)
  ) __2685__ (
    .I5(__118__),
    .I4(__333__),
    .I3(__309__),
    .I2(__261__),
    .I1(__269__),
    .I0(__511__),
    .O(__1314__)
  );
  LUT3 #(
    .INIT(8'hb0)
  ) __2686__ (
    .I2(__254__),
    .I1(g750),
    .I0(__438__),
    .O(__1315__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __2687__ (
    .I1(g109),
    .I0(__92__),
    .O(__1316__)
  );
  LUT6 #(
    .INIT(64'hff00f870ff00ff00)
  ) __2688__ (
    .I5(__680__),
    .I4(__519__),
    .I3(__462__),
    .I2(__394__),
    .I1(g109),
    .I0(__380__),
    .O(__1317__)
  );
  LUT6 #(
    .INIT(64'h7ffffffc7fffffff)
  ) __2689__ (
    .I5(__728__),
    .I4(__479__),
    .I3(__327__),
    .I2(__363__),
    .I1(__33__),
    .I0(__730__),
    .O(__1318__)
  );
  LUT6 #(
    .INIT(64'hfc0355aa00000000)
  ) __2690__ (
    .I5(__805__),
    .I4(__802__),
    .I3(__189__),
    .I2(__732__),
    .I1(__1318__),
    .I0(__446__),
    .O(__1319__)
  );
  LUT2 #(
    .INIT(4'he)
  ) __2691__ (
    .I1(__801__),
    .I0(__1319__),
    .O(__1320__)
  );
  LUT5 #(
    .INIT(32'hfffeffff)
  ) __2692__ (
    .I4(g48),
    .I3(g41),
    .I2(g30),
    .I1(g31),
    .I0(__745__),
    .O(__1321__)
  );
  LUT5 #(
    .INIT(32'h00007800)
  ) __2693__ (
    .I4(__407__),
    .I3(g109),
    .I2(__378__),
    .I1(__497__),
    .I0(__683__),
    .O(__1322__)
  );
  LUT5 #(
    .INIT(32'haaaa0a08)
  ) __2694__ (
    .I4(__273__),
    .I3(__414__),
    .I2(__295__),
    .I1(__112__),
    .I0(__234__),
    .O(__1323__)
  );
  LUT4 #(
    .INIT(16'heeec)
  ) __2695__ (
    .I3(__11__),
    .I2(g1696),
    .I1(__748__),
    .I0(__348__),
    .O(__1324__)
  );
  LUT6 #(
    .INIT(64'hff00f870ff00ff00)
  ) __2696__ (
    .I5(__680__),
    .I4(__519__),
    .I3(__26__),
    .I2(__299__),
    .I1(g109),
    .I0(__380__),
    .O(__1325__)
  );
  LUT6 #(
    .INIT(64'h555555553000cfff)
  ) __2697__ (
    .I5(g18),
    .I4(__161__),
    .I3(__400__),
    .I2(__516__),
    .I1(__149__),
    .I0(__185__),
    .O(__1326__)
  );
  LUT4 #(
    .INIT(16'haaa3)
  ) __2698__ (
    .I3(__11__),
    .I2(g1696),
    .I1(__1326__),
    .I0(__215__),
    .O(__1327__)
  );
  LUT4 #(
    .INIT(16'h88f0)
  ) __2699__ (
    .I3(__679__),
    .I2(__272__),
    .I1(g109),
    .I0(__499__),
    .O(__1328__)
  );
  LUT6 #(
    .INIT(64'hff00f870ff00ff00)
  ) __2700__ (
    .I5(__680__),
    .I4(__519__),
    .I3(__384__),
    .I2(__169__),
    .I1(g109),
    .I0(__380__),
    .O(__1329__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __2701__ (
    .I3(__11__),
    .I2(g1696),
    .I1(__473__),
    .I0(__311__),
    .O(__1330__)
  );
  LUT5 #(
    .INIT(32'h53ac0000)
  ) __2702__ (
    .I4(g109),
    .I3(__105__),
    .I2(g18),
    .I1(__103__),
    .I0(__174__),
    .O(__1331__)
  );
  LUT6 #(
    .INIT(64'hff00bf80aaaaaaaa)
  ) __2703__ (
    .I5(g109),
    .I4(__15__),
    .I3(__4__),
    .I2(g18),
    .I1(__212__),
    .I0(__217__),
    .O(__1332__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __2704__ (
    .I1(__324__),
    .I0(__968__),
    .O(__1333__)
  );
  LUT6 #(
    .INIT(64'h00007fff00008000)
  ) __2705__ (
    .I5(__144__),
    .I4(__154__),
    .I3(__505__),
    .I2(__25__),
    .I1(__280__),
    .I0(__1333__),
    .O(__1334__)
  );
  LUT5 #(
    .INIT(32'hfffeffff)
  ) __2706__ (
    .I4(g48),
    .I3(g41),
    .I2(g30),
    .I1(g31),
    .I0(__675__),
    .O(__1335__)
  );
  LUT4 #(
    .INIT(16'h88f0)
  ) __2707__ (
    .I3(__679__),
    .I2(__162__),
    .I1(g109),
    .I0(__410__),
    .O(__1336__)
  );
  LUT6 #(
    .INIT(64'hff00bf80aaaaaaaa)
  ) __2708__ (
    .I5(g109),
    .I4(__15__),
    .I3(__197__),
    .I2(g18),
    .I1(__212__),
    .I0(__350__),
    .O(__1337__)
  );
  LUT6 #(
    .INIT(64'hff00bf80aaaaaaaa)
  ) __2709__ (
    .I5(g109),
    .I4(__15__),
    .I3(__100__),
    .I2(g18),
    .I1(__212__),
    .I0(__259__),
    .O(__1338__)
  );
  LUT6 #(
    .INIT(64'hff00bf80aaaaaaaa)
  ) __2710__ (
    .I5(g109),
    .I4(__15__),
    .I3(__444__),
    .I2(g18),
    .I1(__212__),
    .I0(__128__),
    .O(__1339__)
  );
  LUT5 #(
    .INIT(32'haaaa0a08)
  ) __2711__ (
    .I4(__37__),
    .I3(__32__),
    .I2(__345__),
    .I1(__12__),
    .I0(__368__),
    .O(__1340__)
  );
  LUT6 #(
    .INIT(64'h0caa0c0c0c0c0c0c)
  ) __2712__ (
    .I5(__56__),
    .I4(__512__),
    .I3(__295__),
    .I2(__511__),
    .I1(__457__),
    .I0(__45__),
    .O(__1341__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __2713__ (
    .I1(g109),
    .I0(__175__),
    .O(__1342__)
  );
  LUT6 #(
    .INIT(64'hff00bf80aaaaaaaa)
  ) __2714__ (
    .I5(g109),
    .I4(__15__),
    .I3(__193__),
    .I2(g18),
    .I1(__212__),
    .I0(__48__),
    .O(__1343__)
  );
  LUT6 #(
    .INIT(64'he4e464e400000000)
  ) __2715__ (
    .I5(g18),
    .I4(__478__),
    .I3(__345__),
    .I2(__32__),
    .I1(__37__),
    .I0(__733__),
    .O(__1344__)
  );
  LUT4 #(
    .INIT(16'h7800)
  ) __2716__ (
    .I3(__702__),
    .I2(__469__),
    .I1(__701__),
    .I0(__336__),
    .O(__1345__)
  );
  LUT4 #(
    .INIT(16'hf800)
  ) __2717__ (
    .I3(g109),
    .I2(__15__),
    .I1(g18),
    .I0(__212__),
    .O(__1346__)
  );
  LUT4 #(
    .INIT(16'h88f0)
  ) __2718__ (
    .I3(__679__),
    .I2(__102__),
    .I1(g109),
    .I0(__341__),
    .O(__1347__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __2719__ (
    .I2(g18),
    .I1(__24__),
    .I0(__117__),
    .O(__1348__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __2720__ (
    .I1(g109),
    .I0(__24__),
    .O(__1349__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __2721__ (
    .I2(g109),
    .I1(__356__),
    .I0(__1326__),
    .O(__1350__)
  );
  LUT5 #(
    .INIT(32'h53ac0000)
  ) __2722__ (
    .I4(g109),
    .I3(__220__),
    .I2(g18),
    .I1(__348__),
    .I0(__494__),
    .O(__1351__)
  );
  LUT4 #(
    .INIT(16'hbf80)
  ) __2723__ (
    .I3(__409__),
    .I2(__38__),
    .I1(__150__),
    .I0(__144__),
    .O(__1352__)
  );
  LUT6 #(
    .INIT(64'h000000003f5f0000)
  ) __2724__ (
    .I5(__438__),
    .I4(g750),
    .I3(__679__),
    .I2(__1286__),
    .I1(__340__),
    .I0(__1220__),
    .O(__1353__)
  );
  LUT3 #(
    .INIT(8'hb0)
  ) __2725__ (
    .I2(__358__),
    .I1(g750),
    .I0(__438__),
    .O(__1354__)
  );
  LUT6 #(
    .INIT(64'hffffffffa88a8aa8)
  ) __2726__ (
    .I5(__1354__),
    .I4(__781__),
    .I3(__1225__),
    .I2(__1224__),
    .I1(__1286__),
    .I0(__1353__),
    .O(__1355__)
  );
  LUT6 #(
    .INIT(64'hff8000ff00000000)
  ) __2727__ (
    .I5(__1178__),
    .I4(__297__),
    .I3(__679__),
    .I2(__468__),
    .I1(__61__),
    .I0(__156__),
    .O(__1356__)
  );
  LUT6 #(
    .INIT(64'hfffffffffffdffff)
  ) __2728__ (
    .I5(g48),
    .I4(g42),
    .I3(g44),
    .I2(g45),
    .I1(g43),
    .I0(__538__),
    .O(__1357__)
  );
  LUT3 #(
    .INIT(8'hb0)
  ) __2729__ (
    .I2(__184__),
    .I1(g750),
    .I0(__438__),
    .O(__1358__)
  );
  LUT6 #(
    .INIT(64'h0f030003aaaaaaaa)
  ) __2730__ (
    .I5(__747__),
    .I4(__602__),
    .I3(__73__),
    .I2(__211__),
    .I1(__1003__),
    .I0(__58__),
    .O(__1359__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __2731__ (
    .I1(g109),
    .I0(__31__),
    .O(__1360__)
  );
  LUT4 #(
    .INIT(16'h88f0)
  ) __2732__ (
    .I3(__679__),
    .I2(__420__),
    .I1(g109),
    .I0(__136__),
    .O(__1361__)
  );
  LUT4 #(
    .INIT(16'hccca)
  ) __2733__ (
    .I3(__11__),
    .I2(g1696),
    .I1(__251__),
    .I0(__40__),
    .O(__1362__)
  );
  LUT5 #(
    .INIT(32'h69960000)
  ) __2734__ (
    .I4(g109),
    .I3(__322__),
    .I2(__107__),
    .I1(__390__),
    .I0(__79__),
    .O(__1363__)
  );
  LUT4 #(
    .INIT(16'hccca)
  ) __2735__ (
    .I3(__11__),
    .I2(g1696),
    .I1(__23__),
    .I0(__134__),
    .O(__1364__)
  );
  LUT6 #(
    .INIT(64'hefffffffffffffff)
  ) __2736__ (
    .I5(g48),
    .I4(__649__),
    .I3(__647__),
    .I2(__642__),
    .I1(__938__),
    .I0(__639__),
    .O(__1365__)
  );
  LUT4 #(
    .INIT(16'hbf80)
  ) __2737__ (
    .I3(__370__),
    .I2(__393__),
    .I1(__701__),
    .I0(__505__),
    .O(__1366__)
  );
  LUT4 #(
    .INIT(16'hccca)
  ) __2738__ (
    .I3(__11__),
    .I2(g1696),
    .I1(__314__),
    .I0(__9__),
    .O(__1367__)
  );
  LUT3 #(
    .INIT(8'h40)
  ) __2739__ (
    .I2(g109),
    .I1(__279__),
    .I0(__183__),
    .O(__1368__)
  );
  LUT2 #(
    .INIT(4'he)
  ) __2740__ (
    .I1(__343__),
    .I0(g82),
    .O(__1369__)
  );
  LUT6 #(
    .INIT(64'hbfffc00000000000)
  ) __2741__ (
    .I5(__1201__),
    .I4(__201__),
    .I3(__98__),
    .I2(__14__),
    .I1(__508__),
    .I0(__411__),
    .O(__1370__)
  );
  assign g7744 = g27;
  assign g6926 = __1258__;
  assign g8562 = __1258__;
  assign g6282 = g102;
  assign g4888 = g1960;
  assign g6264 = g82;
  assign g4193 = g892;
  assign g6284 = g104;
  assign g2601 = __303__;
  assign g2610 = __303__;
  assign g2602 = __331__;
  assign g2607 = __331__;
  assign g4194 = g895;
  assign g6280 = g100;
  assign g8982 = __3__;
  assign g4176 = __456__;
  assign g11163 = __1018__;
  assign g2604 = __233__;
  assign g2609 = __233__;
  assign g4215 = g1191;
  assign g10465 = __1365__;
  assign g4198 = g904;
  assign g4201 = g913;
  assign g10459 = __939__;
  assign g8328 = __841__;
  assign g10461 = __965__;
  assign g8984 = __343__;
  assign g4211 = g1179;
  assign g6920 = __794__;
  assign g8561 = __794__;
  assign g6270 = g88;
  assign g8979 = __254__;
  assign g10457 = __1321__;
  assign g4210 = g1176;
  assign g8313 = __1259__;
  assign g4214 = g1188;
  assign g6279 = g99;
  assign g4887 = g1961;
  assign g6257 = g42;
  assign g8323 = __862__;
  assign g8318 = __783__;
  assign g4180 = __378__;
  assign g4192 = g889;
  assign g8349 = __1308__;
  assign g8335 = __764__;
  assign g4195 = g898;
  assign g4202 = g916;
  assign g4207 = g1200;
  assign g3069 = __106__;
  assign g6259 = g44;
  assign g8977 = __313__;
  assign g4203 = g919;
  assign g6281 = g101;
  assign g6254 = g30;
  assign g6258 = g43;
  assign g4178 = __445__;
  assign g6268 = g86;
  assign g4191 = g886;
  assign g4177 = __405__;
  assign g4205 = g1170;
  assign g6267 = g85;
  assign g10377 = __1335__;
  assign g2648 = __52__;
  assign g6942 = __1251__;
  assign g8564 = __1251__;
  assign g2355 = g18;
  assign g4171 = __985__;
  assign g6932 = __1144__;
  assign g8563 = __1144__;
  assign g10463 = __860__;
  assign g4208 = g1203;
  assign g8340 = __1369__;
  assign g6260 = g45;
  assign g6277 = g95;
  assign g6255 = g31;
  assign g11489 = 1'b0;
  assign g4172 = __438__;
  assign g3007 = __338__;
  assign g10455 = __1296__;
  assign g4173 = __214__;
  assign g5816 = __1__;
  assign g8271 = __1__;
  assign g6275 = g93;
  assign g6265 = g83;
  assign g4209 = g1173;
  assign g6283 = g103;
  assign g6949 = __870__;
  assign g8565 = __870__;
  assign g8316 = __1110__;
  assign g6278 = g96;
  assign g8352 = __933__;
  assign g9451 = __938__;
  assign g9961 = __938__;
  assign g4216 = g1194;
  assign g6276 = g94;
  assign g6263 = g48;
  assign g8985 = __349__;
  assign g11206 = __1301__;
  assign g2986 = __489__;
  assign g6285 = g28;
  assign g6842 = __1215__;
  assign g4179 = __497__;
  assign g4204 = g922;
  assign g10801 = __777__;
  assign g8986 = __184__;
  assign g6273 = g91;
  assign g8347 = __1217__;
  assign g6262 = g47;
  assign g5101 = g872;
  assign g8061 = g872;
  assign g4212 = g1182;
  assign g10379 = __1208__;
  assign g5659 = __895__;
  assign g6253 = g29;
  assign g4206 = g1197;
  assign g6271 = g89;
  assign g5105 = g873;
  assign g8062 = g873;
  assign g8331 = __1032__;
  assign g4196 = g925;
  assign g6266 = g84;
  assign g6272 = g90;
  assign g6955 = __514__;
  assign g8566 = __514__;
  assign g5658 = __1023__;
  assign g6261 = g46;
  assign g4181 = __42__;
  assign g4213 = g1185;
  assign g8980 = __41__;
  assign g4200 = g910;
  assign g3327 = __2__;
  assign g1957 = __196__;
  assign g4174 = __453__;
  assign g6274 = g92;
  assign g8978 = __228__;
  assign g8981 = __30__;
  assign g2603 = __158__;
  assign g2608 = __158__;
  assign g8976 = __351__;
  assign g2606 = __153__;
  assign g2612 = __153__;
  assign g2605 = __180__;
  assign g2611 = __180__;
  assign g6269 = g87;
  assign g10628 = __1056__;
  assign g4175 = __237__;
  assign g6256 = g41;
  assign g8983 = __353__;
  assign g4197 = g901;
  assign g4199 = g907;
endmodule
