module prom2 (
    x0,
    x1,
    x2,
    x3,
    x4,
    x5,
    x6,
    x7,
    x8,
    y0,
    y1,
    y2,
    y3,
    y4,
    y5,
    y6,
    y7,
    y8,
    y9,
    y10,
    y11,
    y12,
    y13,
    y14,
    y15,
    y16,
    y17,
    y18,
    y19,
    y20
);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 ;
  wire n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 ;
  assign n10 = x7 & ~x8;
  assign n11 = ~x5 & n10;
  assign n12 = ~x3 & n11;
  assign n13 = (x2 & ~x4) | (x2 & n12) | (~x4 & n12);
  assign n14 = ~x2 & n13;
  assign n15 = x1 | x2;
  assign n24 = x3 | n15;
  assign n25 = x0 & n24;
  assign n26 = x0 | n24;
  assign n27 = ~n25 & n26;
  assign n28 = x7 | x8;
  assign n29 = (~x7 & n10) | (~x7 & n28) | (n10 & n28);
  assign n16 = ~x4 & x5;
  assign n17 = ~x3 & n16;
  assign n18 = ~x0 & n17;
  assign n19 = ~n15 & n18;
  assign n20 = ~x3 & x4;
  assign n21 = ~x2 & n20;
  assign n22 = ~x0 & n21;
  assign n23 = ~x1 & n22;
  assign n30 = (n19 & n23) | (n19 & n29) | (n23 & n29);
  assign n31 = ~n27 & n30;
  assign n32 = (n27 & n29) | (n27 & n31) | (n29 & n31);
  assign n33 = (x0 & x1) | (x0 & ~n32) | (x1 & ~n32);
  assign n34 = n14 & n33;
  assign n35 = (n14 & n32) | (n14 & ~n34) | (n32 & ~n34);
  assign n42 = x2 & x3;
  assign n53 = ~x3 & x5;
  assign n54 = x5 | x8;
  assign n55 = x2 & n54;
  assign n56 = (n42 & n53) | (n42 & ~n55) | (n53 & ~n55);
  assign n57 = x1 | x7;
  assign n58 = (x4 & n56) | (x4 & n57) | (n56 & n57);
  assign n59 = n56 & ~n58;
  assign n65 = (x2 & ~x5) | (x2 & x7) | (~x5 & x7);
  assign n66 = (~x4 & x7) | (~x4 & n65) | (x7 & n65);
  assign n67 = x7 & ~n66;
  assign n68 = n66 | n67;
  assign n69 = (~x7 & n67) | (~x7 & n68) | (n67 & n68);
  assign n70 = ~x6 & x8;
  assign n71 = (x1 & ~n69) | (x1 & n70) | (~n69 & n70);
  assign n72 = n69 & n71;
  assign n37 = ~x5 & x6;
  assign n73 = x2 | x4;
  assign n74 = n37 & ~n73;
  assign n75 = (x1 & ~n28) | (x1 & n74) | (~n28 & n74);
  assign n76 = ~x1 & n75;
  assign n79 = ~x1 & x2;
  assign n77 = x6 | n28;
  assign n78 = x5 & ~n77;
  assign n80 = x3 & ~x4;
  assign n81 = n78 & n80;
  assign n82 = n79 & n81;
  assign n83 = (~n72 & n76) | (~n72 & n82) | (n76 & n82);
  assign n84 = x3 & ~n82;
  assign n85 = (n72 & n83) | (n72 & ~n84) | (n83 & ~n84);
  assign n45 = x2 | x3;
  assign n61 = x4 & ~x5;
  assign n60 = x7 & x8;
  assign n62 = x1 & n60;
  assign n63 = (n45 & n61) | (n45 & n62) | (n61 & n62);
  assign n64 = ~n45 & n63;
  assign n94 = (x1 & x2) | (x1 & ~x7) | (x2 & ~x7);
  assign n95 = x7 | n94;
  assign n96 = ~x1 & x3;
  assign n97 = (~x2 & n94) | (~x2 & n96) | (n94 & n96);
  assign n98 = (~x1 & n95) | (~x1 & n97) | (n95 & n97);
  assign n99 = x8 & n98;
  assign n91 = (x2 & x3) | (x2 & ~x7) | (x3 & ~x7);
  assign n92 = (x2 & x3) | (x2 & x8) | (x3 & x8);
  assign n93 = n91 & ~n92;
  assign n100 = n93 | n99;
  assign n101 = (~x1 & n99) | (~x1 & n100) | (n99 & n100);
  assign n86 = x4 & ~x7;
  assign n87 = x1 & x7;
  assign n88 = ~x4 & x8;
  assign n89 = x1 & ~n88;
  assign n90 = (n86 & n87) | (n86 & ~n89) | (n87 & ~n89);
  assign n102 = (~x2 & n90) | (~x2 & n101) | (n90 & n101);
  assign n103 = x3 | n102;
  assign n104 = (~x3 & n101) | (~x3 & n103) | (n101 & n103);
  assign n105 = n64 | n104;
  assign n106 = (~n59 & n85) | (~n59 & n105) | (n85 & n105);
  assign n107 = n59 | n106;
  assign n108 = ~x0 & n107;
  assign n36 = x3 | x4;
  assign n38 = ~n36 & n37;
  assign n41 = x2 & n20;
  assign n44 = x0 & ~x1;
  assign n46 = n44 & ~n45;
  assign n47 = (~n41 & n42) | (~n41 & n46) | (n42 & n46);
  assign n43 = ~x0 & x1;
  assign n48 = n43 | n46;
  assign n49 = (n41 & n47) | (n41 & n48) | (n47 & n48);
  assign n50 = (~n17 & n38) | (~n17 & n49) | (n38 & n49);
  assign n39 = x1 & x2;
  assign n40 = ~x0 & n39;
  assign n51 = n40 | n49;
  assign n52 = (n17 & n50) | (n17 & n51) | (n50 & n51);
  assign n109 = n52 | n108;
  assign n110 = (n29 & n108) | (n29 & n109) | (n108 & n109);
  assign n111 = (x4 & x5) | (x4 & ~x6) | (x5 & ~x6);
  assign n112 = (~x3 & x6) | (~x3 & n111) | (x6 & n111);
  assign n113 = (x3 & ~x4) | (x3 & n111) | (~x4 & n111);
  assign n114 = n112 | n113;
  assign n115 = x2 & ~n114;
  assign n116 = (x0 & x1) | (x0 & n115) | (x1 & n115);
  assign n117 = ~x0 & n116;
  assign n118 = x4 & x5;
  assign n119 = x3 & n118;
  assign n120 = x0 & ~x3;
  assign n121 = x1 & ~x3;
  assign n122 = (n43 & n120) | (n43 & ~n121) | (n120 & ~n121);
  assign n123 = (n17 & ~n20) | (n17 & n122) | (~n20 & n122);
  assign n124 = n43 | n122;
  assign n125 = (n20 & n123) | (n20 & n124) | (n123 & n124);
  assign n126 = ~x2 & n125;
  assign n127 = n40 | n126;
  assign n128 = (n119 & n126) | (n119 & n127) | (n126 & n127);
  assign n186 = x3 & ~x7;
  assign n187 = x5 & ~x7;
  assign n188 = (n53 & n186) | (n53 & ~n187) | (n186 & ~n187);
  assign n189 = x8 & n188;
  assign n190 = x2 & ~n189;
  assign n185 = x5 | n28;
  assign n191 = x3 & ~n185;
  assign n192 = x2 | n191;
  assign n193 = ~n190 & n192;
  assign n197 = (~x4 & x6) | (~x4 & n193) | (x6 & n193);
  assign n194 = x6 & n53;
  assign n195 = (x2 & n60) | (x2 & n194) | (n60 & n194);
  assign n196 = ~x2 & n195;
  assign n198 = x4 & n196;
  assign n199 = (n193 & ~n197) | (n193 & n198) | (~n197 & n198);
  assign n183 = x2 & ~n36;
  assign n184 = ~x7 & x8;
  assign n200 = (n183 & n184) | (n183 & n199) | (n184 & n199);
  assign n201 = n37 & ~n200;
  assign n202 = (n37 & n199) | (n37 & ~n201) | (n199 & ~n201);
  assign n203 = x1 & ~n202;
  assign n172 = (x3 & x6) | (x3 & x8) | (x6 & x8);
  assign n174 = (~x7 & x8) | (~x7 & n172) | (x8 & n172);
  assign n175 = x8 & ~n174;
  assign n176 = n174 | n175;
  assign n177 = (~x8 & n175) | (~x8 & n176) | (n175 & n176);
  assign n178 = x2 & ~x5;
  assign n179 = x2 & ~n178;
  assign n180 = n177 & n179;
  assign n171 = (x3 & x6) | (x3 & ~x7) | (x6 & ~x7);
  assign n173 = n171 & ~n172;
  assign n181 = (n173 & ~n178) | (n173 & n179) | (~n178 & n179);
  assign n182 = (~x5 & n180) | (~x5 & n181) | (n180 & n181);
  assign n204 = ~x4 & n182;
  assign n205 = x1 | n204;
  assign n206 = ~n203 & n205;
  assign n130 = (~x1 & x5) | (~x1 & x7) | (x5 & x7);
  assign n131 = (x2 & x5) | (x2 & n130) | (x5 & n130);
  assign n132 = (x1 & ~x2) | (x1 & n131) | (~x2 & n131);
  assign n133 = ~x7 & n132;
  assign n134 = (~x5 & n131) | (~x5 & n133) | (n131 & n133);
  assign n135 = x4 | n134;
  assign n129 = ~x5 & x7;
  assign n136 = n39 & n129;
  assign n137 = x4 & ~n136;
  assign n138 = n135 & ~n137;
  assign n142 = (x3 & ~x8) | (x3 & n138) | (~x8 & n138);
  assign n139 = x5 & ~n28;
  assign n140 = (x1 & ~n73) | (x1 & n139) | (~n73 & n139);
  assign n141 = ~x1 & n140;
  assign n143 = ~x3 & n141;
  assign n144 = (n138 & ~n142) | (n138 & n143) | (~n142 & n143);
  assign n155 = (x1 & x4) | (x1 & ~x8) | (x4 & ~x8);
  assign n156 = (x2 & x8) | (x2 & n155) | (x8 & n155);
  assign n157 = (x1 & x4) | (x1 & n156) | (x4 & n156);
  assign n158 = n155 & ~n157;
  assign n159 = (n156 & ~n157) | (n156 & n158) | (~n157 & n158);
  assign n160 = x3 | n159;
  assign n153 = x4 & x8;
  assign n154 = (x2 & x4) | (x2 & n153) | (x4 & n153);
  assign n161 = ~x1 & n154;
  assign n162 = x3 & ~n161;
  assign n163 = n160 & ~n162;
  assign n164 = x3 & x4;
  assign n150 = (x2 & ~x8) | (x2 & n15) | (~x8 & n15);
  assign n151 = (x2 & x8) | (x2 & ~n15) | (x8 & ~n15);
  assign n152 = (~x2 & n150) | (~x2 & n151) | (n150 & n151);
  assign n165 = (x3 & x4) | (x3 & n152) | (x4 & n152);
  assign n166 = (n163 & ~n164) | (n163 & n165) | (~n164 & n165);
  assign n167 = x7 | n166;
  assign n145 = (x1 & ~x2) | (x1 & x3) | (~x2 & x3);
  assign n146 = x1 & ~n145;
  assign n147 = x2 & x4;
  assign n148 = (~x3 & n145) | (~x3 & n147) | (n145 & n147);
  assign n149 = (x2 & ~n146) | (x2 & n148) | (~n146 & n148);
  assign n168 = x8 & ~n149;
  assign n169 = x7 & ~n168;
  assign n170 = n167 & ~n169;
  assign n207 = (~x0 & n144) | (~x0 & n170) | (n144 & n170);
  assign n208 = ~n206 & n207;
  assign n209 = (~x0 & n206) | (~x0 & n208) | (n206 & n208);
  assign n210 = (~n117 & n128) | (~n117 & n209) | (n128 & n209);
  assign n211 = n29 | n209;
  assign n212 = (n117 & n210) | (n117 & n211) | (n210 & n211);
  assign n233 = (x3 & x5) | (x3 & ~x7) | (x5 & ~x7);
  assign n234 = x5 & ~n233;
  assign n235 = (~x7 & x8) | (~x7 & n234) | (x8 & n234);
  assign n236 = (~n233 & n234) | (~n233 & n235) | (n234 & n235);
  assign n242 = x2 & n236;
  assign n237 = (x3 & ~x7) | (x3 & x8) | (~x7 & x8);
  assign n238 = (~x5 & x8) | (~x5 & n237) | (x8 & n237);
  assign n239 = x8 & ~n238;
  assign n240 = n238 | n239;
  assign n241 = (~x8 & n239) | (~x8 & n240) | (n239 & n240);
  assign n243 = x2 | n241;
  assign n244 = (~x2 & n242) | (~x2 & n243) | (n242 & n243);
  assign n245 = x1 & ~n244;
  assign n231 = x5 & n10;
  assign n232 = x2 & ~x3;
  assign n246 = n231 & n232;
  assign n247 = x1 | n246;
  assign n248 = ~n245 & n247;
  assign n249 = x4 & ~n248;
  assign n225 = (x3 & x5) | (x3 & x7) | (x5 & x7);
  assign n226 = (x3 & x8) | (x3 & ~n225) | (x8 & ~n225);
  assign n227 = (~x7 & x8) | (~x7 & n225) | (x8 & n225);
  assign n228 = ~n226 & n227;
  assign n229 = x2 & ~n228;
  assign n230 = n192 & ~n229;
  assign n250 = ~x1 & n230;
  assign n251 = x4 | n250;
  assign n252 = ~n249 & n251;
  assign n253 = x6 & ~n252;
  assign n214 = x4 | x7;
  assign n215 = (~x4 & n86) | (~x4 & n214) | (n86 & n214);
  assign n216 = x8 | n215;
  assign n217 = x5 | n216;
  assign n218 = x2 & n217;
  assign n213 = x5 & n60;
  assign n219 = x4 & n213;
  assign n220 = x2 | n219;
  assign n221 = ~n218 & n220;
  assign n222 = x3 & n221;
  assign n223 = n11 | n222;
  assign n224 = (n183 & n222) | (n183 & n223) | (n222 & n223);
  assign n254 = x1 & n224;
  assign n255 = x6 | n254;
  assign n256 = ~n253 & n255;
  assign n327 = x0 & n256;
  assign n257 = x6 & n10;
  assign n258 = n16 & n46;
  assign n259 = n257 & n258;
  assign n260 = x2 & n80;
  assign n261 = x0 & x1;
  assign n262 = x1 & ~n261;
  assign n263 = n260 & n262;
  assign n264 = (n21 & ~n261) | (n21 & n262) | (~n261 & n262);
  assign n265 = (x0 & n263) | (x0 & n264) | (n263 & n264);
  assign n324 = ~n29 & n265;
  assign n281 = (x3 & ~x5) | (x3 & x8) | (~x5 & x8);
  assign n282 = n237 & ~n281;
  assign n283 = (x3 & x7) | (x3 & ~x8) | (x7 & ~x8);
  assign n284 = (x4 & ~x8) | (x4 & n283) | (~x8 & n283);
  assign n285 = x8 & n284;
  assign n286 = n284 & ~n285;
  assign n287 = (x8 & ~n285) | (x8 & n286) | (~n285 & n286);
  assign n290 = (x2 & ~x5) | (x2 & n287) | (~x5 & n287);
  assign n288 = x4 & n10;
  assign n289 = ~n45 & n288;
  assign n291 = ~x5 & n289;
  assign n292 = (~n287 & n290) | (~n287 & n291) | (n290 & n291);
  assign n293 = (x2 & x4) | (x2 & ~n292) | (x4 & ~n292);
  assign n294 = n282 & n293;
  assign n295 = (n282 & n292) | (n282 & ~n294) | (n292 & ~n294);
  assign n296 = (~x0 & x1) | (~x0 & n295) | (x1 & n295);
  assign n271 = x5 & n184;
  assign n272 = ~x2 & x4;
  assign n273 = x4 & ~n272;
  assign n274 = n271 & n273;
  assign n275 = (n11 & ~n272) | (n11 & n273) | (~n272 & n273);
  assign n276 = (~x2 & n274) | (~x2 & n275) | (n274 & n275);
  assign n277 = x3 | n276;
  assign n266 = (x4 & x7) | (x4 & x8) | (x7 & x8);
  assign n267 = (x5 & ~x8) | (x5 & n266) | (~x8 & n266);
  assign n268 = (x4 & x7) | (x4 & n267) | (x7 & n267);
  assign n269 = ~n266 & n268;
  assign n270 = (~n267 & n268) | (~n267 & n269) | (n268 & n269);
  assign n278 = ~x2 & n270;
  assign n279 = x3 & ~n278;
  assign n280 = n277 & ~n279;
  assign n297 = (x0 & x1) | (x0 & ~n280) | (x1 & ~n280);
  assign n298 = n296 & ~n297;
  assign n303 = (x3 & x8) | (x3 & n214) | (x8 & n214);
  assign n304 = x7 & ~n303;
  assign n305 = (~x4 & n214) | (~x4 & n303) | (n214 & n303);
  assign n306 = (~x7 & n304) | (~x7 & n305) | (n304 & n305);
  assign n307 = (~x1 & x2) | (~x1 & n306) | (x2 & n306);
  assign n299 = ~x3 & x8;
  assign n300 = (~x4 & x7) | (~x4 & n299) | (x7 & n299);
  assign n301 = (x4 & ~x8) | (x4 & n299) | (~x8 & n299);
  assign n302 = (x3 & n300) | (x3 & n301) | (n300 & n301);
  assign n308 = (x1 & x2) | (x1 & ~n302) | (x2 & ~n302);
  assign n309 = n307 & ~n308;
  assign n311 = x2 | x8;
  assign n312 = (x4 & ~x7) | (x4 & n311) | (~x7 & n311);
  assign n313 = (x2 & x4) | (x2 & ~n311) | (x4 & ~n311);
  assign n314 = (x8 & ~n312) | (x8 & n313) | (~n312 & n313);
  assign n315 = (x1 & ~x3) | (x1 & n314) | (~x3 & n314);
  assign n310 = (~x2 & n28) | (~x2 & n73) | (n28 & n73);
  assign n316 = (x1 & x3) | (x1 & ~n310) | (x3 & ~n310);
  assign n317 = n315 & n316;
  assign n318 = x0 & ~n15;
  assign n319 = ~n36 & n318;
  assign n320 = n184 & n319;
  assign n321 = (~n309 & n317) | (~n309 & n320) | (n317 & n320);
  assign n322 = x0 & ~n320;
  assign n323 = (n309 & n321) | (n309 & ~n322) | (n321 & ~n322);
  assign n325 = n298 | n323;
  assign n326 = (n265 & ~n324) | (n265 & n325) | (~n324 & n325);
  assign n328 = n259 | n326;
  assign n329 = (n256 & ~n327) | (n256 & n328) | (~n327 & n328);
  assign n377 = x4 & ~x6;
  assign n354 = ~x5 & n60;
  assign n355 = (~x3 & x5) | (~x3 & x8) | (x5 & x8);
  assign n356 = (x4 & ~x8) | (x4 & n355) | (~x8 & n355);
  assign n357 = (x4 & x5) | (x4 & ~n355) | (x5 & ~n355);
  assign n358 = n356 & ~n357;
  assign n362 = (~x1 & x7) | (~x1 & n358) | (x7 & n358);
  assign n359 = x4 & n96;
  assign n360 = (x5 & x8) | (x5 & n359) | (x8 & n359);
  assign n361 = ~x8 & n360;
  assign n363 = ~x7 & n361;
  assign n364 = (n358 & ~n362) | (n358 & n363) | (~n362 & n363);
  assign n365 = (~x1 & n80) | (~x1 & n364) | (n80 & n364);
  assign n366 = n354 & ~n365;
  assign n367 = (n354 & n364) | (n354 & ~n366) | (n364 & ~n366);
  assign n368 = x2 & ~n367;
  assign n350 = (x3 & x4) | (x3 & x7) | (x4 & x7);
  assign n351 = (x3 & x4) | (x3 & ~x8) | (x4 & ~x8);
  assign n352 = n350 & ~n351;
  assign n353 = x5 & n352;
  assign n369 = ~x1 & n353;
  assign n370 = x2 | n369;
  assign n371 = ~n368 & n370;
  assign n372 = (~x0 & x6) | (~x0 & n371) | (x6 & n371);
  assign n338 = ~x1 & x4;
  assign n339 = x4 & ~n338;
  assign n340 = n188 & n339;
  assign n337 = x5 | x7;
  assign n341 = (n337 & n338) | (n337 & ~n339) | (n338 & ~n339);
  assign n342 = (x1 & ~n340) | (x1 & n341) | (~n340 & n341);
  assign n343 = ~x2 & n342;
  assign n332 = (x1 & x3) | (x1 & x5) | (x3 & x5);
  assign n333 = (~x3 & x7) | (~x3 & n332) | (x7 & n332);
  assign n334 = (x1 & x5) | (x1 & n333) | (x5 & n333);
  assign n335 = n332 & ~n334;
  assign n336 = (n333 & ~n334) | (n333 & n335) | (~n334 & n335);
  assign n344 = ~x4 & n336;
  assign n345 = x2 & ~n344;
  assign n346 = n343 | n345;
  assign n347 = x8 | n346;
  assign n330 = ~x3 & n213;
  assign n331 = ~x4 & n330;
  assign n348 = ~n331 & n347;
  assign n349 = (x1 & n347) | (x1 & n348) | (n347 & n348);
  assign n373 = (x0 & x6) | (x0 & n349) | (x6 & n349);
  assign n374 = n372 & ~n373;
  assign n398 = x3 | x5;
  assign n399 = x4 | n398;
  assign n400 = x0 & x2;
  assign n401 = x0 & ~n400;
  assign n402 = ~n399 & n401;
  assign n403 = (n119 & ~n400) | (n119 & n401) | (~n400 & n401);
  assign n404 = (x2 & n402) | (x2 & n403) | (n402 & n403);
  assign n405 = x1 | n404;
  assign n394 = (x2 & x4) | (x2 & ~x5) | (x4 & ~x5);
  assign n395 = x5 | n394;
  assign n396 = (x2 & x3) | (x2 & ~n395) | (x3 & ~n395);
  assign n397 = (n394 & n395) | (n394 & ~n396) | (n395 & ~n396);
  assign n406 = x0 | n397;
  assign n407 = x1 & n406;
  assign n408 = n405 & ~n407;
  assign n460 = ~x7 & n408;
  assign n409 = n40 & ~n337;
  assign n410 = ~n36 & n409;
  assign n437 = x4 & x7;
  assign n438 = (x4 & x8) | (x4 & ~n272) | (x8 & ~n272);
  assign n439 = (x7 & ~x8) | (x7 & n272) | (~x8 & n272);
  assign n440 = (~n437 & n438) | (~n437 & n439) | (n438 & n439);
  assign n441 = x5 & n440;
  assign n434 = (~x2 & x7) | (~x2 & x8) | (x7 & x8);
  assign n435 = ~x7 & n434;
  assign n436 = (x2 & n434) | (x2 & n435) | (n434 & n435);
  assign n442 = x4 & n436;
  assign n443 = x5 | n442;
  assign n444 = ~n441 & n443;
  assign n445 = (n16 & n86) | (n16 & ~n187) | (n86 & ~n187);
  assign n446 = (x2 & x8) | (x2 & n445) | (x8 & n445);
  assign n447 = (x0 & ~x8) | (x0 & n446) | (~x8 & n446);
  assign n448 = (x0 & x2) | (x0 & ~n446) | (x2 & ~n446);
  assign n449 = n447 & ~n448;
  assign n450 = x0 & ~n449;
  assign n451 = (n444 & n449) | (n444 & ~n450) | (n449 & ~n450);
  assign n452 = x3 | n451;
  assign n428 = x8 & n73;
  assign n429 = (n60 & n86) | (n60 & ~n428) | (n86 & ~n428);
  assign n430 = x5 | n429;
  assign n431 = n28 | n73;
  assign n432 = x5 & n431;
  assign n433 = n430 & ~n432;
  assign n453 = ~x0 & n433;
  assign n454 = x3 & ~n453;
  assign n455 = n452 & ~n454;
  assign n456 = x1 | n455;
  assign n425 = n183 & ~n271;
  assign n411 = (~x2 & x4) | (~x2 & x5) | (x4 & x5);
  assign n412 = (x2 & ~x7) | (x2 & n411) | (~x7 & n411);
  assign n413 = (x4 & x5) | (x4 & n412) | (x5 & n412);
  assign n414 = ~n411 & n413;
  assign n415 = (~n412 & n413) | (~n412 & n414) | (n413 & n414);
  assign n418 = (~x3 & x8) | (~x3 & n415) | (x8 & n415);
  assign n416 = x4 & ~n45;
  assign n417 = ~n337 & n416;
  assign n419 = ~x8 & n417;
  assign n420 = (n415 & ~n418) | (n415 & n419) | (~n418 & n419);
  assign n421 = x2 & ~n147;
  assign n422 = n354 & n421;
  assign n423 = (n139 & ~n147) | (n139 & n421) | (~n147 & n421);
  assign n424 = (x4 & n422) | (x4 & n423) | (n422 & n423);
  assign n426 = n420 | n424;
  assign n427 = (n183 & ~n425) | (n183 & n426) | (~n425 & n426);
  assign n457 = ~x0 & n427;
  assign n458 = x1 & ~n457;
  assign n459 = n456 & ~n458;
  assign n461 = n410 | n459;
  assign n462 = (n408 & ~n460) | (n408 & n461) | (~n460 & n461);
  assign n378 = x4 | x6;
  assign n379 = (~x4 & n377) | (~x4 & n378) | (n377 & n378);
  assign n380 = ~x2 & x8;
  assign n381 = (x3 & n379) | (x3 & ~n380) | (n379 & ~n380);
  assign n382 = n379 & ~n381;
  assign n383 = x1 | n382;
  assign n375 = x6 | x8;
  assign n376 = x4 & ~n375;
  assign n384 = n42 & n376;
  assign n385 = x1 & ~n384;
  assign n386 = n383 & ~n385;
  assign n390 = (~x5 & n187) | (~x5 & n337) | (n187 & n337);
  assign n391 = (x0 & n386) | (x0 & ~n390) | (n386 & ~n390);
  assign n387 = x8 & n20;
  assign n388 = (x6 & n318) | (x6 & n387) | (n318 & n387);
  assign n389 = ~x6 & n388;
  assign n392 = n389 & n390;
  assign n393 = (n386 & ~n391) | (n386 & n392) | (~n391 & n392);
  assign n463 = ~x4 & x6;
  assign n464 = n184 & n463;
  assign n465 = (x1 & x2) | (x1 & ~x8) | (x2 & ~x8);
  assign n466 = n94 & ~n465;
  assign n467 = (n10 & ~n15) | (n10 & n466) | (~n15 & n466);
  assign n468 = x3 & ~n467;
  assign n469 = (x3 & n466) | (x3 & ~n468) | (n466 & ~n468);
  assign n476 = x4 & x6;
  assign n477 = x6 & ~n476;
  assign n478 = n469 & n477;
  assign n470 = (x2 & x3) | (x2 & ~x8) | (x3 & ~x8);
  assign n471 = ~x3 & n470;
  assign n472 = (x1 & x2) | (x1 & ~n471) | (x2 & ~n471);
  assign n473 = (n470 & n471) | (n470 & ~n472) | (n471 & ~n472);
  assign n474 = x7 | n466;
  assign n475 = (n466 & n473) | (n466 & n474) | (n473 & n474);
  assign n479 = (n475 & ~n476) | (n475 & n477) | (~n476 & n477);
  assign n480 = (x4 & n478) | (x4 & n479) | (n478 & n479);
  assign n481 = ~x0 & n480;
  assign n482 = n46 | n481;
  assign n483 = (n464 & n481) | (n464 & n482) | (n481 & n482);
  assign n484 = n393 | n483;
  assign n485 = (~n374 & n462) | (~n374 & n484) | (n462 & n484);
  assign n486 = n374 | n485;
  assign n500 = (x2 & x7) | (x2 & ~x8) | (x7 & ~x8);
  assign n501 = (x5 & x7) | (x5 & x8) | (x7 & x8);
  assign n502 = ~n500 & n501;
  assign n503 = (x2 & x5) | (x2 & n29) | (x5 & n29);
  assign n504 = (x0 & ~x5) | (x0 & n503) | (~x5 & n503);
  assign n505 = (x0 & x2) | (x0 & ~n503) | (x2 & ~n503);
  assign n506 = n504 & ~n505;
  assign n507 = x0 & ~n506;
  assign n508 = (n502 & n506) | (n502 & ~n507) | (n506 & ~n507);
  assign n509 = x1 | n508;
  assign n495 = (x5 & x7) | (x5 & ~n434) | (x7 & ~n434);
  assign n496 = (~x7 & x8) | (~x7 & n495) | (x8 & n495);
  assign n497 = n434 & n496;
  assign n498 = x5 & ~n497;
  assign n499 = (n495 & n497) | (n495 & ~n498) | (n497 & ~n498);
  assign n510 = ~x0 & n499;
  assign n511 = x1 & ~n510;
  assign n512 = n509 & ~n511;
  assign n513 = x3 | n512;
  assign n488 = (x1 & x2) | (x1 & x8) | (x2 & x8);
  assign n489 = (x7 & ~x8) | (x7 & n488) | (~x8 & n488);
  assign n490 = (x1 & x2) | (x1 & n489) | (x2 & n489);
  assign n491 = n488 & ~n490;
  assign n492 = (n489 & ~n490) | (n489 & n491) | (~n490 & n491);
  assign n487 = x1 & ~x2;
  assign n493 = n487 | n492;
  assign n494 = (n213 & n492) | (n213 & n493) | (n492 & n493);
  assign n514 = ~x0 & n494;
  assign n515 = x3 & ~n514;
  assign n516 = n513 & ~n515;
  assign n517 = (x4 & ~x6) | (x4 & n516) | (~x6 & n516);
  assign n518 = (~n377 & n486) | (~n377 & n517) | (n486 & n517);
  assign n534 = (x0 & ~x4) | (x0 & x5) | (~x4 & x5);
  assign n535 = (~x3 & x5) | (~x3 & n534) | (x5 & n534);
  assign n536 = x5 & ~n535;
  assign n537 = n535 | n536;
  assign n538 = (~x5 & n536) | (~x5 & n537) | (n536 & n537);
  assign n539 = x2 | n538;
  assign n530 = (x3 & ~x4) | (x3 & x5) | (~x4 & x5);
  assign n531 = x6 | n530;
  assign n532 = (~x5 & x6) | (~x5 & n530) | (x6 & n530);
  assign n533 = (x5 & ~n531) | (x5 & n532) | (~n531 & n532);
  assign n540 = ~x0 & n533;
  assign n541 = x2 & ~n540;
  assign n542 = n539 & ~n541;
  assign n543 = x1 | n542;
  assign n521 = (~x2 & x3) | (~x2 & x5) | (x3 & x5);
  assign n522 = (x2 & ~x4) | (x2 & n521) | (~x4 & n521);
  assign n523 = (x3 & x5) | (x3 & n522) | (x5 & n522);
  assign n524 = ~n521 & n523;
  assign n525 = (~n522 & n523) | (~n522 & n524) | (n523 & n524);
  assign n526 = x6 & ~n525;
  assign n519 = x2 & ~x4;
  assign n520 = (x4 & ~n20) | (x4 & n519) | (~n20 & n519);
  assign n527 = x5 | n520;
  assign n528 = ~x6 & n527;
  assign n529 = n526 | n528;
  assign n544 = x0 | n529;
  assign n545 = x1 & n544;
  assign n546 = n543 & ~n545;
  assign n735 = n29 & n546;
  assign n551 = ~x6 & n390;
  assign n556 = x4 & ~n147;
  assign n557 = n551 & n556;
  assign n552 = ~x6 & x7;
  assign n553 = ~x5 & n552;
  assign n554 = x6 & n187;
  assign n555 = n553 | n554;
  assign n558 = (~n147 & n555) | (~n147 & n556) | (n555 & n556);
  assign n559 = (x2 & n557) | (x2 & n558) | (n557 & n558);
  assign n560 = x1 & ~n559;
  assign n547 = (x4 & x5) | (x4 & ~x7) | (x5 & ~x7);
  assign n548 = x4 & ~n547;
  assign n549 = (x5 & x6) | (x5 & n548) | (x6 & n548);
  assign n550 = (~n547 & n548) | (~n547 & n549) | (n548 & n549);
  assign n561 = ~x2 & n550;
  assign n562 = x1 | n561;
  assign n563 = ~n560 & n562;
  assign n568 = (x0 & ~x3) | (x0 & n563) | (~x3 & n563);
  assign n564 = x6 | x7;
  assign n565 = ~n45 & n61;
  assign n566 = (x1 & ~n564) | (x1 & n565) | (~n564 & n565);
  assign n567 = ~x1 & n566;
  assign n569 = ~x0 & n567;
  assign n570 = (n563 & ~n568) | (n563 & n569) | (~n568 & n569);
  assign n583 = x6 & x7;
  assign n584 = n46 & n583;
  assign n585 = n61 & n584;
  assign n572 = x6 & n184;
  assign n573 = ~x1 & x5;
  assign n574 = (n96 & n232) | (n96 & ~n573) | (n232 & ~n573);
  assign n575 = (~x2 & n232) | (~x2 & n574) | (n232 & n574);
  assign n576 = ~x4 & n575;
  assign n577 = ~x0 & n576;
  assign n578 = (~x3 & n118) | (~x3 & n577) | (n118 & n577);
  assign n579 = n318 & ~n578;
  assign n580 = (n318 & n577) | (n318 & ~n579) | (n577 & ~n579);
  assign n571 = ~x6 & n10;
  assign n581 = n571 & n580;
  assign n582 = (n572 & n580) | (n572 & n581) | (n580 & n581);
  assign n632 = x5 | x6;
  assign n633 = (x2 & x6) | (x2 & x8) | (x6 & x8);
  assign n634 = x5 & x8;
  assign n635 = (~x6 & n633) | (~x6 & n634) | (n633 & n634);
  assign n636 = (~x2 & x6) | (~x2 & x7) | (x6 & x7);
  assign n637 = x2 & n636;
  assign n638 = (x5 & x6) | (x5 & ~n637) | (x6 & ~n637);
  assign n639 = (n636 & n637) | (n636 & ~n638) | (n637 & ~n638);
  assign n644 = (x4 & ~x8) | (x4 & n639) | (~x8 & n639);
  assign n591 = x5 & x6;
  assign n640 = x6 & ~x7;
  assign n641 = (~x2 & n591) | (~x2 & n640) | (n591 & n640);
  assign n642 = (~x2 & x7) | (~x2 & n591) | (x7 & n591);
  assign n643 = (x7 & n641) | (x7 & ~n642) | (n641 & ~n642);
  assign n645 = (x4 & x8) | (x4 & ~n643) | (x8 & ~n643);
  assign n646 = n644 & ~n645;
  assign n647 = (x4 & x7) | (x4 & ~n646) | (x7 & ~n646);
  assign n648 = n635 & n647;
  assign n649 = (n635 & n646) | (n635 & ~n648) | (n646 & ~n648);
  assign n671 = (~x0 & x3) | (~x0 & n649) | (x3 & n649);
  assign n658 = (x5 & ~x7) | (x5 & x8) | (~x7 & x8);
  assign n659 = (x2 & x7) | (x2 & n658) | (x7 & n658);
  assign n660 = (x7 & x8) | (x7 & ~n659) | (x8 & ~n659);
  assign n661 = n658 & n660;
  assign n662 = (x2 & ~n659) | (x2 & n661) | (~n659 & n661);
  assign n663 = x6 | n662;
  assign n655 = x5 & ~x8;
  assign n656 = (~x5 & n54) | (~x5 & n655) | (n54 & n655);
  assign n657 = x7 & n656;
  assign n664 = x2 & n657;
  assign n665 = x6 & ~n664;
  assign n666 = n663 & ~n665;
  assign n667 = x4 | n666;
  assign n650 = (x5 & x6) | (x5 & ~x8) | (x6 & ~x8);
  assign n651 = (x2 & ~x5) | (x2 & n650) | (~x5 & n650);
  assign n652 = (x5 & x8) | (x5 & n651) | (x8 & n651);
  assign n653 = n650 & ~n652;
  assign n654 = (x2 & ~n651) | (x2 & n653) | (~n651 & n653);
  assign n668 = x7 & n654;
  assign n669 = x4 & ~n668;
  assign n670 = n667 & ~n669;
  assign n672 = (x0 & x3) | (x0 & ~n670) | (x3 & ~n670);
  assign n673 = n671 & ~n672;
  assign n624 = x2 | n36;
  assign n631 = x0 & ~n624;
  assign n674 = (n184 & n631) | (n184 & n673) | (n631 & n673);
  assign n675 = n632 | n674;
  assign n676 = (~n632 & n673) | (~n632 & n675) | (n673 & n675);
  assign n677 = x1 | n676;
  assign n594 = (x4 & ~x5) | (x4 & x6) | (~x5 & x6);
  assign n595 = (x5 & ~x7) | (x5 & n594) | (~x7 & n594);
  assign n596 = (x4 & x6) | (x4 & n595) | (x6 & n595);
  assign n597 = n594 & ~n596;
  assign n598 = (n595 & ~n596) | (n595 & n597) | (~n596 & n597);
  assign n599 = x3 & n598;
  assign n586 = (x4 & x5) | (x4 & x6) | (x5 & x6);
  assign n592 = (x4 & ~x7) | (x4 & n591) | (~x7 & n591);
  assign n593 = n586 & ~n592;
  assign n600 = x3 | n593;
  assign n601 = (~x3 & n599) | (~x3 & n600) | (n599 & n600);
  assign n602 = x8 | n601;
  assign n587 = (x6 & x7) | (x6 & ~n586) | (x7 & ~n586);
  assign n588 = (x4 & x5) | (x4 & ~n587) | (x5 & ~n587);
  assign n589 = ~n586 & n588;
  assign n590 = (n587 & n588) | (n587 & n589) | (n588 & n589);
  assign n603 = ~x3 & n590;
  assign n604 = x8 & ~n603;
  assign n605 = n602 & ~n604;
  assign n623 = x2 & n164;
  assign n625 = n11 & ~n624;
  assign n626 = n271 | n625;
  assign n627 = (n623 & n625) | (n623 & n626) | (n625 & n626);
  assign n628 = (x2 & n605) | (x2 & n627) | (n605 & n627);
  assign n609 = (~x3 & x4) | (~x3 & x6) | (x4 & x6);
  assign n610 = (x4 & x7) | (x4 & ~n609) | (x7 & ~n609);
  assign n611 = (x3 & ~x6) | (x3 & n610) | (~x6 & n610);
  assign n612 = n609 & n611;
  assign n613 = (~n610 & n611) | (~n610 & n612) | (n611 & n612);
  assign n614 = x8 | n613;
  assign n606 = (x3 & x7) | (x3 & n80) | (x7 & n80);
  assign n607 = (~x3 & x7) | (~x3 & n80) | (x7 & n80);
  assign n608 = (x3 & ~n606) | (x3 & n607) | (~n606 & n607);
  assign n615 = x6 & n608;
  assign n616 = x8 & ~n615;
  assign n617 = n614 & ~n616;
  assign n618 = x3 & ~x5;
  assign n619 = (x4 & n571) | (x4 & n618) | (n571 & n618);
  assign n620 = ~x4 & n619;
  assign n621 = x5 | n620;
  assign n622 = (n617 & n620) | (n617 & n621) | (n620 & n621);
  assign n629 = (~x2 & n622) | (~x2 & n627) | (n622 & n627);
  assign n630 = n628 | n629;
  assign n678 = ~x0 & n630;
  assign n679 = x1 & ~n678;
  assign n680 = n677 & ~n679;
  assign n681 = n582 | n680;
  assign n682 = (~n570 & n585) | (~n570 & n681) | (n585 & n681);
  assign n683 = n570 | n682;
  assign n708 = (x2 & x6) | (x2 & ~x8) | (x6 & ~x8);
  assign n709 = (~x2 & x4) | (~x2 & n708) | (x4 & n708);
  assign n710 = (~x4 & x8) | (~x4 & n708) | (x8 & n708);
  assign n711 = n709 & n710;
  assign n712 = x4 & ~x8;
  assign n713 = (x0 & x2) | (x0 & n712) | (x2 & n712);
  assign n714 = (x2 & x4) | (x2 & ~n713) | (x4 & ~n713);
  assign n715 = (x0 & ~x8) | (x0 & n714) | (~x8 & n714);
  assign n716 = ~n713 & n715;
  assign n721 = (~x5 & x6) | (~x5 & n716) | (x6 & n716);
  assign n717 = ~x5 & x8;
  assign n718 = x4 & n717;
  assign n719 = (x0 & x2) | (x0 & n718) | (x2 & n718);
  assign n720 = ~x0 & n719;
  assign n722 = ~x6 & n720;
  assign n723 = (n716 & ~n721) | (n716 & n722) | (~n721 & n722);
  assign n724 = (x0 & x5) | (x0 & ~n723) | (x5 & ~n723);
  assign n725 = n711 & n724;
  assign n726 = (n711 & n723) | (n711 & ~n725) | (n723 & ~n725);
  assign n727 = x3 | n726;
  assign n702 = (~x2 & x5) | (~x2 & x6) | (x5 & x6);
  assign n703 = (x2 & x4) | (x2 & n702) | (x4 & n702);
  assign n704 = (x5 & x6) | (x5 & n703) | (x6 & n703);
  assign n705 = n702 & ~n704;
  assign n706 = (n703 & ~n704) | (n703 & n705) | (~n704 & n705);
  assign n707 = ~x8 & n706;
  assign n728 = ~x0 & n707;
  assign n729 = x3 & ~n728;
  assign n730 = n727 & ~n729;
  assign n731 = x1 | n730;
  assign n685 = x2 & ~x8;
  assign n686 = x2 & ~n685;
  assign n687 = x4 & n686;
  assign n688 = (x6 & ~n685) | (x6 & n686) | (~n685 & n686);
  assign n689 = (~x8 & n687) | (~x8 & n688) | (n687 & n688);
  assign n695 = x3 & n689;
  assign n690 = (x2 & x4) | (x2 & x8) | (x4 & x8);
  assign n691 = (x4 & ~x6) | (x4 & n690) | (~x6 & n690);
  assign n692 = x4 & ~n691;
  assign n693 = n691 | n692;
  assign n694 = (~x4 & n692) | (~x4 & n693) | (n692 & n693);
  assign n696 = x3 | n694;
  assign n697 = (~x3 & n695) | (~x3 & n696) | (n695 & n696);
  assign n698 = x5 | n697;
  assign n684 = x6 & ~x8;
  assign n699 = n623 & n684;
  assign n700 = x5 & ~n699;
  assign n701 = n698 & ~n700;
  assign n732 = ~x0 & n701;
  assign n733 = x1 & ~n732;
  assign n734 = n731 & ~n733;
  assign n736 = n683 | n734;
  assign n737 = (n546 & ~n735) | (n546 & n736) | (~n735 & n736);
  assign n755 = x5 & x7;
  assign n756 = (~x5 & n20) | (~x5 & n755) | (n20 & n755);
  assign n757 = ~x1 & n756;
  assign n758 = ~x2 & n757;
  assign n759 = x0 & n758;
  assign n739 = (~x1 & x2) | (~x1 & x7) | (x2 & x7);
  assign n740 = ~x2 & n739;
  assign n741 = (x1 & ~x5) | (x1 & n740) | (~x5 & n740);
  assign n742 = (n739 & n740) | (n739 & n741) | (n740 & n741);
  assign n747 = (~x3 & x4) | (~x3 & n742) | (x4 & n742);
  assign n743 = (x1 & ~x2) | (x1 & x5) | (~x2 & x5);
  assign n744 = n65 & ~n743;
  assign n745 = x7 & ~n744;
  assign n746 = (n743 & n744) | (n743 & ~n745) | (n744 & ~n745);
  assign n748 = (x3 & x4) | (x3 & n746) | (x4 & n746);
  assign n749 = n747 & ~n748;
  assign n750 = (~n118 & n187) | (~n118 & n214) | (n187 & n214);
  assign n751 = (x2 & x3) | (x2 & ~n750) | (x3 & ~n750);
  assign n752 = (x1 & ~x3) | (x1 & n751) | (~x3 & n751);
  assign n753 = (x1 & x2) | (x1 & ~n751) | (x2 & ~n751);
  assign n754 = n752 & ~n753;
  assign n760 = n749 | n754;
  assign n761 = ~x0 & n760;
  assign n762 = n759 | n761;
  assign n738 = (~x6 & n375) | (~x6 & n684) | (n375 & n684);
  assign n917 = n738 & n762;
  assign n765 = x4 | x5;
  assign n766 = (x2 & x3) | (x2 & n765) | (x3 & n765);
  assign n767 = (x2 & x3) | (x2 & ~n765) | (x3 & ~n765);
  assign n768 = (x4 & x5) | (x4 & n767) | (x5 & n767);
  assign n769 = n766 & ~n768;
  assign n770 = x1 & n769;
  assign n763 = x2 | x5;
  assign n764 = (x2 & n80) | (x2 & ~n763) | (n80 & ~n763);
  assign n771 = x1 | n764;
  assign n772 = (~x1 & n770) | (~x1 & n771) | (n770 & n771);
  assign n781 = (~x0 & x7) | (~x0 & n772) | (x7 & n772);
  assign n773 = x2 | n53;
  assign n774 = (x2 & ~x4) | (x2 & n53) | (~x4 & n53);
  assign n775 = n773 & ~n774;
  assign n776 = (~x2 & n773) | (~x2 & n775) | (n773 & n775);
  assign n777 = x1 | n776;
  assign n778 = x2 & n119;
  assign n779 = x1 & ~n778;
  assign n780 = n777 & ~n779;
  assign n782 = (x0 & x7) | (x0 & ~n780) | (x7 & ~n780);
  assign n783 = n781 & ~n782;
  assign n790 = ~x4 & x7;
  assign n784 = x2 & x5;
  assign n785 = (x3 & ~n43) | (x3 & n784) | (~n43 & n784);
  assign n786 = n43 & n785;
  assign n787 = ~x3 & n44;
  assign n788 = (x2 & ~x5) | (x2 & n787) | (~x5 & n787);
  assign n789 = ~x2 & n788;
  assign n791 = n786 | n789;
  assign n792 = (~x4 & x7) | (~x4 & n791) | (x7 & n791);
  assign n793 = (n790 & n791) | (n790 & ~n792) | (n791 & ~n792);
  assign n794 = n783 | n793;
  assign n795 = (~x6 & x8) | (~x6 & n794) | (x8 & n794);
  assign n796 = (n70 & n794) | (n70 & ~n795) | (n794 & ~n795);
  assign n797 = (x2 & x3) | (x2 & x7) | (x3 & x7);
  assign n798 = (~x5 & x7) | (~x5 & n797) | (x7 & n797);
  assign n799 = x7 & ~n798;
  assign n800 = n798 | n799;
  assign n801 = (~x7 & n799) | (~x7 & n800) | (n799 & n800);
  assign n804 = (x1 & x6) | (x1 & ~n801) | (x6 & ~n801);
  assign n802 = x3 & n79;
  assign n803 = ~n337 & n802;
  assign n805 = x6 & n803;
  assign n806 = (n801 & n804) | (n801 & n805) | (n804 & n805);
  assign n807 = x3 | n632;
  assign n808 = (x1 & x2) | (x1 & ~n807) | (x2 & ~n807);
  assign n809 = ~x1 & n808;
  assign n860 = x5 & ~n564;
  assign n813 = ~x2 & x5;
  assign n861 = (~x3 & x4) | (~x3 & n813) | (x4 & n813);
  assign n862 = (x2 & x3) | (x2 & n861) | (x3 & n861);
  assign n863 = (x4 & x5) | (x4 & ~n862) | (x5 & ~n862);
  assign n864 = ~n861 & n863;
  assign n865 = x4 & n232;
  assign n866 = n129 & n865;
  assign n867 = x7 & ~n866;
  assign n868 = (n864 & n866) | (n864 & ~n867) | (n866 & ~n867);
  assign n869 = x6 & n868;
  assign n870 = n260 | n869;
  assign n871 = (n860 & n869) | (n860 & n870) | (n869 & n870);
  assign n872 = x8 & n871;
  assign n851 = x5 & ~x6;
  assign n852 = (~n16 & n463) | (~n16 & n851) | (n463 & n851);
  assign n853 = (~x2 & x7) | (~x2 & n852) | (x7 & n852);
  assign n854 = ~x7 & n853;
  assign n855 = (x2 & x3) | (x2 & n854) | (x3 & n854);
  assign n856 = (n853 & n854) | (n853 & n855) | (n854 & n855);
  assign n846 = (x2 & ~x5) | (x2 & n20) | (~x5 & n20);
  assign n847 = (x2 & x3) | (x2 & ~x5) | (x3 & ~x5);
  assign n848 = (~x3 & x4) | (~x3 & n846) | (x4 & n846);
  assign n849 = (n20 & n847) | (n20 & ~n848) | (n847 & ~n848);
  assign n850 = n846 & ~n849;
  assign n857 = (~x6 & n850) | (~x6 & n856) | (n850 & n856);
  assign n858 = x7 | n857;
  assign n859 = (~x7 & n856) | (~x7 & n858) | (n856 & n858);
  assign n873 = x8 | n859;
  assign n874 = (~x8 & n872) | (~x8 & n873) | (n872 & n873);
  assign n875 = x1 & n874;
  assign n812 = ~x2 & x3;
  assign n814 = (x2 & x7) | (x2 & n813) | (x7 & n813);
  assign n815 = (x3 & x7) | (x3 & n813) | (x7 & n813);
  assign n816 = (n812 & n814) | (n812 & ~n815) | (n814 & ~n815);
  assign n817 = ~n45 & n553;
  assign n818 = x6 | n817;
  assign n819 = (n816 & n817) | (n816 & n818) | (n817 & n818);
  assign n822 = (x4 & ~x8) | (x4 & n819) | (~x8 & n819);
  assign n820 = x2 & ~n77;
  assign n821 = n53 & n820;
  assign n823 = ~x4 & n821;
  assign n824 = (n819 & ~n822) | (n819 & n823) | (~n822 & n823);
  assign n836 = (x5 & x6) | (x5 & ~n658) | (x6 & ~n658);
  assign n837 = (x7 & ~x8) | (x7 & n836) | (~x8 & n836);
  assign n838 = n658 & n837;
  assign n839 = (~n836 & n837) | (~n836 & n838) | (n837 & n838);
  assign n840 = x2 & n839;
  assign n833 = (~x6 & x7) | (~x6 & x8) | (x7 & x8);
  assign n834 = (x5 & x6) | (x5 & ~n833) | (x6 & ~n833);
  assign n835 = (~x6 & n717) | (~x6 & n834) | (n717 & n834);
  assign n841 = x2 | n835;
  assign n842 = (~x2 & n840) | (~x2 & n841) | (n840 & n841);
  assign n843 = (~x3 & x4) | (~x3 & n842) | (x4 & n842);
  assign n825 = (x6 & ~x7) | (x6 & x8) | (~x7 & x8);
  assign n826 = (x2 & ~x8) | (x2 & n825) | (~x8 & n825);
  assign n827 = (x2 & x6) | (x2 & ~n825) | (x6 & ~n825);
  assign n828 = n826 & ~n827;
  assign n829 = x5 & ~n828;
  assign n830 = ~x2 & n60;
  assign n831 = x5 | n830;
  assign n832 = ~n829 & n831;
  assign n844 = (x3 & x4) | (x3 & n832) | (x4 & n832);
  assign n845 = n843 & n844;
  assign n876 = n824 | n845;
  assign n877 = ~x1 & n876;
  assign n878 = n875 | n877;
  assign n879 = (~n806 & n809) | (~n806 & n878) | (n809 & n878);
  assign n810 = x4 | x8;
  assign n811 = (~x4 & n712) | (~x4 & n810) | (n712 & n810);
  assign n880 = n811 | n878;
  assign n881 = (n806 & n879) | (n806 & n880) | (n879 & n880);
  assign n914 = x0 & n881;
  assign n882 = ~x6 & n60;
  assign n883 = n258 & n882;
  assign n897 = x0 & x5;
  assign n898 = (x3 & ~x6) | (x3 & n897) | (~x6 & n897);
  assign n899 = (x0 & x3) | (x0 & ~n898) | (x3 & ~n898);
  assign n900 = (x5 & ~x6) | (x5 & n899) | (~x6 & n899);
  assign n901 = ~n898 & n900;
  assign n902 = ~x7 & n901;
  assign n903 = x1 | n902;
  assign n896 = (x3 & ~n398) | (x3 & n583) | (~n398 & n583);
  assign n904 = ~x0 & n896;
  assign n905 = x1 & ~n904;
  assign n906 = n903 & ~n905;
  assign n907 = x2 | n906;
  assign n890 = (x1 & x5) | (x1 & x6) | (x5 & x6);
  assign n891 = (~x1 & x3) | (~x1 & n890) | (x3 & n890);
  assign n892 = (x5 & x6) | (x5 & n891) | (x6 & n891);
  assign n893 = ~n890 & n892;
  assign n894 = (~n891 & n892) | (~n891 & n893) | (n892 & n893);
  assign n895 = x7 & n894;
  assign n908 = ~x0 & n895;
  assign n909 = x2 & ~n908;
  assign n910 = n907 & ~n909;
  assign n911 = ~x4 & n910;
  assign n884 = (x2 & x6) | (x2 & ~x7) | (x6 & ~x7);
  assign n885 = (x2 & ~x5) | (x2 & x6) | (~x5 & x6);
  assign n886 = ~n884 & n885;
  assign n887 = x1 & x4;
  assign n888 = (x3 & ~n886) | (x3 & n887) | (~n886 & n887);
  assign n889 = n886 & n888;
  assign n912 = n889 | n911;
  assign n913 = (~x0 & n911) | (~x0 & n912) | (n911 & n912);
  assign n915 = n883 | n913;
  assign n916 = (n881 & ~n914) | (n881 & n915) | (~n914 & n915);
  assign n918 = n796 | n916;
  assign n919 = (n762 & ~n917) | (n762 & n918) | (~n917 & n918);
  assign n994 = x6 & x8;
  assign n1061 = x1 & ~x4;
  assign n1062 = x3 & n1061;
  assign n1063 = (~x1 & x2) | (~x1 & n1061) | (x2 & n1061);
  assign n1064 = (~x3 & n487) | (~x3 & n1063) | (n487 & n1063);
  assign n1065 = (x3 & ~n1062) | (x3 & n1064) | (~n1062 & n1064);
  assign n1066 = (x1 & x2) | (x1 & ~x4) | (x2 & ~x4);
  assign n1067 = (x1 & ~x5) | (x1 & n1066) | (~x5 & n1066);
  assign n1068 = x1 & ~n1067;
  assign n1069 = n1067 | n1068;
  assign n1070 = (~x1 & n1068) | (~x1 & n1069) | (n1068 & n1069);
  assign n1071 = x5 & ~n1070;
  assign n1072 = (n1065 & ~n1070) | (n1065 & n1071) | (~n1070 & n1071);
  assign n1079 = x8 & ~n1072;
  assign n1074 = (n20 & ~n178) | (n20 & n767) | (~n178 & n767);
  assign n1075 = x1 | n1074;
  assign n1073 = x3 & n16;
  assign n1076 = x2 & n1073;
  assign n1077 = x1 & ~n1076;
  assign n1078 = n1075 & ~n1077;
  assign n1080 = x8 | n1078;
  assign n1081 = (~x8 & n1079) | (~x8 & n1080) | (n1079 & n1080);
  assign n1082 = (~x0 & x6) | (~x0 & n1081) | (x6 & n1081);
  assign n1045 = (~x2 & x3) | (~x2 & x8) | (x3 & x8);
  assign n1046 = n521 & ~n1045;
  assign n1047 = (x2 & x3) | (x2 & ~n42) | (x3 & ~n42);
  assign n1048 = (x1 & ~x4) | (x1 & n1047) | (~x4 & n1047);
  assign n1049 = ~n42 & n1048;
  assign n1055 = (~x5 & x8) | (~x5 & n1049) | (x8 & n1049);
  assign n1050 = (x1 & x3) | (x1 & x4) | (x3 & x4);
  assign n1051 = (~x2 & x4) | (~x2 & n1050) | (x4 & n1050);
  assign n1052 = x4 & ~n1051;
  assign n1053 = n1051 | n1052;
  assign n1054 = (~x4 & n1052) | (~x4 & n1053) | (n1052 & n1053);
  assign n1056 = (x5 & x8) | (x5 & n1054) | (x8 & n1054);
  assign n1057 = n1055 & n1056;
  assign n1058 = (x1 & ~x4) | (x1 & n1057) | (~x4 & n1057);
  assign n1059 = n1046 & ~n1058;
  assign n1060 = (n1046 & n1057) | (n1046 & ~n1059) | (n1057 & ~n1059);
  assign n1083 = (x0 & x6) | (x0 & ~n1060) | (x6 & ~n1060);
  assign n1084 = n1082 & ~n1083;
  assign n1036 = ~x4 & n299;
  assign n1037 = (x1 & ~x4) | (x1 & x8) | (~x4 & x8);
  assign n1038 = x8 & ~n1037;
  assign n1039 = (x1 & x2) | (x1 & n1038) | (x2 & n1038);
  assign n1040 = (~n1037 & n1038) | (~n1037 & n1039) | (n1038 & n1039);
  assign n1041 = x3 & n1040;
  assign n1042 = ~x0 & n1041;
  assign n1043 = n15 & ~n1042;
  assign n1044 = (n1036 & n1042) | (n1036 & ~n1043) | (n1042 & ~n1043);
  assign n1085 = (x5 & x6) | (x5 & ~n1044) | (x6 & ~n1044);
  assign n1086 = (n632 & n1084) | (n632 & ~n1085) | (n1084 & ~n1085);
  assign n1087 = x7 & ~n1086;
  assign n1013 = (~x4 & x5) | (~x4 & x6) | (x5 & x6);
  assign n1014 = x4 & n1013;
  assign n1015 = (x3 & ~x6) | (x3 & n1014) | (~x6 & n1014);
  assign n1016 = (n1013 & n1014) | (n1013 & n1015) | (n1014 & n1015);
  assign n1029 = ~x2 & n1016;
  assign n1017 = (x4 & x5) | (x4 & ~x8) | (x5 & ~x8);
  assign n1018 = (~x5 & x6) | (~x5 & x8) | (x6 & x8);
  assign n1019 = ~x4 & n1018;
  assign n1020 = n1017 | n1019;
  assign n1024 = (x2 & x3) | (x2 & ~n1020) | (x3 & ~n1020);
  assign n1021 = x5 | n375;
  assign n1022 = x4 & ~n1021;
  assign n1023 = x2 & n1022;
  assign n1025 = ~x3 & n1023;
  assign n1026 = (n1020 & n1024) | (n1020 & ~n1025) | (n1024 & ~n1025);
  assign n1027 = ~x4 & n812;
  assign n1028 = ~n632 & n1027;
  assign n1030 = n1026 & ~n1028;
  assign n1031 = (~n1016 & n1029) | (~n1016 & n1030) | (n1029 & n1030);
  assign n1032 = x1 & ~n1031;
  assign n995 = (~x6 & n272) | (~x6 & n656) | (n272 & n656);
  assign n996 = ~n656 & n995;
  assign n997 = (n519 & n994) | (n519 & n996) | (n994 & n996);
  assign n998 = x5 & ~n997;
  assign n999 = (x5 & n996) | (x5 & ~n998) | (n996 & ~n998);
  assign n1000 = (x4 & x6) | (x4 & x8) | (x6 & x8);
  assign n1001 = x8 & n1000;
  assign n1002 = (x2 & x4) | (x2 & n1000) | (x4 & n1000);
  assign n1003 = x8 | n1002;
  assign n1004 = ~n1001 & n1003;
  assign n1005 = x3 | n1004;
  assign n1006 = x2 & n153;
  assign n1007 = x3 & ~n1006;
  assign n1008 = n1005 & ~n1007;
  assign n1009 = x5 | n1008;
  assign n1010 = ~n624 & n994;
  assign n1011 = x5 & ~n1010;
  assign n1012 = n1009 & ~n1011;
  assign n1033 = n999 | n1012;
  assign n1034 = ~x1 & n1033;
  assign n1035 = n1032 | n1034;
  assign n1088 = ~x0 & n1035;
  assign n1089 = x7 | n1088;
  assign n1090 = ~n1087 & n1089;
  assign n972 = (x0 & x4) | (x0 & x5) | (x4 & x5);
  assign n973 = (x4 & x7) | (x4 & ~n972) | (x7 & ~n972);
  assign n974 = (x0 & x5) | (x0 & ~n973) | (x5 & ~n973);
  assign n975 = ~n972 & n974;
  assign n976 = (n973 & n974) | (n973 & n975) | (n974 & n975);
  assign n983 = x1 & n976;
  assign n977 = (x0 & x4) | (x0 & n390) | (x4 & n390);
  assign n978 = (x1 & ~x4) | (x1 & n977) | (~x4 & n977);
  assign n979 = (x0 & x1) | (x0 & ~n977) | (x1 & ~n977);
  assign n980 = n978 & ~n979;
  assign n981 = ~x4 & n43;
  assign n982 = ~n337 & n981;
  assign n984 = n980 | n982;
  assign n985 = (n976 & ~n983) | (n976 & n984) | (~n983 & n984);
  assign n986 = x2 | n985;
  assign n968 = (x1 & x5) | (x1 & ~n437) | (x5 & ~n437);
  assign n969 = (x1 & ~x5) | (x1 & x7) | (~x5 & x7);
  assign n970 = x1 & ~n969;
  assign n971 = n968 & ~n970;
  assign n987 = ~x0 & n971;
  assign n988 = x2 & ~n987;
  assign n989 = n986 & ~n988;
  assign n990 = x3 | n989;
  assign n941 = x5 & n790;
  assign n963 = ~x2 & n941;
  assign n964 = (~x2 & n61) | (~x2 & n963) | (n61 & n963);
  assign n965 = x1 & ~n964;
  assign n960 = (x2 & x5) | (x2 & x7) | (x5 & x7);
  assign n961 = x4 & n960;
  assign n962 = (n73 & n755) | (n73 & ~n961) | (n755 & ~n961);
  assign n966 = x1 | n962;
  assign n967 = (~x1 & n965) | (~x1 & n966) | (n965 & n966);
  assign n991 = x0 | n967;
  assign n992 = x3 & n991;
  assign n993 = n990 & ~n992;
  assign n1091 = (x6 & x8) | (x6 & n993) | (x8 & n993);
  assign n1092 = (~n994 & n1090) | (~n994 & n1091) | (n1090 & n1091);
  assign n930 = (~x1 & x2) | (~x1 & x5) | (x2 & x5);
  assign n931 = (x5 & x7) | (x5 & ~n930) | (x7 & ~n930);
  assign n932 = (~x2 & x7) | (~x2 & n930) | (x7 & n930);
  assign n933 = n931 & ~n932;
  assign n953 = x0 & n933;
  assign n934 = x7 & n44;
  assign n935 = (x2 & x5) | (x2 & n934) | (x5 & n934);
  assign n936 = ~x2 & n935;
  assign n942 = (x0 & x1) | (x0 & x4) | (x1 & x4);
  assign n943 = (x0 & x7) | (x0 & ~n942) | (x7 & ~n942);
  assign n944 = (~x1 & x7) | (~x1 & n942) | (x7 & n942);
  assign n945 = ~n943 & n944;
  assign n946 = (x0 & x1) | (x0 & ~n945) | (x1 & ~n945);
  assign n947 = n941 & n946;
  assign n948 = (n941 & n945) | (n941 & ~n947) | (n945 & ~n947);
  assign n949 = x2 | n948;
  assign n937 = (x1 & x4) | (x1 & ~x7) | (x4 & ~x7);
  assign n938 = (~x4 & x5) | (~x4 & n937) | (x5 & n937);
  assign n939 = (x1 & x5) | (x1 & ~n937) | (x5 & ~n937);
  assign n940 = n938 & ~n939;
  assign n950 = ~x0 & n940;
  assign n951 = x2 & ~n950;
  assign n952 = n949 & ~n951;
  assign n954 = n936 | n952;
  assign n955 = (n933 & ~n953) | (n933 & n954) | (~n953 & n954);
  assign n956 = x3 | n955;
  assign n920 = x2 & ~x7;
  assign n921 = (~x2 & n61) | (~x2 & n920) | (n61 & n920);
  assign n927 = x1 & n921;
  assign n922 = (x2 & ~x4) | (x2 & x7) | (~x4 & x7);
  assign n923 = (x5 & ~x7) | (x5 & n922) | (~x7 & n922);
  assign n924 = (x2 & ~x4) | (x2 & n923) | (~x4 & n923);
  assign n925 = ~n922 & n924;
  assign n926 = (~n923 & n924) | (~n923 & n925) | (n924 & n925);
  assign n928 = x1 | n926;
  assign n929 = (~x1 & n927) | (~x1 & n928) | (n927 & n928);
  assign n957 = ~x0 & n929;
  assign n958 = x3 & ~n957;
  assign n959 = n956 & ~n958;
  assign n1093 = n959 | n1092;
  assign n1094 = (~n738 & n1092) | (~n738 & n1093) | (n1092 & n1093);
  assign n1132 = x0 & ~x6;
  assign n1133 = (~x4 & x7) | (~x4 & n1132) | (x7 & n1132);
  assign n1134 = (x6 & ~x7) | (x6 & n1132) | (~x7 & n1132);
  assign n1135 = (~x0 & x4) | (~x0 & n1134) | (x4 & n1134);
  assign n1136 = n1133 | n1135;
  assign n1137 = ~x3 & n1136;
  assign n1131 = ~x4 & n552;
  assign n1138 = ~x0 & n1131;
  assign n1139 = x3 & ~n1138;
  assign n1140 = n1137 | n1139;
  assign n1141 = ~x2 & n1140;
  assign n1127 = (x3 & x4) | (x3 & ~x7) | (x4 & ~x7);
  assign n1128 = (~x3 & x6) | (~x3 & n1127) | (x6 & n1127);
  assign n1129 = (~x6 & x7) | (~x6 & n1127) | (x7 & n1127);
  assign n1130 = n1128 & n1129;
  assign n1142 = ~x0 & n1130;
  assign n1143 = x2 & ~n1142;
  assign n1144 = n1141 | n1143;
  assign n1145 = ~x1 & n1144;
  assign n1122 = x4 & n186;
  assign n1123 = x2 & ~n1122;
  assign n1121 = ~x4 & n583;
  assign n1124 = ~x3 & n1121;
  assign n1125 = x2 | n1124;
  assign n1126 = ~n1123 & n1125;
  assign n1146 = ~x0 & n1126;
  assign n1147 = x1 & ~n1146;
  assign n1148 = n1145 | n1147;
  assign n1282 = n656 | n1148;
  assign n1163 = (~x0 & x5) | (~x0 & x7) | (x5 & x7);
  assign n1164 = (x7 & x8) | (x7 & ~n1163) | (x8 & ~n1163);
  assign n1165 = (x0 & ~x5) | (x0 & n1164) | (~x5 & n1164);
  assign n1166 = n1163 & n1165;
  assign n1167 = (~n1164 & n1165) | (~n1164 & n1166) | (n1165 & n1166);
  assign n1168 = ~x4 & n1167;
  assign n1169 = x1 | n1168;
  assign n1161 = x7 & ~n656;
  assign n1162 = x4 & n1161;
  assign n1170 = ~x0 & n1162;
  assign n1171 = x1 & ~n1170;
  assign n1172 = n1169 & ~n1171;
  assign n1173 = x3 | n1172;
  assign n1159 = x1 & ~n61;
  assign n1160 = (n60 & n61) | (n60 & n1159) | (n61 & n1159);
  assign n1174 = ~x0 & n1160;
  assign n1175 = x3 & ~n1174;
  assign n1176 = n1173 & ~n1175;
  assign n1177 = x2 | n1176;
  assign n1154 = (x4 & n60) | (x4 & ~n765) | (n60 & ~n765);
  assign n1155 = ~x3 & n1154;
  assign n1156 = x1 & n1155;
  assign n1149 = (x1 & x7) | (x1 & ~x8) | (x7 & ~x8);
  assign n1150 = (x5 & ~x8) | (x5 & n1149) | (~x8 & n1149);
  assign n1151 = x8 & n1150;
  assign n1152 = n1150 & ~n1151;
  assign n1153 = (x8 & ~n1151) | (x8 & n1152) | (~n1151 & n1152);
  assign n1157 = (~x3 & x4) | (~x3 & n1153) | (x4 & n1153);
  assign n1158 = (n80 & ~n1156) | (n80 & n1157) | (~n1156 & n1157);
  assign n1178 = x0 | n1158;
  assign n1179 = x2 & n1178;
  assign n1180 = n1177 & ~n1179;
  assign n1222 = (n54 & ~n591) | (n54 & n684) | (~n591 & n684);
  assign n1224 = x3 & ~n164;
  assign n1225 = ~n1222 & n1224;
  assign n1223 = ~x5 & n994;
  assign n1226 = (~n164 & n1223) | (~n164 & n1224) | (n1223 & n1224);
  assign n1227 = (x4 & n1225) | (x4 & n1226) | (n1225 & n1226);
  assign n1228 = x2 | n1227;
  assign n1221 = ~x5 & n684;
  assign n1229 = n20 & n1221;
  assign n1230 = x2 & ~n1229;
  assign n1231 = n1228 & ~n1230;
  assign n1250 = (x6 & x7) | (x6 & n86) | (x7 & n86);
  assign n1251 = (x6 & ~x8) | (x6 & n86) | (~x8 & n86);
  assign n1252 = (n28 & ~n1250) | (n28 & n1251) | (~n1250 & n1251);
  assign n1253 = x5 & n1252;
  assign n1254 = x4 & n882;
  assign n1255 = x5 | n1254;
  assign n1256 = ~n1253 & n1255;
  assign n1257 = x2 & ~n1256;
  assign n1258 = n16 & n572;
  assign n1259 = x2 | n1258;
  assign n1260 = ~n1257 & n1259;
  assign n1262 = (x2 & x4) | (x2 & x7) | (x4 & x7);
  assign n1263 = (x2 & x3) | (x2 & ~n1262) | (x3 & ~n1262);
  assign n1264 = (x4 & x7) | (x4 & ~n1263) | (x7 & ~n1263);
  assign n1265 = ~n1262 & n1264;
  assign n1266 = (n1263 & n1264) | (n1263 & n1265) | (n1264 & n1265);
  assign n1261 = x5 & n70;
  assign n1267 = n1261 & n1266;
  assign n1268 = (n1221 & n1266) | (n1221 & n1267) | (n1266 & n1267);
  assign n1269 = (~x3 & n1260) | (~x3 & n1268) | (n1260 & n1268);
  assign n1236 = x2 & ~x6;
  assign n1237 = x7 & n73;
  assign n1238 = (n583 & n1236) | (n583 & ~n1237) | (n1236 & ~n1237);
  assign n1239 = (x2 & x4) | (x2 & ~x6) | (x4 & ~x6);
  assign n1240 = (x2 & ~x7) | (x2 & n1239) | (~x7 & n1239);
  assign n1241 = x2 & ~n1240;
  assign n1242 = n1240 | n1241;
  assign n1243 = (~x2 & n1241) | (~x2 & n1242) | (n1241 & n1242);
  assign n1244 = x8 | n1243;
  assign n1245 = (n1238 & n1243) | (n1238 & n1244) | (n1243 & n1244);
  assign n1246 = x5 | n1245;
  assign n1232 = (x6 & x7) | (x6 & ~x8) | (x7 & ~x8);
  assign n1233 = (x2 & ~x6) | (x2 & x8) | (~x6 & x8);
  assign n1234 = x7 & ~n1233;
  assign n1235 = n1232 & ~n1234;
  assign n1247 = ~x4 & n1235;
  assign n1248 = x5 & ~n1247;
  assign n1249 = n1246 & ~n1248;
  assign n1270 = (x3 & n1249) | (x3 & n1268) | (n1249 & n1268);
  assign n1271 = n1269 | n1270;
  assign n1272 = x0 & n16;
  assign n1273 = (n45 & ~n375) | (n45 & n1272) | (~n375 & n1272);
  assign n1274 = ~n45 & n1273;
  assign n1275 = (~n1231 & n1271) | (~n1231 & n1274) | (n1271 & n1274);
  assign n1276 = x0 & ~n1274;
  assign n1277 = (n1231 & n1275) | (n1231 & ~n1276) | (n1275 & ~n1276);
  assign n1278 = x1 | n1277;
  assign n1206 = (x2 & ~x4) | (x2 & x5) | (~x4 & x5);
  assign n1207 = (x2 & ~x7) | (x2 & n1206) | (~x7 & n1206);
  assign n1208 = x2 & ~n1207;
  assign n1209 = n1207 | n1208;
  assign n1210 = (~x2 & n1208) | (~x2 & n1209) | (n1208 & n1209);
  assign n1211 = x8 & n1210;
  assign n1203 = (x7 & n519) | (x7 & ~n765) | (n519 & ~n765);
  assign n1204 = (x2 & ~x7) | (x2 & n765) | (~x7 & n765);
  assign n1205 = (~x2 & n1203) | (~x2 & n1204) | (n1203 & n1204);
  assign n1212 = x8 | n1205;
  assign n1213 = (~x8 & n1211) | (~x8 & n1212) | (n1211 & n1212);
  assign n1214 = x3 & ~n1213;
  assign n1200 = (x4 & ~x5) | (x4 & x8) | (~x5 & x8);
  assign n1201 = ~x2 & n1200;
  assign n1202 = (n411 & n717) | (n411 & ~n1201) | (n717 & ~n1201);
  assign n1215 = x7 | n1202;
  assign n1216 = ~x3 & n1215;
  assign n1217 = n1214 | n1216;
  assign n1218 = x6 & ~n1217;
  assign n1188 = (x2 & x5) | (x2 & ~n501) | (x5 & ~n501);
  assign n1189 = (~x5 & x7) | (~x5 & n1188) | (x7 & n1188);
  assign n1190 = n501 | n1189;
  assign n1191 = (~x2 & n1188) | (~x2 & n1190) | (n1188 & n1190);
  assign n1192 = x3 & n1191;
  assign n1185 = (x5 & x7) | (x5 & ~x8) | (x7 & ~x8);
  assign n1186 = x8 & n1185;
  assign n1187 = (~n755 & n1185) | (~n755 & n1186) | (n1185 & n1186);
  assign n1193 = ~x2 & n1187;
  assign n1194 = x3 | n1193;
  assign n1195 = ~n1192 & n1194;
  assign n1196 = x4 | n1195;
  assign n1181 = (x2 & x3) | (x2 & ~n755) | (x3 & ~n755);
  assign n1182 = (~x2 & x5) | (~x2 & n1181) | (x5 & n1181);
  assign n1183 = (~x3 & x7) | (~x3 & n1182) | (x7 & n1182);
  assign n1184 = n1181 & n1183;
  assign n1197 = ~x8 & n1184;
  assign n1198 = x4 & ~n1197;
  assign n1199 = n1196 & ~n1198;
  assign n1219 = x6 | n1199;
  assign n1220 = (~x6 & n1218) | (~x6 & n1219) | (n1218 & n1219);
  assign n1279 = ~x0 & n1220;
  assign n1280 = x1 & ~n1279;
  assign n1281 = n1278 & ~n1280;
  assign n1283 = n1180 | n1281;
  assign n1284 = (~n1148 & n1282) | (~n1148 & n1283) | (n1282 & n1283);
  assign n1104 = ~x0 & x2;
  assign n1107 = x0 & ~x5;
  assign n1108 = (~n178 & n1104) | (~n178 & n1107) | (n1104 & n1107);
  assign n1109 = x6 | n1108;
  assign n1105 = ~x0 & x4;
  assign n1106 = (n272 & n1104) | (n272 & ~n1105) | (n1104 & ~n1105);
  assign n1110 = ~x5 & n1106;
  assign n1111 = x6 & ~n1110;
  assign n1112 = n1109 & ~n1111;
  assign n1113 = x1 | n1112;
  assign n1102 = x6 & ~n519;
  assign n1103 = (n37 & n118) | (n37 & ~n1102) | (n118 & ~n1102);
  assign n1114 = ~x0 & n1103;
  assign n1115 = x1 & ~n1114;
  assign n1116 = n1113 & ~n1115;
  assign n1117 = x3 | n1116;
  assign n1095 = (x1 & x4) | (x1 & ~n765) | (x4 & ~n765);
  assign n1096 = (x1 & x2) | (x1 & ~n765) | (x2 & ~n765);
  assign n1097 = (n519 & n1095) | (n519 & ~n1096) | (n1095 & ~n1096);
  assign n1098 = ~x6 & n16;
  assign n1099 = n487 & n1098;
  assign n1100 = x6 | n1099;
  assign n1101 = (n1097 & n1099) | (n1097 & n1100) | (n1099 & n1100);
  assign n1118 = ~x0 & n1101;
  assign n1119 = x3 & ~n1118;
  assign n1120 = n1117 & ~n1119;
  assign n1285 = n1120 | n1284;
  assign n1286 = (n29 & n1284) | (n29 & n1285) | (n1284 & n1285);
  assign n1287 = x2 | x6;
  assign n1288 = (~n147 & n377) | (~n147 & n1287) | (n377 & n1287);
  assign n1289 = x1 & ~n1288;
  assign n1290 = ~x0 & n1289;
  assign n1291 = (x2 & n44) | (x2 & n463) | (n44 & n463);
  assign n1292 = ~x2 & n1291;
  assign n1293 = x4 & ~n15;
  assign n1294 = (x6 & x7) | (x6 & n1293) | (x7 & n1293);
  assign n1295 = ~x7 & n1294;
  assign n1296 = n39 | n1295;
  assign n1297 = (n1131 & n1295) | (n1131 & n1296) | (n1295 & n1296);
  assign n1321 = x0 & n1297;
  assign n1298 = ~x4 & n318;
  assign n1299 = ~n564 & n1298;
  assign n1305 = (x6 & ~x7) | (x6 & n922) | (~x7 & n922);
  assign n1306 = (x2 & x6) | (x2 & ~n922) | (x6 & ~n922);
  assign n1307 = n1305 & ~n1306;
  assign n1311 = (x0 & x8) | (x0 & n1307) | (x8 & n1307);
  assign n1308 = x0 & x4;
  assign n1309 = (x2 & ~n564) | (x2 & n1308) | (~n564 & n1308);
  assign n1310 = ~x2 & n1309;
  assign n1312 = x8 & n1310;
  assign n1313 = (~x0 & n1311) | (~x0 & n1312) | (n1311 & n1312);
  assign n1302 = (~x4 & x6) | (~x4 & x7) | (x6 & x7);
  assign n1303 = (~x4 & x6) | (~x4 & x8) | (x6 & x8);
  assign n1304 = n1302 & ~n1303;
  assign n1314 = (~x0 & n1304) | (~x0 & n1313) | (n1304 & n1313);
  assign n1315 = x2 & ~n1314;
  assign n1316 = (x2 & n1313) | (x2 & ~n1315) | (n1313 & ~n1315);
  assign n1317 = x1 | n1316;
  assign n1300 = (~x2 & x8) | (~x2 & n379) | (x8 & n379);
  assign n1301 = n500 & n1300;
  assign n1318 = ~x0 & n1301;
  assign n1319 = x1 & ~n1318;
  assign n1320 = n1317 & ~n1319;
  assign n1322 = n1299 | n1320;
  assign n1323 = (n1297 & ~n1321) | (n1297 & n1322) | (~n1321 & n1322);
  assign n1324 = (~n1290 & n1292) | (~n1290 & n1323) | (n1292 & n1323);
  assign n1325 = n29 & ~n1323;
  assign n1326 = (n1290 & n1324) | (n1290 & ~n1325) | (n1324 & ~n1325);
  assign n1477 = x3 & n1326;
  assign n1336 = (x1 & x2) | (x1 & x4) | (x2 & x4);
  assign n1337 = (x2 & x6) | (x2 & ~n1336) | (x6 & ~n1336);
  assign n1338 = (x1 & x4) | (x1 & ~n1337) | (x4 & ~n1337);
  assign n1339 = n1336 & ~n1338;
  assign n1340 = (n1337 & n1338) | (n1337 & ~n1339) | (n1338 & ~n1339);
  assign n1345 = (~x7 & x8) | (~x7 & n1340) | (x8 & n1340);
  assign n1341 = ~x2 & x6;
  assign n1342 = (x2 & x4) | (x2 & n1341) | (x4 & n1341);
  assign n1343 = (x1 & x4) | (x1 & n1341) | (x4 & n1341);
  assign n1344 = (n487 & n1342) | (n487 & ~n1343) | (n1342 & ~n1343);
  assign n1346 = (x7 & x8) | (x7 & ~n1344) | (x8 & ~n1344);
  assign n1347 = n1345 | n1346;
  assign n1327 = (~x2 & x4) | (~x2 & n884) | (x4 & n884);
  assign n1328 = (x4 & x6) | (x4 & ~n884) | (x6 & ~n884);
  assign n1329 = n1327 & ~n1328;
  assign n1333 = (x1 & x8) | (x1 & ~n1329) | (x8 & ~n1329);
  assign n1330 = (x2 & x4) | (x2 & ~n94) | (x4 & ~n94);
  assign n1331 = (~x1 & x4) | (~x1 & n94) | (x4 & n94);
  assign n1332 = n1330 & ~n1331;
  assign n1334 = x8 & n1332;
  assign n1335 = (n1329 & n1333) | (n1329 & n1334) | (n1333 & n1334);
  assign n1348 = n1335 & n1347;
  assign n1349 = ~x0 & x3;
  assign n1350 = (~n1347 & n1348) | (~n1347 & n1349) | (n1348 & n1349);
  assign n1351 = (~x1 & n20) | (~x1 & n632) | (n20 & n632);
  assign n1352 = x1 & n1073;
  assign n1353 = (n20 & ~n1351) | (n20 & n1352) | (~n1351 & n1352);
  assign n1358 = (x0 & ~x2) | (x0 & n1353) | (~x2 & n1353);
  assign n1354 = x1 | x3;
  assign n1355 = x0 & ~n1354;
  assign n1356 = x4 & n591;
  assign n1357 = n1355 & n1356;
  assign n1359 = ~x2 & n1357;
  assign n1360 = (~x0 & n1358) | (~x0 & n1359) | (n1358 & n1359);
  assign n1361 = (n40 & n164) | (n40 & n1360) | (n164 & n1360);
  assign n1362 = n591 & ~n1361;
  assign n1363 = (n591 & n1360) | (n591 & ~n1362) | (n1360 & ~n1362);
  assign n1474 = n29 & n1363;
  assign n1375 = n46 & ~n375;
  assign n1376 = n118 & n1375;
  assign n1369 = ~x4 & n591;
  assign n1370 = (x1 & n232) | (x1 & n1369) | (n232 & n1369);
  assign n1371 = ~x1 & n1370;
  assign n1364 = (x1 & ~x3) | (x1 & x4) | (~x3 & x4);
  assign n1365 = (x1 & x6) | (x1 & ~n1364) | (x6 & ~n1364);
  assign n1366 = (x3 & ~x4) | (x3 & n1365) | (~x4 & n1365);
  assign n1367 = n1364 | n1366;
  assign n1368 = (~n1365 & n1366) | (~n1365 & n1367) | (n1366 & n1367);
  assign n1372 = (x2 & n1368) | (x2 & ~n1371) | (n1368 & ~n1371);
  assign n1373 = ~x5 & n1372;
  assign n1374 = (x5 & ~n1371) | (x5 & n1373) | (~n1371 & n1373);
  assign n1377 = (x0 & n1374) | (x0 & ~n1376) | (n1374 & ~n1376);
  assign n1378 = x8 & n1377;
  assign n1379 = (x8 & n1376) | (x8 & ~n1378) | (n1376 & ~n1378);
  assign n1417 = x1 & ~n487;
  assign n1418 = n376 & n1417;
  assign n1416 = ~x4 & n994;
  assign n1419 = (~n487 & n1416) | (~n487 & n1417) | (n1416 & n1417);
  assign n1420 = (~x2 & n1418) | (~x2 & n1419) | (n1418 & n1419);
  assign n1415 = (~x3 & n398) | (~x3 & n618) | (n398 & n618);
  assign n1465 = n1415 & n1420;
  assign n1384 = (x2 & x3) | (x2 & x5) | (x3 & x5);
  assign n1421 = (x3 & ~x4) | (x3 & n1384) | (~x4 & n1384);
  assign n1422 = x3 & ~n1421;
  assign n1423 = n1421 | n1422;
  assign n1424 = (~x3 & n1422) | (~x3 & n1423) | (n1422 & n1423);
  assign n1425 = (x1 & ~x8) | (x1 & n1424) | (~x8 & n1424);
  assign n1426 = x8 & n1425;
  assign n1427 = (x1 & x6) | (x1 & ~n1426) | (x6 & ~n1426);
  assign n1428 = (n1425 & n1426) | (n1425 & ~n1427) | (n1426 & ~n1427);
  assign n1448 = (x2 & x3) | (x2 & ~x4) | (x3 & ~x4);
  assign n1449 = (x4 & x6) | (x4 & n1448) | (x6 & n1448);
  assign n1450 = (x2 & x3) | (x2 & n1449) | (x3 & n1449);
  assign n1451 = ~n1448 & n1450;
  assign n1452 = (~n1449 & n1450) | (~n1449 & n1451) | (n1450 & n1451);
  assign n1453 = x5 & ~n1452;
  assign n1454 = ~x3 & n379;
  assign n1455 = x5 | n1454;
  assign n1456 = ~n1453 & n1455;
  assign n1457 = x1 | n1456;
  assign n1458 = ~n45 & n1356;
  assign n1459 = x1 & ~n1458;
  assign n1460 = n1457 & ~n1459;
  assign n1461 = ~x8 & n1460;
  assign n1429 = (x2 & x6) | (x2 & n111) | (x6 & n111);
  assign n1430 = (x5 & x6) | (x5 & ~n1429) | (x6 & ~n1429);
  assign n1431 = n111 | n1430;
  assign n1432 = (x2 & ~n1429) | (x2 & n1431) | (~n1429 & n1431);
  assign n1434 = (~x1 & x3) | (~x1 & n1432) | (x3 & n1432);
  assign n1433 = n416 & ~n632;
  assign n1435 = ~x1 & n1433;
  assign n1436 = (~n1432 & n1434) | (~n1432 & n1435) | (n1434 & n1435);
  assign n1437 = x3 & x6;
  assign n1438 = (~x2 & x5) | (~x2 & n1437) | (x5 & n1437);
  assign n1439 = (x5 & x6) | (x5 & ~n1437) | (x6 & ~n1437);
  assign n1440 = (~x2 & x3) | (~x2 & n1439) | (x3 & n1439);
  assign n1441 = ~n1438 & n1440;
  assign n1445 = (~x1 & x4) | (~x1 & n1441) | (x4 & n1441);
  assign n1442 = (~x5 & n632) | (~x5 & n851) | (n632 & n851);
  assign n1443 = (x2 & n20) | (x2 & n1442) | (n20 & n1442);
  assign n1444 = ~n1442 & n1443;
  assign n1446 = x1 & n1444;
  assign n1447 = (n1441 & ~n1445) | (n1441 & n1446) | (~n1445 & n1446);
  assign n1462 = n1436 | n1447;
  assign n1463 = x8 & n1462;
  assign n1464 = n1461 | n1463;
  assign n1466 = n1428 | n1464;
  assign n1467 = (n1420 & ~n1465) | (n1420 & n1466) | (~n1465 & n1466);
  assign n1468 = (~x0 & x7) | (~x0 & n1467) | (x7 & n1467);
  assign n1392 = (x1 & x3) | (x1 & x6) | (x3 & x6);
  assign n1393 = (x3 & n591) | (x3 & ~n1392) | (n591 & ~n1392);
  assign n1394 = (~x5 & n1392) | (~x5 & n1393) | (n1392 & n1393);
  assign n1395 = (~x3 & n1393) | (~x3 & n1394) | (n1393 & n1394);
  assign n1399 = (~x2 & x8) | (~x2 & n1395) | (x8 & n1395);
  assign n1396 = x6 | n15;
  assign n1397 = (x3 & x5) | (x3 & ~n1396) | (x5 & ~n1396);
  assign n1398 = ~x3 & n1397;
  assign n1400 = ~x8 & n1398;
  assign n1401 = (n1395 & ~n1399) | (n1395 & n1400) | (~n1399 & n1400);
  assign n1402 = (~x1 & n1261) | (~x1 & n1401) | (n1261 & n1401);
  assign n1403 = n812 & ~n1402;
  assign n1404 = (n812 & n1401) | (n812 & ~n1403) | (n1401 & ~n1403);
  assign n1405 = (x3 & x8) | (x3 & ~n810) | (x8 & ~n810);
  assign n1406 = (x3 & x5) | (x3 & ~n810) | (x5 & ~n810);
  assign n1407 = (n655 & n1405) | (n655 & ~n1406) | (n1405 & ~n1406);
  assign n1408 = (x2 & x6) | (x2 & n1407) | (x6 & n1407);
  assign n1409 = (x1 & ~x2) | (x1 & n1408) | (~x2 & n1408);
  assign n1410 = (x1 & x6) | (x1 & ~n1408) | (x6 & ~n1408);
  assign n1411 = n1409 & ~n1410;
  assign n1412 = (~x4 & n1404) | (~x4 & n1411) | (n1404 & n1411);
  assign n1380 = (x3 & ~x6) | (x3 & n1287) | (~x6 & n1287);
  assign n1381 = (x3 & ~x5) | (x3 & n1287) | (~x5 & n1287);
  assign n1382 = (n851 & ~n1380) | (n851 & n1381) | (~n1380 & n1381);
  assign n1387 = x1 & x8;
  assign n1388 = x8 & ~n1387;
  assign n1389 = n1382 & n1388;
  assign n1383 = (x2 & x5) | (x2 & x6) | (x5 & x6);
  assign n1385 = ~x3 & x6;
  assign n1386 = (~n1383 & n1384) | (~n1383 & n1385) | (n1384 & n1385);
  assign n1390 = (n1386 & ~n1387) | (n1386 & n1388) | (~n1387 & n1388);
  assign n1391 = (x1 & n1389) | (x1 & n1390) | (n1389 & n1390);
  assign n1413 = (x4 & n1391) | (x4 & n1411) | (n1391 & n1411);
  assign n1414 = n1412 | n1413;
  assign n1469 = (x0 & x7) | (x0 & ~n1414) | (x7 & ~n1414);
  assign n1470 = n1468 & ~n1469;
  assign n1471 = (n46 & n257) | (n46 & n1470) | (n257 & n1470);
  assign n1472 = n61 & ~n1471;
  assign n1473 = (n61 & n1470) | (n61 & ~n1472) | (n1470 & ~n1472);
  assign n1475 = n1379 | n1473;
  assign n1476 = (n1363 & ~n1474) | (n1363 & n1475) | (~n1474 & n1475);
  assign n1478 = n1350 | n1476;
  assign n1479 = (n1326 & ~n1477) | (n1326 & n1478) | (~n1477 & n1478);
  assign n1519 = ~x3 & n351;
  assign n1520 = (x1 & ~x4) | (x1 & n1519) | (~x4 & n1519);
  assign n1521 = (n351 & n1519) | (n351 & n1520) | (n1519 & n1520);
  assign n1524 = x6 & n1521;
  assign n1522 = x1 | x8;
  assign n1523 = (n712 & ~n887) | (n712 & n1522) | (~n887 & n1522);
  assign n1525 = (x3 & x6) | (x3 & ~n1523) | (x6 & ~n1523);
  assign n1526 = (~n1437 & n1524) | (~n1437 & n1525) | (n1524 & n1525);
  assign n1527 = x5 & ~n1526;
  assign n1515 = (x4 & x6) | (x4 & ~x8) | (x6 & ~x8);
  assign n1516 = ~x4 & n1515;
  assign n1517 = (~x3 & x8) | (~x3 & n1516) | (x8 & n1516);
  assign n1518 = (n1515 & n1516) | (n1515 & n1517) | (n1516 & n1517);
  assign n1528 = x1 & n1518;
  assign n1529 = x5 | n1528;
  assign n1530 = ~n1527 & n1529;
  assign n1553 = (x2 & ~x7) | (x2 & n1530) | (~x7 & n1530);
  assign n1542 = x3 & ~n54;
  assign n1543 = (x5 & x6) | (x5 & ~n54) | (x6 & ~n54);
  assign n1544 = (x3 & n632) | (x3 & ~n1543) | (n632 & ~n1543);
  assign n1545 = (~x3 & n1542) | (~x3 & n1544) | (n1542 & n1544);
  assign n1546 = x1 | n1545;
  assign n1541 = x5 & ~n375;
  assign n1547 = ~x3 & n1541;
  assign n1548 = x1 & ~n1547;
  assign n1549 = n1546 & ~n1548;
  assign n1550 = x4 & n1549;
  assign n1532 = (x1 & ~x3) | (x1 & x6) | (~x3 & x6);
  assign n1533 = (x3 & x5) | (x3 & n1532) | (x5 & n1532);
  assign n1534 = x3 & n1532;
  assign n1535 = x5 | n1532;
  assign n1536 = (~n1533 & n1534) | (~n1533 & n1535) | (n1534 & n1535);
  assign n1537 = x8 & ~n1536;
  assign n1531 = (n53 & n96) | (n53 & ~n573) | (n96 & ~n573);
  assign n1538 = x6 & n1531;
  assign n1539 = x8 | n1538;
  assign n1540 = ~n1537 & n1539;
  assign n1551 = x4 | n1540;
  assign n1552 = (~x4 & n1550) | (~x4 & n1551) | (n1550 & n1551);
  assign n1554 = (x2 & x7) | (x2 & n1552) | (x7 & n1552);
  assign n1555 = n1553 & n1554;
  assign n1661 = x0 & n1555;
  assign n1558 = n1121 & ~n1354;
  assign n1556 = (x3 & n564) | (x3 & n887) | (n564 & n887);
  assign n1557 = ~n564 & n1556;
  assign n1559 = n1557 | n1558;
  assign n1560 = (~x0 & n1558) | (~x0 & n1559) | (n1558 & n1559);
  assign n1620 = (x2 & n656) | (x2 & n1560) | (n656 & n1560);
  assign n1593 = (n53 & ~n299) | (n53 & n717) | (~n299 & n717);
  assign n1594 = x7 & n1593;
  assign n1598 = x3 & x8;
  assign n1599 = (x4 & ~x5) | (x4 & n1598) | (~x5 & n1598);
  assign n1600 = (~x3 & x5) | (~x3 & n1599) | (x5 & n1599);
  assign n1601 = (x4 & x8) | (x4 & ~n1600) | (x8 & ~n1600);
  assign n1602 = ~n1599 & n1601;
  assign n1603 = x7 | n1602;
  assign n1595 = x5 & n153;
  assign n1596 = x5 | n810;
  assign n1597 = ~n1595 & n1596;
  assign n1604 = x3 & ~n1597;
  assign n1605 = x7 & ~n1604;
  assign n1606 = n1603 & ~n1605;
  assign n1607 = ~x3 & n139;
  assign n1608 = x0 & n1607;
  assign n1609 = (~n1594 & n1606) | (~n1594 & n1608) | (n1606 & n1608);
  assign n1610 = x0 & ~n1608;
  assign n1611 = (n1594 & n1609) | (n1594 & ~n1610) | (n1609 & ~n1610);
  assign n1612 = x6 & ~n1611;
  assign n1585 = (x3 & ~n790) | (x3 & n810) | (~n790 & n810);
  assign n1586 = (~x3 & x7) | (~x3 & n1585) | (x7 & n1585);
  assign n1587 = (~x4 & n810) | (~x4 & n1586) | (n810 & n1586);
  assign n1588 = (~n810 & n1585) | (~n810 & n1587) | (n1585 & n1587);
  assign n1589 = x5 & n1588;
  assign n1582 = (x3 & x7) | (x3 & x8) | (x7 & x8);
  assign n1583 = ~x3 & n1582;
  assign n1584 = (~n60 & n1582) | (~n60 & n1583) | (n1582 & n1583);
  assign n1590 = x4 & n1584;
  assign n1591 = x5 | n1590;
  assign n1592 = ~n1589 & n1591;
  assign n1613 = ~x0 & n1592;
  assign n1614 = x6 | n1613;
  assign n1615 = ~n1612 & n1614;
  assign n1616 = x1 | n1615;
  assign n1571 = (x3 & ~x4) | (x3 & x7) | (~x4 & x7);
  assign n1572 = (x3 & ~x6) | (x3 & n1571) | (~x6 & n1571);
  assign n1573 = x3 & ~n1572;
  assign n1574 = n1572 | n1573;
  assign n1575 = (~x3 & n1573) | (~x3 & n1574) | (n1573 & n1574);
  assign n1576 = x8 & n1575;
  assign n1568 = (x4 & x6) | (x4 & ~x7) | (x6 & ~x7);
  assign n1569 = x4 & ~n1568;
  assign n1570 = (n552 & n1568) | (n552 & ~n1569) | (n1568 & ~n1569);
  assign n1577 = ~x8 & n1570;
  assign n1578 = (x8 & ~n1576) | (x8 & n1577) | (~n1576 & n1577);
  assign n1579 = x5 & ~n1578;
  assign n1561 = x3 | x7;
  assign n1562 = x6 & n1561;
  assign n1563 = (n60 & n684) | (n60 & ~n1562) | (n684 & ~n1562);
  assign n1565 = ~x4 & n1563;
  assign n1564 = (n10 & n375) | (n10 & ~n583) | (n375 & ~n583);
  assign n1566 = (x3 & x4) | (x3 & n1564) | (x4 & n1564);
  assign n1567 = (n36 & n1565) | (n36 & ~n1566) | (n1565 & ~n1566);
  assign n1580 = x5 | n1567;
  assign n1581 = (~x5 & n1579) | (~x5 & n1580) | (n1579 & n1580);
  assign n1617 = ~x0 & n1581;
  assign n1618 = x1 & ~n1617;
  assign n1619 = n1616 & ~n1618;
  assign n1621 = ~x2 & n1619;
  assign n1622 = (n1560 & ~n1620) | (n1560 & n1621) | (~n1620 & n1621);
  assign n1644 = ~n394 & n1239;
  assign n1647 = (~x0 & x1) | (~x0 & n1644) | (x1 & n1644);
  assign n1645 = x4 & n37;
  assign n1646 = n487 & n1645;
  assign n1648 = ~x0 & n1646;
  assign n1649 = (~x1 & n1647) | (~x1 & n1648) | (n1647 & n1648);
  assign n1650 = (~n40 & n318) | (~n40 & n1649) | (n318 & n1649);
  assign n1643 = (n16 & n37) | (n16 & ~n463) | (n37 & ~n463);
  assign n1651 = n1643 | n1649;
  assign n1652 = (n40 & n1650) | (n40 & n1651) | (n1650 & n1651);
  assign n1653 = x8 | n1652;
  assign n1635 = (x2 & ~x4) | (x2 & x6) | (~x4 & x6);
  assign n1636 = (x2 & ~x5) | (x2 & n1635) | (~x5 & n1635);
  assign n1637 = x2 & ~n1636;
  assign n1638 = n1636 | n1637;
  assign n1639 = (~x2 & n1637) | (~x2 & n1638) | (n1637 & n1638);
  assign n1640 = x1 & n1639;
  assign n1631 = (x2 & ~x4) | (x2 & n702) | (~x4 & n702);
  assign n1632 = (x5 & x6) | (x5 & n1631) | (x6 & n1631);
  assign n1633 = n702 & ~n1632;
  assign n1634 = (n1631 & ~n1632) | (n1631 & n1633) | (~n1632 & n1633);
  assign n1641 = x1 | n1634;
  assign n1642 = (~x1 & n1640) | (~x1 & n1641) | (n1640 & n1641);
  assign n1654 = ~x0 & n1642;
  assign n1655 = x8 & ~n1654;
  assign n1656 = n1653 & ~n1655;
  assign n1657 = x3 | n1656;
  assign n1626 = (x2 & n887) | (x2 & n1221) | (n887 & n1221);
  assign n1627 = ~x2 & n1626;
  assign n1623 = (x1 & x4) | (x1 & x8) | (x4 & x8);
  assign n1624 = (x6 & x8) | (x6 & n887) | (x8 & n887);
  assign n1625 = n1623 & ~n1624;
  assign n1628 = (x2 & n1625) | (x2 & n1627) | (n1625 & n1627);
  assign n1629 = x5 & ~n1628;
  assign n1630 = (x5 & n1627) | (x5 & ~n1629) | (n1627 & ~n1629);
  assign n1658 = ~x0 & n1630;
  assign n1659 = x3 & ~n1658;
  assign n1660 = n1657 & ~n1659;
  assign n1662 = n1622 | n1660;
  assign n1663 = (n1555 & ~n1661) | (n1555 & n1662) | (~n1661 & n1662);
  assign n1480 = (x1 & x3) | (x1 & x7) | (x3 & x7);
  assign n1481 = (x1 & x4) | (x1 & x7) | (x4 & x7);
  assign n1482 = (n80 & ~n1480) | (n80 & n1481) | (~n1480 & n1481);
  assign n1486 = (x2 & x8) | (x2 & ~n1482) | (x8 & ~n1482);
  assign n1483 = x1 & x3;
  assign n1484 = (x4 & x8) | (x4 & n1483) | (x8 & n1483);
  assign n1485 = ~x8 & n1484;
  assign n1487 = x2 & n1485;
  assign n1488 = (n1482 & n1486) | (n1482 & n1487) | (n1486 & n1487);
  assign n1489 = (~x3 & x4) | (~x3 & x8) | (x4 & x8);
  assign n1490 = (x3 & x7) | (x3 & n1489) | (x7 & n1489);
  assign n1491 = (x4 & x8) | (x4 & n1490) | (x8 & n1490);
  assign n1492 = n1489 & ~n1491;
  assign n1493 = (n1490 & ~n1491) | (n1490 & n1492) | (~n1491 & n1492);
  assign n1499 = (x1 & ~x2) | (x1 & n1493) | (~x2 & n1493);
  assign n1494 = (x3 & x4) | (x3 & x8) | (x4 & x8);
  assign n1495 = (x4 & ~x7) | (x4 & n1494) | (~x7 & n1494);
  assign n1496 = x4 & ~n1495;
  assign n1497 = n1495 | n1496;
  assign n1498 = (~x4 & n1496) | (~x4 & n1497) | (n1496 & n1497);
  assign n1500 = (x1 & x2) | (x1 & ~n1498) | (x2 & ~n1498);
  assign n1501 = n1499 & ~n1500;
  assign n1502 = (x3 & ~x7) | (x3 & n39) | (~x7 & n39);
  assign n1503 = (x1 & x3) | (x1 & ~n39) | (x3 & ~n39);
  assign n1504 = (x2 & ~x7) | (x2 & n1503) | (~x7 & n1503);
  assign n1505 = ~n1502 & n1504;
  assign n1509 = (x0 & n811) | (x0 & n1505) | (n811 & n1505);
  assign n1506 = ~x3 & x7;
  assign n1507 = (x2 & n44) | (x2 & n1506) | (n44 & n1506);
  assign n1508 = ~x2 & n1507;
  assign n1510 = ~n811 & n1508;
  assign n1511 = (n1505 & ~n1509) | (n1505 & n1510) | (~n1509 & n1510);
  assign n1512 = (~n1488 & n1501) | (~n1488 & n1511) | (n1501 & n1511);
  assign n1513 = x0 & ~n1511;
  assign n1514 = (n1488 & n1512) | (n1488 & ~n1513) | (n1512 & ~n1513);
  assign n1664 = n1514 | n1663;
  assign n1665 = (~n1442 & n1663) | (~n1442 & n1664) | (n1663 & n1664);
  assign n1687 = (n36 & ~n118) | (n36 & n784) | (~n118 & n784);
  assign n1688 = (~x3 & n36) | (~x3 & n1687) | (n36 & n1687);
  assign n1689 = x1 & ~n1688;
  assign n1690 = ~x0 & n1689;
  assign n1691 = n399 & ~n1690;
  assign n1692 = (n318 & n1690) | (n318 & ~n1691) | (n1690 & ~n1691);
  assign n1666 = n318 & n591;
  assign n1667 = n20 & n1666;
  assign n1676 = x5 | n79;
  assign n1677 = (~n765 & n887) | (~n765 & n1676) | (n887 & n1676);
  assign n1678 = (n16 & n377) | (n16 & ~n851) | (n377 & ~n851);
  assign n1679 = (x1 & ~x2) | (x1 & n1678) | (~x2 & n1678);
  assign n1680 = ~x1 & n1679;
  assign n1681 = (x2 & n1679) | (x2 & n1680) | (n1679 & n1680);
  assign n1682 = x6 | n1681;
  assign n1683 = (n1677 & n1681) | (n1677 & n1682) | (n1681 & n1682);
  assign n1684 = (~x0 & x3) | (~x0 & n1683) | (x3 & n1683);
  assign n1670 = (x1 & x4) | (x1 & ~n15) | (x4 & ~n15);
  assign n1671 = (x4 & x5) | (x4 & ~n15) | (x5 & ~n15);
  assign n1672 = (n573 & n1670) | (n573 & ~n1671) | (n1670 & ~n1671);
  assign n1673 = ~x6 & n1672;
  assign n1668 = (x1 & ~x2) | (x1 & x6) | (~x2 & x6);
  assign n1669 = n930 & n1668;
  assign n1674 = n1669 | n1673;
  assign n1675 = (~x4 & n1673) | (~x4 & n1674) | (n1673 & n1674);
  assign n1685 = (x0 & x3) | (x0 & ~n1675) | (x3 & ~n1675);
  assign n1686 = n1684 & ~n1685;
  assign n1693 = (~n29 & n1667) | (~n29 & n1686) | (n1667 & n1686);
  assign n1694 = ~n1692 & n1693;
  assign n1695 = (~n29 & n1692) | (~n29 & n1694) | (n1692 & n1694);
  assign n1806 = (x0 & x3) | (x0 & n712) | (x3 & n712);
  assign n1807 = (x0 & x3) | (x0 & ~n712) | (x3 & ~n712);
  assign n1808 = (x4 & ~x8) | (x4 & n1807) | (~x8 & n1807);
  assign n1809 = ~n1806 & n1808;
  assign n1810 = ~x3 & n184;
  assign n1811 = (x0 & ~x4) | (x0 & n1810) | (~x4 & n1810);
  assign n1812 = ~x0 & n1811;
  assign n1813 = x7 | n1812;
  assign n1814 = (n1809 & n1812) | (n1809 & n1813) | (n1812 & n1813);
  assign n1815 = x1 | n1814;
  assign n1803 = x3 & x7;
  assign n1804 = x3 & ~n88;
  assign n1805 = (n86 & n1803) | (n86 & ~n1804) | (n1803 & ~n1804);
  assign n1816 = ~x0 & n1805;
  assign n1817 = x1 & ~n1816;
  assign n1818 = n1815 & ~n1817;
  assign n1819 = x2 | n1818;
  assign n1796 = (x1 & ~x4) | (x1 & n60) | (~x4 & n60);
  assign n1797 = (x4 & ~x7) | (x4 & n60) | (~x7 & n60);
  assign n1798 = (x1 & x8) | (x1 & ~n1797) | (x8 & ~n1797);
  assign n1799 = ~n1796 & n1798;
  assign n1800 = (~x4 & n184) | (~x4 & n1799) | (n184 & n1799);
  assign n1801 = n121 & ~n1800;
  assign n1802 = (n121 & n1799) | (n121 & ~n1801) | (n1799 & ~n1801);
  assign n1820 = ~x0 & n1802;
  assign n1821 = x2 & ~n1820;
  assign n1822 = n1819 & ~n1821;
  assign n1823 = x5 | n1822;
  assign n1784 = (n10 & n299) | (n10 & ~n1506) | (n299 & ~n1506);
  assign n1786 = x2 & ~n39;
  assign n1787 = n1784 & n1786;
  assign n1785 = ~x3 & n10;
  assign n1788 = (~n39 & n1785) | (~n39 & n1786) | (n1785 & n1786);
  assign n1789 = (x1 & n1787) | (x1 & n1788) | (n1787 & n1788);
  assign n1791 = n1785 & n1786;
  assign n1790 = x3 & n184;
  assign n1792 = (~n39 & n1786) | (~n39 & n1790) | (n1786 & n1790);
  assign n1793 = (x1 & n1791) | (x1 & n1792) | (n1791 & n1792);
  assign n1794 = x4 & ~n1793;
  assign n1795 = (n1789 & n1793) | (n1789 & ~n1794) | (n1793 & ~n1794);
  assign n1824 = ~x0 & n1795;
  assign n1825 = x5 & ~n1824;
  assign n1826 = n1823 & ~n1825;
  assign n1736 = ~n28 & n463;
  assign n1759 = (x4 & ~x7) | (x4 & n690) | (~x7 & n690);
  assign n1760 = x4 & ~n1759;
  assign n1761 = n1759 | n1760;
  assign n1762 = (~x4 & n1760) | (~x4 & n1761) | (n1760 & n1761);
  assign n1766 = ~x1 & n1762;
  assign n1767 = ~x1 & x7;
  assign n1763 = (~x2 & x4) | (~x2 & x8) | (x4 & x8);
  assign n1764 = x2 & n1763;
  assign n1765 = (~n153 & n1763) | (~n153 & n1764) | (n1763 & n1764);
  assign n1768 = (~x1 & x7) | (~x1 & n1765) | (x7 & n1765);
  assign n1769 = (n1766 & ~n1767) | (n1766 & n1768) | (~n1767 & n1768);
  assign n1770 = x3 & n1769;
  assign n1750 = (x1 & ~x4) | (x1 & x7) | (~x4 & x7);
  assign n1751 = (x4 & ~x8) | (x4 & n1750) | (~x8 & n1750);
  assign n1752 = (x1 & x7) | (x1 & n1751) | (x7 & n1751);
  assign n1753 = n1750 & ~n1752;
  assign n1754 = (n1751 & ~n1752) | (n1751 & n1753) | (~n1752 & n1753);
  assign n1755 = x2 & ~n1754;
  assign n1756 = x1 & n184;
  assign n1757 = x2 | n1756;
  assign n1758 = ~n1755 & n1757;
  assign n1771 = x3 | n1758;
  assign n1772 = (~x3 & n1770) | (~x3 & n1771) | (n1770 & n1771);
  assign n1773 = x6 & n1772;
  assign n1737 = x2 & n1571;
  assign n1738 = x3 | n1571;
  assign n1739 = (x2 & ~x4) | (x2 & n1738) | (~x4 & n1738);
  assign n1740 = ~n1737 & n1739;
  assign n1745 = (x1 & ~x8) | (x1 & n1740) | (~x8 & n1740);
  assign n1741 = ~x7 & n42;
  assign n1742 = (x3 & x4) | (x3 & ~n42) | (x4 & ~n42);
  assign n1743 = (x7 & n164) | (x7 & ~n1742) | (n164 & ~n1742);
  assign n1744 = (x7 & n1741) | (x7 & ~n1743) | (n1741 & ~n1743);
  assign n1746 = (x1 & x8) | (x1 & ~n1744) | (x8 & ~n1744);
  assign n1747 = n1745 & ~n1746;
  assign n1748 = (x1 & ~n184) | (x1 & n865) | (~n184 & n865);
  assign n1749 = n184 & n1748;
  assign n1774 = n1747 | n1749;
  assign n1775 = ~x6 & n1774;
  assign n1776 = n1773 | n1775;
  assign n1777 = ~x0 & n1776;
  assign n1778 = n46 | n1777;
  assign n1779 = (n1736 & n1777) | (n1736 & n1778) | (n1777 & n1778);
  assign n1780 = x5 & ~n1779;
  assign n1696 = (x2 & ~x7) | (x2 & x8) | (~x7 & x8);
  assign n1697 = (~x2 & x4) | (~x2 & n1696) | (x4 & n1696);
  assign n1698 = (x4 & x8) | (x4 & ~n1696) | (x8 & ~n1696);
  assign n1699 = n1697 & ~n1698;
  assign n1702 = (x1 & x6) | (x1 & ~n1699) | (x6 & ~n1699);
  assign n1700 = x4 & n79;
  assign n1701 = n60 & n1700;
  assign n1703 = x6 & n1701;
  assign n1704 = (n1699 & n1702) | (n1699 & n1703) | (n1702 & n1703);
  assign n1729 = (x1 & x4) | (x1 & x6) | (x4 & x6);
  assign n1724 = (x2 & x7) | (x2 & x8) | (x7 & x8);
  assign n1725 = (~x3 & x8) | (~x3 & n1724) | (x8 & n1724);
  assign n1726 = x8 & ~n1725;
  assign n1727 = n1725 | n1726;
  assign n1728 = (~x8 & n1726) | (~x8 & n1727) | (n1726 & n1727);
  assign n1730 = x1 | x4;
  assign n1731 = (x6 & n1728) | (x6 & n1730) | (n1728 & n1730);
  assign n1732 = ~n1729 & n1731;
  assign n1733 = (~x3 & n1704) | (~x3 & n1732) | (n1704 & n1732);
  assign n1712 = ~x2 & x7;
  assign n1713 = (x2 & x6) | (x2 & n1712) | (x6 & n1712);
  assign n1714 = (x1 & x6) | (x1 & n1712) | (x6 & n1712);
  assign n1715 = (n487 & n1713) | (n487 & ~n1714) | (n1713 & ~n1714);
  assign n1716 = x8 & ~n1715;
  assign n1709 = ~x1 & x6;
  assign n1710 = x1 & n640;
  assign n1711 = (x1 & n1709) | (x1 & ~n1710) | (n1709 & ~n1710);
  assign n1717 = x2 & ~n1711;
  assign n1718 = x8 | n1717;
  assign n1719 = ~n1716 & n1718;
  assign n1720 = x4 & ~n1719;
  assign n1705 = (x6 & ~x8) | (x6 & n87) | (~x8 & n87);
  assign n1706 = (~x1 & x8) | (~x1 & n1705) | (x8 & n1705);
  assign n1707 = (x6 & x7) | (x6 & ~n1706) | (x7 & ~n1706);
  assign n1708 = ~n1705 & n1707;
  assign n1721 = x2 & n1708;
  assign n1722 = x4 | n1721;
  assign n1723 = ~n1720 & n1722;
  assign n1734 = (x3 & n1723) | (x3 & n1732) | (n1723 & n1732);
  assign n1735 = n1733 | n1734;
  assign n1781 = ~x0 & n1735;
  assign n1782 = x5 | n1781;
  assign n1783 = ~n1780 & n1782;
  assign n1827 = n42 & n118;
  assign n1828 = (x1 & n583) | (x1 & n1827) | (n583 & n1827);
  assign n1829 = ~x1 & n1828;
  assign n1830 = (x2 & x6) | (x2 & n86) | (x6 & n86);
  assign n1831 = ~x2 & n1830;
  assign n1845 = (x1 & ~x3) | (x1 & n1831) | (~x3 & n1831);
  assign n1832 = (x1 & x4) | (x1 & ~x5) | (x4 & ~x5);
  assign n1833 = (x1 & ~x7) | (x1 & n1832) | (~x7 & n1832);
  assign n1834 = x1 & ~n1833;
  assign n1835 = n1833 | n1834;
  assign n1836 = (~x1 & n1834) | (~x1 & n1835) | (n1834 & n1835);
  assign n1842 = (~x2 & x6) | (~x2 & n1836) | (x6 & n1836);
  assign n1837 = (~x4 & x5) | (~x4 & x7) | (x5 & x7);
  assign n1838 = ~x5 & n1837;
  assign n1839 = (x4 & n1837) | (x4 & n1838) | (n1837 & n1838);
  assign n1840 = ~x1 & n1839;
  assign n1841 = ~x2 & n1840;
  assign n1843 = ~x6 & n1841;
  assign n1844 = (n1836 & ~n1842) | (n1836 & n1843) | (~n1842 & n1843);
  assign n1846 = ~x3 & n1844;
  assign n1847 = (~x1 & n1845) | (~x1 & n1846) | (n1845 & n1846);
  assign n1848 = n46 & n552;
  assign n1849 = n16 & n1848;
  assign n1850 = (~n1829 & n1847) | (~n1829 & n1849) | (n1847 & n1849);
  assign n1851 = x0 & ~n1849;
  assign n1852 = (n1829 & n1850) | (n1829 & ~n1851) | (n1850 & ~n1851);
  assign n1853 = n1783 | n1852;
  assign n1854 = (~n1695 & n1826) | (~n1695 & n1853) | (n1826 & n1853);
  assign n1855 = n1695 | n1854;
  assign n1861 = x1 & ~x5;
  assign n1862 = (~x0 & x3) | (~x0 & n1861) | (x3 & n1861);
  assign n1863 = (x1 & x3) | (x1 & ~n1861) | (x3 & ~n1861);
  assign n1864 = (x5 & n1862) | (x5 & ~n1863) | (n1862 & ~n1863);
  assign n1865 = (x1 & ~x7) | (x1 & n120) | (~x7 & n120);
  assign n1866 = ~x1 & n1865;
  assign n1867 = x7 | n1866;
  assign n1868 = (n1864 & n1866) | (n1864 & n1867) | (n1866 & n1867);
  assign n1869 = x2 | n1868;
  assign n1857 = (~x1 & x5) | (~x1 & n1803) | (x5 & n1803);
  assign n1858 = (x1 & ~x3) | (x1 & n1803) | (~x3 & n1803);
  assign n1859 = (x5 & x7) | (x5 & ~n1858) | (x7 & ~n1858);
  assign n1860 = ~n1857 & n1859;
  assign n1870 = ~x0 & n1860;
  assign n1871 = x2 & ~n1870;
  assign n1872 = n1869 & ~n1871;
  assign n1856 = (n88 & ~n463) | (n88 & n684) | (~n463 & n684);
  assign n2043 = ~n1856 & n1872;
  assign n1918 = (x1 & x3) | (x1 & ~x7) | (x3 & ~x7);
  assign n1919 = n1050 & ~n1918;
  assign n1920 = x0 | n1919;
  assign n1917 = x4 | n1561;
  assign n1921 = x1 | n1917;
  assign n1922 = x0 & n1921;
  assign n1923 = n1920 & ~n1922;
  assign n1976 = n1222 & n1923;
  assign n1924 = n37 & n44;
  assign n1925 = (n20 & ~n184) | (n20 & n1924) | (~n184 & n1924);
  assign n1926 = n184 & n1925;
  assign n1927 = (~x3 & x7) | (~x3 & x8) | (x7 & x8);
  assign n1928 = (x3 & ~x8) | (x3 & n1927) | (~x8 & n1927);
  assign n1929 = ~x6 & n1927;
  assign n1930 = (~x7 & n1927) | (~x7 & n1929) | (n1927 & n1929);
  assign n1931 = n1928 | n1930;
  assign n1932 = x1 & n1931;
  assign n1933 = x3 | n77;
  assign n1934 = ~x1 & n1933;
  assign n1935 = n1932 | n1934;
  assign n1944 = x4 & ~n1935;
  assign n1936 = ~x1 & x8;
  assign n1937 = (x6 & n299) | (x6 & n1936) | (n299 & n1936);
  assign n1938 = (x3 & ~x6) | (x3 & n1937) | (~x6 & n1937);
  assign n1939 = (~x8 & n1936) | (~x8 & n1938) | (n1936 & n1938);
  assign n1940 = (~n1936 & n1937) | (~n1936 & n1939) | (n1937 & n1939);
  assign n1941 = ~n77 & n121;
  assign n1942 = x7 | n1941;
  assign n1943 = (n1940 & n1941) | (n1940 & n1942) | (n1941 & n1942);
  assign n1945 = x4 | n1943;
  assign n1946 = (~x4 & n1944) | (~x4 & n1945) | (n1944 & n1945);
  assign n1973 = (~x0 & x5) | (~x0 & n1946) | (x5 & n1946);
  assign n1955 = x7 & ~n811;
  assign n1956 = ~x6 & n1955;
  assign n1964 = ~x3 & n1956;
  assign n1957 = x6 & n20;
  assign n1958 = ~n28 & n1957;
  assign n1959 = (x3 & ~x4) | (x3 & x8) | (~x4 & x8);
  assign n1960 = (~x3 & x7) | (~x3 & n1959) | (x7 & n1959);
  assign n1961 = (~x4 & x8) | (~x4 & n1960) | (x8 & n1960);
  assign n1962 = ~n1959 & n1961;
  assign n1963 = (~n1960 & n1961) | (~n1960 & n1962) | (n1961 & n1962);
  assign n1965 = n1958 | n1963;
  assign n1966 = (n1956 & ~n1964) | (n1956 & n1965) | (~n1964 & n1965);
  assign n1967 = x1 | n1966;
  assign n1951 = x3 & ~x8;
  assign n1952 = (x3 & ~x7) | (x3 & n351) | (~x7 & n351);
  assign n1953 = n351 | n1952;
  assign n1954 = ~n1951 & n1953;
  assign n1968 = ~x6 & n1954;
  assign n1969 = x1 & ~n1968;
  assign n1970 = n1967 & ~n1969;
  assign n1947 = (x6 & ~x8) | (x6 & n1149) | (~x8 & n1149);
  assign n1948 = x8 & n1947;
  assign n1949 = n1947 & ~n1948;
  assign n1950 = (x8 & ~n1948) | (x8 & n1949) | (~n1948 & n1949);
  assign n1971 = (x3 & ~x4) | (x3 & n1950) | (~x4 & n1950);
  assign n1972 = (n20 & ~n1970) | (n20 & n1971) | (~n1970 & n1971);
  assign n1974 = (x0 & x5) | (x0 & n1972) | (x5 & n1972);
  assign n1975 = n1973 & ~n1974;
  assign n1977 = n1926 | n1975;
  assign n1978 = (n1923 & ~n1976) | (n1923 & n1977) | (~n1976 & n1977);
  assign n1979 = x2 | n1978;
  assign n1900 = (~x3 & x8) | (~x3 & n225) | (x8 & n225);
  assign n1901 = (x5 & x7) | (x5 & n1900) | (x7 & n1900);
  assign n1902 = ~n225 & n1901;
  assign n1903 = (~n1900 & n1901) | (~n1900 & n1902) | (n1901 & n1902);
  assign n1904 = x1 | n1903;
  assign n1905 = x3 | n185;
  assign n1906 = x1 & n1905;
  assign n1907 = n1904 & ~n1906;
  assign n1908 = x4 & n1907;
  assign n1891 = (~x3 & x5) | (~x3 & x7) | (x5 & x7);
  assign n1892 = (x1 & x5) | (x1 & ~n1891) | (x5 & ~n1891);
  assign n1893 = (~x5 & x7) | (~x5 & n1892) | (x7 & n1892);
  assign n1894 = n1891 & n1893;
  assign n1895 = x1 & ~n1894;
  assign n1896 = (n1892 & n1894) | (n1892 & ~n1895) | (n1894 & ~n1895);
  assign n1897 = x8 & n1896;
  assign n1888 = (x1 & ~x3) | (x1 & x7) | (~x3 & x7);
  assign n1889 = (~x1 & x3) | (~x1 & x8) | (x3 & x8);
  assign n1890 = n1888 | n1889;
  assign n1898 = n1890 & ~n1897;
  assign n1899 = (x5 & n1897) | (x5 & ~n1898) | (n1897 & ~n1898);
  assign n1909 = x4 | n1899;
  assign n1910 = (~x4 & n1908) | (~x4 & n1909) | (n1908 & n1909);
  assign n1911 = x6 & ~n1910;
  assign n1881 = x1 & x5;
  assign n1882 = x3 & x5;
  assign n1883 = (x1 & ~x7) | (x1 & n1882) | (~x7 & n1882);
  assign n1884 = (n755 & ~n1881) | (n755 & n1883) | (~n1881 & n1883);
  assign n1885 = x4 & n1884;
  assign n1886 = (x4 & ~x7) | (x4 & n1531) | (~x7 & n1531);
  assign n1887 = (~n86 & n1885) | (~n86 & n1886) | (n1885 & n1886);
  assign n1912 = x8 & n1887;
  assign n1913 = x6 | n1912;
  assign n1914 = ~n1911 & n1913;
  assign n1873 = (~x1 & x8) | (~x1 & n437) | (x8 & n437);
  assign n1874 = (x7 & x8) | (x7 & ~n437) | (x8 & ~n437);
  assign n1875 = (~x1 & x4) | (~x1 & n1874) | (x4 & n1874);
  assign n1876 = ~n1873 & n1875;
  assign n1877 = x5 & ~n1876;
  assign n1878 = n10 & ~n1730;
  assign n1879 = x5 | n1878;
  assign n1880 = ~n1877 & n1879;
  assign n1915 = (~x3 & x6) | (~x3 & n1880) | (x6 & n1880);
  assign n1916 = (~n1385 & n1914) | (~n1385 & n1915) | (n1914 & n1915);
  assign n1980 = ~x0 & n1916;
  assign n1981 = x2 & ~n1980;
  assign n1982 = n1979 & ~n1981;
  assign n2022 = (~x3 & x4) | (~x3 & x7) | (x4 & x7);
  assign n2023 = (x1 & x3) | (x1 & n2022) | (x3 & n2022);
  assign n2024 = (x3 & x7) | (x3 & ~n2023) | (x7 & ~n2023);
  assign n2025 = n2022 & n2024;
  assign n2026 = (x1 & ~n2023) | (x1 & n2025) | (~n2023 & n2025);
  assign n2027 = x2 & ~n2026;
  assign n2020 = x3 & ~n350;
  assign n2021 = (x4 & ~n350) | (x4 & n2020) | (~n350 & n2020);
  assign n2028 = x1 & n2021;
  assign n2029 = x2 | n2028;
  assign n2030 = ~n2027 & n2029;
  assign n2031 = x6 & ~n2030;
  assign n2016 = (x1 & x3) | (x1 & ~n1336) | (x3 & ~n1336);
  assign n2017 = (x2 & x4) | (x2 & ~n2016) | (x4 & ~n2016);
  assign n2018 = ~n1336 & n2017;
  assign n2019 = (n2016 & n2017) | (n2016 & n2018) | (n2017 & n2018);
  assign n2032 = ~x7 & n2019;
  assign n2033 = x6 | n2032;
  assign n2034 = ~n2031 & n2033;
  assign n2035 = x0 | n2034;
  assign n2015 = n20 & ~n564;
  assign n2036 = ~n15 & n2015;
  assign n2037 = x0 & ~n2036;
  assign n2038 = n2035 & ~n2037;
  assign n2039 = x5 & n2038;
  assign n1983 = (x2 & ~x3) | (x2 & x6) | (~x3 & x6);
  assign n1984 = x6 & ~n1983;
  assign n1985 = (x1 & x2) | (x1 & n1984) | (x2 & n1984);
  assign n1986 = (~n1983 & n1984) | (~n1983 & n1985) | (n1984 & n1985);
  assign n1989 = (x0 & ~n215) | (x0 & n1986) | (~n215 & n1986);
  assign n1987 = (x2 & n44) | (x2 & n1385) | (n44 & n1385);
  assign n1988 = ~x2 & n1987;
  assign n1990 = ~n215 & n1988;
  assign n1991 = (~x0 & n1989) | (~x0 & n1990) | (n1989 & n1990);
  assign n1992 = ~x6 & n20;
  assign n2012 = n318 & ~n1992;
  assign n1993 = (x4 & n40) | (x4 & n1437) | (n40 & n1437);
  assign n1994 = ~x4 & n1993;
  assign n2002 = (x1 & x7) | (x1 & ~n1437) | (x7 & ~n1437);
  assign n2003 = (~x1 & x3) | (~x1 & n2002) | (x3 & n2002);
  assign n2004 = (x6 & ~x7) | (x6 & n2003) | (~x7 & n2003);
  assign n2005 = n2002 & n2004;
  assign n2006 = ~x1 & n1122;
  assign n2007 = x4 & ~n2006;
  assign n2008 = (n2005 & n2006) | (n2005 & ~n2007) | (n2006 & ~n2007);
  assign n2009 = (~x0 & x2) | (~x0 & n2008) | (x2 & n2008);
  assign n1995 = (x1 & x7) | (x1 & ~n1561) | (x7 & ~n1561);
  assign n1996 = (x1 & x6) | (x1 & ~n1561) | (x6 & ~n1561);
  assign n1997 = (n640 & n1995) | (n640 & ~n1996) | (n1995 & ~n1996);
  assign n1998 = x4 | n1997;
  assign n1999 = n121 & n552;
  assign n2000 = x4 & ~n1999;
  assign n2001 = n1998 & ~n2000;
  assign n2010 = (x0 & x2) | (x0 & ~n2001) | (x2 & ~n2001);
  assign n2011 = n2009 & ~n2010;
  assign n2013 = n1994 | n2011;
  assign n2014 = (n318 & ~n2012) | (n318 & n2013) | (~n2012 & n2013);
  assign n2040 = n1991 | n2014;
  assign n2041 = ~x5 & n2040;
  assign n2042 = n2039 | n2041;
  assign n2044 = n1982 | n2042;
  assign n2045 = (n1872 & ~n2043) | (n1872 & n2044) | (~n2043 & n2044);
  assign n2046 = (x3 & ~x5) | (x3 & x6) | (~x5 & x6);
  assign n2047 = (x4 & ~x6) | (x4 & n2046) | (~x6 & n2046);
  assign n2048 = (x3 & x4) | (x3 & ~n2046) | (x4 & ~n2046);
  assign n2049 = n2047 & ~n2048;
  assign n2051 = (x0 & ~x1) | (x0 & n2049) | (~x1 & n2049);
  assign n2050 = n1098 & ~n1354;
  assign n2052 = ~x0 & n2050;
  assign n2053 = (n2049 & ~n2051) | (n2049 & n2052) | (~n2051 & n2052);
  assign n2054 = (x3 & x5) | (x3 & x6) | (x5 & x6);
  assign n2055 = (~x4 & x6) | (~x4 & n2054) | (x6 & n2054);
  assign n2056 = x6 & ~n2055;
  assign n2057 = n2055 | n2056;
  assign n2058 = (~x6 & n2056) | (~x6 & n2057) | (n2056 & n2057);
  assign n2059 = (x1 & n1104) | (x1 & ~n2058) | (n1104 & ~n2058);
  assign n2060 = n2058 & n2059;
  assign n2061 = (n1357 & ~n2053) | (n1357 & n2060) | (~n2053 & n2060);
  assign n2062 = x2 & ~n2060;
  assign n2063 = (n2053 & n2061) | (n2053 & ~n2062) | (n2061 & ~n2062);
  assign n2209 = ~n29 & n2063;
  assign n2086 = (x5 & x8) | (x5 & ~n400) | (x8 & ~n400);
  assign n2087 = (~x0 & x5) | (~x0 & n400) | (x5 & n400);
  assign n2088 = (~x2 & x8) | (~x2 & n2087) | (x8 & n2087);
  assign n2089 = n2086 & ~n2088;
  assign n2090 = ~x7 & n2089;
  assign n2085 = (~x5 & n634) | (~x5 & n1712) | (n634 & n1712);
  assign n2091 = n2085 | n2090;
  assign n2092 = (x0 & n2090) | (x0 & n2091) | (n2090 & n2091);
  assign n2093 = x4 & ~n2092;
  assign n2082 = ~x7 & n1185;
  assign n2083 = (x2 & x5) | (x2 & ~n2082) | (x5 & ~n2082);
  assign n2084 = (n1185 & n2082) | (n1185 & ~n2083) | (n2082 & ~n2083);
  assign n2094 = ~x0 & n2084;
  assign n2095 = x4 | n2094;
  assign n2096 = ~n2093 & n2095;
  assign n2110 = x1 & n2096;
  assign n2097 = (n129 & n184) | (n129 & n763) | (n184 & n763);
  assign n2098 = (~x8 & n184) | (~x8 & n2097) | (n184 & n2097);
  assign n2099 = (x4 & ~n43) | (x4 & n2098) | (~n43 & n2098);
  assign n2100 = n2098 & ~n2099;
  assign n2101 = (x1 & n811) | (x1 & n813) | (n811 & n813);
  assign n2102 = ~n811 & n2101;
  assign n2103 = (~x4 & n717) | (~x4 & n2102) | (n717 & n2102);
  assign n2104 = n79 & ~n2103;
  assign n2105 = (n79 & n2102) | (n79 & ~n2104) | (n2102 & ~n2104);
  assign n2106 = x0 | n2105;
  assign n2107 = n15 | n1596;
  assign n2108 = x0 & n2107;
  assign n2109 = n2106 & ~n2108;
  assign n2111 = n2100 | n2109;
  assign n2112 = (n2096 & ~n2110) | (n2096 & n2111) | (~n2110 & n2111);
  assign n2113 = x3 | n2112;
  assign n2064 = (x5 & ~x7) | (x5 & n178) | (~x7 & n178);
  assign n2065 = (x7 & x8) | (x7 & ~n178) | (x8 & ~n178);
  assign n2066 = (~n54 & n2064) | (~n54 & n2065) | (n2064 & n2065);
  assign n2067 = x4 & ~n2066;
  assign n2068 = x2 & n60;
  assign n2069 = x4 | n2068;
  assign n2070 = ~n2067 & n2069;
  assign n2079 = x1 & n2070;
  assign n2071 = (x5 & n311) | (x5 & ~n1712) | (n311 & ~n1712);
  assign n2072 = (~x5 & x7) | (~x5 & n2071) | (x7 & n2071);
  assign n2073 = (~x2 & n311) | (~x2 & n2072) | (n311 & n2072);
  assign n2074 = (~n311 & n2071) | (~n311 & n2073) | (n2071 & n2073);
  assign n2075 = ~x4 & n2074;
  assign n2076 = ~x2 & n213;
  assign n2077 = x4 & ~n2076;
  assign n2078 = n2075 | n2077;
  assign n2080 = ~x1 & n2078;
  assign n2081 = (x1 & ~n2079) | (x1 & n2080) | (~n2079 & n2080);
  assign n2114 = x0 | n2081;
  assign n2115 = x3 & n2114;
  assign n2116 = n2113 & ~n2115;
  assign n2161 = (x2 & ~x3) | (x2 & n1061) | (~x3 & n1061);
  assign n2162 = x2 | n2161;
  assign n2163 = x2 & n2161;
  assign n2164 = n2162 & ~n2163;
  assign n2166 = (x0 & ~x7) | (x0 & n2164) | (~x7 & n2164);
  assign n2165 = ~n15 & n1122;
  assign n2167 = ~x0 & n2165;
  assign n2168 = (n2164 & ~n2166) | (n2164 & n2167) | (~n2166 & n2167);
  assign n2169 = (x3 & n318) | (x3 & n790) | (n318 & n790);
  assign n2170 = ~x3 & n2169;
  assign n2196 = n183 & ~n860;
  assign n2183 = (x5 & x7) | (x5 & n1127) | (x7 & n1127);
  assign n2184 = (x4 & x7) | (x4 & ~n2183) | (x7 & ~n2183);
  assign n2185 = n1127 | n2184;
  assign n2186 = (x5 & ~n2183) | (x5 & n2185) | (~n2183 & n2185);
  assign n2187 = x6 & ~n2186;
  assign n2188 = ~x2 & n2187;
  assign n2189 = (x2 & ~x7) | (x2 & n1448) | (~x7 & n1448);
  assign n2190 = x2 & ~n2189;
  assign n2191 = n2189 | n2190;
  assign n2192 = (~x2 & n2190) | (~x2 & n2191) | (n2190 & n2191);
  assign n2193 = ~x2 & n1992;
  assign n2194 = x6 | n2193;
  assign n2195 = (n2192 & n2193) | (n2192 & n2194) | (n2193 & n2194);
  assign n2197 = n2188 | n2195;
  assign n2198 = (n183 & ~n2196) | (n183 & n2197) | (~n2196 & n2197);
  assign n2199 = (~x0 & x1) | (~x0 & n2198) | (x1 & n2198);
  assign n2171 = (~x3 & x6) | (~x3 & x7) | (x6 & x7);
  assign n2172 = x7 & n2171;
  assign n2173 = (~x3 & x4) | (~x3 & n2172) | (x4 & n2172);
  assign n2174 = (n377 & n2171) | (n377 & ~n2173) | (n2171 & ~n2173);
  assign n2175 = x5 | n2174;
  assign n2176 = n80 & ~n564;
  assign n2177 = x5 & ~n2176;
  assign n2178 = n2175 & ~n2177;
  assign n2179 = x2 | n2178;
  assign n2180 = n20 & n553;
  assign n2181 = x2 & ~n2180;
  assign n2182 = n2179 & ~n2181;
  assign n2200 = (x0 & x1) | (x0 & ~n2182) | (x1 & ~n2182);
  assign n2201 = n2199 & ~n2200;
  assign n2202 = (~n2168 & n2170) | (~n2168 & n2201) | (n2170 & n2201);
  assign n2203 = n1442 & ~n2201;
  assign n2204 = (n2168 & n2202) | (n2168 & ~n2203) | (n2202 & ~n2203);
  assign n2205 = x8 & ~n2204;
  assign n2117 = x3 | n797;
  assign n2118 = x3 & n798;
  assign n2119 = n2117 & ~n2118;
  assign n2120 = x4 & ~n2119;
  assign n2121 = x3 & n129;
  assign n2122 = x4 | n2121;
  assign n2123 = ~n2120 & n2122;
  assign n2124 = ~x5 & n183;
  assign n2125 = n583 & n2124;
  assign n2126 = x6 & ~n2125;
  assign n2127 = (n2123 & n2125) | (n2123 & ~n2126) | (n2125 & ~n2126);
  assign n2149 = (x3 & x4) | (x3 & ~x5) | (x4 & ~x5);
  assign n2150 = (x3 & ~x7) | (x3 & n2149) | (~x7 & n2149);
  assign n2151 = x3 & ~n2150;
  assign n2152 = n2150 | n2151;
  assign n2153 = (~x3 & n2151) | (~x3 & n2152) | (n2151 & n2152);
  assign n2154 = (x2 & x6) | (x2 & n2153) | (x6 & n2153);
  assign n2155 = (x1 & ~x6) | (x1 & n2154) | (~x6 & n2154);
  assign n2156 = (x1 & x2) | (x1 & ~n2154) | (x2 & ~n2154);
  assign n2157 = n2155 & ~n2156;
  assign n2158 = (~x1 & n2127) | (~x1 & n2157) | (n2127 & n2157);
  assign n2131 = x3 & ~x6;
  assign n2132 = (~x4 & x7) | (~x4 & n2131) | (x7 & n2131);
  assign n2133 = (x6 & ~x7) | (x6 & n2131) | (~x7 & n2131);
  assign n2134 = (~x3 & x4) | (~x3 & n2133) | (x4 & n2133);
  assign n2135 = n2132 | n2134;
  assign n2142 = x2 | n2135;
  assign n2136 = n416 & n552;
  assign n2137 = (x2 & x3) | (x2 & ~x6) | (x3 & ~x6);
  assign n2138 = (x2 & ~x7) | (x2 & n2137) | (~x7 & n2137);
  assign n2139 = x2 & ~n2138;
  assign n2140 = n2138 | n2139;
  assign n2141 = (~x2 & n2139) | (~x2 & n2140) | (n2139 & n2140);
  assign n2143 = n2136 | n2141;
  assign n2144 = (~n2135 & n2142) | (~n2135 & n2143) | (n2142 & n2143);
  assign n2145 = x5 & ~n2144;
  assign n2128 = (x7 & n73) | (x7 & ~n2022) | (n73 & ~n2022);
  assign n2129 = (~x2 & n2022) | (~x2 & n2128) | (n2022 & n2128);
  assign n2130 = (~x7 & n2128) | (~x7 & n2129) | (n2128 & n2129);
  assign n2146 = x6 | n2130;
  assign n2147 = ~x5 & n2146;
  assign n2148 = n2145 | n2147;
  assign n2159 = (x1 & ~n2148) | (x1 & n2157) | (~n2148 & n2157);
  assign n2160 = n2158 | n2159;
  assign n2206 = ~x0 & n2160;
  assign n2207 = x8 | n2206;
  assign n2208 = ~n2205 & n2207;
  assign n2210 = n2116 | n2208;
  assign n2211 = (n2063 & ~n2209) | (n2063 & n2210) | (~n2209 & n2210);
  assign n2212 = x0 & x3;
  assign n2213 = (~x4 & x5) | (~x4 & n2212) | (x5 & n2212);
  assign n2214 = (x3 & x5) | (x3 & ~n2212) | (x5 & ~n2212);
  assign n2215 = (x0 & ~x4) | (x0 & n2214) | (~x4 & n2214);
  assign n2216 = ~n2213 & n2215;
  assign n2219 = (x1 & x2) | (x1 & n2216) | (x2 & n2216);
  assign n2217 = (x4 & n43) | (x4 & n618) | (n43 & n618);
  assign n2218 = ~x4 & n2217;
  assign n2220 = ~x2 & n2218;
  assign n2221 = (n2216 & ~n2219) | (n2216 & n2220) | (~n2219 & n2220);
  assign n2222 = (~x3 & n61) | (~x3 & n2221) | (n61 & n2221);
  assign n2223 = n40 & ~n2222;
  assign n2224 = (n40 & n2221) | (n40 & ~n2223) | (n2221 & ~n2223);
  assign n2407 = n738 & n2224;
  assign n2303 = (~n573 & n655) | (~n573 & n1936) | (n655 & n1936);
  assign n2304 = (x3 & ~x7) | (x3 & n2303) | (~x7 & n2303);
  assign n2305 = ~x3 & n2304;
  assign n2306 = (x7 & n2304) | (x7 & n2305) | (n2304 & n2305);
  assign n2307 = n1354 & ~n2306;
  assign n2308 = (n271 & n2306) | (n271 & ~n2307) | (n2306 & ~n2307);
  assign n2309 = x6 & ~n2308;
  assign n2310 = x5 & ~n1890;
  assign n2311 = x6 | n2310;
  assign n2312 = ~n2309 & n2311;
  assign n2313 = ~x2 & n2312;
  assign n2292 = (x5 & ~x6) | (x5 & x8) | (~x6 & x8);
  assign n2293 = (x7 & x8) | (x7 & ~n2292) | (x8 & ~n2292);
  assign n2294 = (~x5 & x7) | (~x5 & n2292) | (x7 & n2292);
  assign n2295 = n2293 & ~n2294;
  assign n2298 = (~x1 & x3) | (~x1 & n2295) | (x3 & n2295);
  assign n2296 = x5 & n29;
  assign n2297 = ~x6 & n2296;
  assign n2299 = (x1 & x3) | (x1 & n2297) | (x3 & n2297);
  assign n2300 = n2298 & n2299;
  assign n2301 = ~x1 & n882;
  assign n2302 = n53 & n2301;
  assign n2314 = n2300 | n2302;
  assign n2315 = x2 & n2314;
  assign n2316 = n2313 | n2315;
  assign n2277 = (x2 & ~x6) | (x2 & n847) | (~x6 & n847);
  assign n2278 = x2 & ~n2277;
  assign n2279 = n2277 | n2278;
  assign n2280 = (~x2 & n2278) | (~x2 & n2279) | (n2278 & n2279);
  assign n2283 = (x1 & n29) | (x1 & n2280) | (n29 & n2280);
  assign n2281 = ~x3 & n39;
  assign n2282 = n591 & n2281;
  assign n2284 = ~n29 & n2282;
  assign n2285 = (n2280 & ~n2283) | (n2280 & n2284) | (~n2283 & n2284);
  assign n2286 = ~x5 & n79;
  assign n2287 = x6 & ~n28;
  assign n2288 = n2286 & n2287;
  assign n2289 = (x1 & ~x2) | (x1 & n2288) | (~x2 & n2288);
  assign n2290 = n882 & ~n2289;
  assign n2291 = (n882 & n2288) | (n882 & ~n2290) | (n2288 & ~n2290);
  assign n2317 = (~x0 & n2285) | (~x0 & n2291) | (n2285 & n2291);
  assign n2318 = ~n2316 & n2317;
  assign n2319 = (~x0 & n2316) | (~x0 & n2318) | (n2316 & n2318);
  assign n2320 = (n46 & n184) | (n46 & n2319) | (n184 & n2319);
  assign n2321 = n37 & ~n2320;
  assign n2322 = (n37 & n2319) | (n37 & ~n2321) | (n2319 & ~n2321);
  assign n2329 = (x5 & ~x7) | (x5 & n171) | (~x7 & n171);
  assign n2330 = x7 & n2329;
  assign n2331 = n2329 & ~n2330;
  assign n2332 = (x7 & ~n2330) | (x7 & n2331) | (~n2330 & n2331);
  assign n2333 = x4 & ~n2332;
  assign n2334 = x2 & n2333;
  assign n2335 = n860 | n2334;
  assign n2336 = (~n624 & n2334) | (~n624 & n2335) | (n2334 & n2335);
  assign n2337 = (~x0 & x1) | (~x0 & n2336) | (x1 & n2336);
  assign n2323 = (x5 & x7) | (x5 & ~n1302) | (x7 & ~n1302);
  assign n2324 = (x4 & ~x6) | (x4 & n2323) | (~x6 & n2323);
  assign n2325 = n1302 | n2324;
  assign n2326 = (~n2323 & n2324) | (~n2323 & n2325) | (n2324 & n2325);
  assign n2327 = x3 | n2326;
  assign n2328 = x2 | n2327;
  assign n2338 = (x0 & x1) | (x0 & n2328) | (x1 & n2328);
  assign n2339 = n2337 & ~n2338;
  assign n2340 = (n16 & n46) | (n16 & n2339) | (n46 & n2339);
  assign n2341 = n564 | n2340;
  assign n2342 = (~n564 & n2339) | (~n564 & n2341) | (n2339 & n2341);
  assign n2343 = (x4 & n2322) | (x4 & n2342) | (n2322 & n2342);
  assign n2255 = (x6 & ~x8) | (x6 & n1927) | (~x8 & n1927);
  assign n2256 = (~x7 & x8) | (~x7 & n2255) | (x8 & n2255);
  assign n2257 = ~n1927 & n2256;
  assign n2258 = (~x6 & n2255) | (~x6 & n2257) | (n2255 & n2257);
  assign n2259 = x1 | n2258;
  assign n2260 = ~x3 & n257;
  assign n2261 = x1 & ~n2260;
  assign n2262 = n2259 & ~n2261;
  assign n2263 = (x7 & x8) | (x7 & n122) | (x8 & n122);
  assign n2264 = (x6 & ~x7) | (x6 & n2263) | (~x7 & n2263);
  assign n2265 = (x6 & x8) | (x6 & ~n2263) | (x8 & ~n2263);
  assign n2266 = n2264 & ~n2265;
  assign n2267 = x0 & ~n2266;
  assign n2268 = (n2262 & n2266) | (n2262 & ~n2267) | (n2266 & ~n2267);
  assign n2269 = x2 | n2268;
  assign n2252 = ~n96 & n571;
  assign n2242 = x3 | x8;
  assign n2243 = (~x1 & x3) | (~x1 & n1385) | (x3 & n1385);
  assign n2244 = (x1 & x8) | (x1 & ~n1385) | (x8 & ~n1385);
  assign n2245 = (~n2242 & n2243) | (~n2242 & n2244) | (n2243 & n2244);
  assign n2246 = ~x7 & n2245;
  assign n2247 = (~x6 & n564) | (~x6 & n640) | (n564 & n640);
  assign n2248 = (x3 & x8) | (x3 & ~n2247) | (x8 & ~n2247);
  assign n2249 = (x1 & ~x3) | (x1 & n2248) | (~x3 & n2248);
  assign n2250 = (x1 & x8) | (x1 & ~n2248) | (x8 & ~n2248);
  assign n2251 = n2249 & ~n2250;
  assign n2253 = n2246 | n2251;
  assign n2254 = (n571 & ~n2252) | (n571 & n2253) | (~n2252 & n2253);
  assign n2270 = ~x0 & n2254;
  assign n2271 = x2 & ~n2270;
  assign n2272 = n2269 & ~n2271;
  assign n2273 = x5 | n2272;
  assign n2231 = (x8 & n552) | (x8 & n1803) | (n552 & n1803);
  assign n2232 = (x3 & x8) | (x3 & ~n2231) | (x8 & ~n2231);
  assign n2233 = (x7 & ~n552) | (x7 & n2232) | (~n552 & n2232);
  assign n2234 = (n552 & ~n2231) | (n552 & n2233) | (~n2231 & n2233);
  assign n2235 = x1 & ~n2234;
  assign n2227 = x7 & n172;
  assign n2228 = x6 | n172;
  assign n2229 = (x7 & x8) | (x7 & n2228) | (x8 & n2228);
  assign n2230 = ~n2227 & n2229;
  assign n2236 = x1 | n2230;
  assign n2237 = (~x1 & n2235) | (~x1 & n2236) | (n2235 & n2236);
  assign n2238 = x2 & ~n2237;
  assign n2225 = x6 & ~n29;
  assign n2226 = (x3 & ~n29) | (x3 & n2225) | (~n29 & n2225);
  assign n2239 = ~x1 & n2226;
  assign n2240 = x2 | n2239;
  assign n2241 = ~n2238 & n2240;
  assign n2274 = ~x0 & n2241;
  assign n2275 = x5 & ~n2274;
  assign n2276 = n2273 & ~n2275;
  assign n2344 = (~x4 & n2276) | (~x4 & n2342) | (n2276 & n2342);
  assign n2345 = n2343 | n2344;
  assign n2374 = x2 & x6;
  assign n2375 = (x4 & x8) | (x4 & n2374) | (x8 & n2374);
  assign n2376 = x4 | n2375;
  assign n2377 = x4 & n2375;
  assign n2378 = n2376 & ~n2377;
  assign n2379 = x5 | n2378;
  assign n2372 = x8 & n476;
  assign n2373 = (x8 & n712) | (x8 & ~n2372) | (n712 & ~n2372);
  assign n2380 = x2 | n2373;
  assign n2381 = x5 & n2380;
  assign n2382 = n2379 & ~n2381;
  assign n2383 = x1 & ~n2382;
  assign n2368 = (x2 & x4) | (x2 & ~n591) | (x4 & ~n591);
  assign n2369 = (x2 & ~x6) | (x2 & n591) | (~x6 & n591);
  assign n2370 = (x4 & ~x5) | (x4 & n2369) | (~x5 & n2369);
  assign n2371 = n2368 & ~n2370;
  assign n2384 = ~x8 & n2371;
  assign n2385 = x1 | n2384;
  assign n2386 = ~n2383 & n2385;
  assign n2387 = x3 & n2386;
  assign n2346 = (x4 & x5) | (x4 & x8) | (x5 & x8);
  assign n2347 = (~x6 & x8) | (~x6 & n2346) | (x8 & n2346);
  assign n2348 = x8 & ~n2347;
  assign n2349 = n2347 | n2348;
  assign n2350 = (~x8 & n2348) | (~x8 & n2349) | (n2348 & n2349);
  assign n2351 = x1 & ~n2350;
  assign n2352 = ~x4 & n717;
  assign n2353 = x1 | n2352;
  assign n2354 = ~n2351 & n2353;
  assign n2355 = ~x6 & n717;
  assign n2356 = x1 & n519;
  assign n2357 = n2355 & n2356;
  assign n2358 = x2 & ~n2357;
  assign n2359 = (n2354 & n2357) | (n2354 & ~n2358) | (n2357 & ~n2358);
  assign n2360 = (x2 & x4) | (x2 & ~x8) | (x4 & ~x8);
  assign n2361 = (~x4 & x6) | (~x4 & n2360) | (x6 & n2360);
  assign n2362 = (x2 & x6) | (x2 & ~n2360) | (x6 & ~n2360);
  assign n2363 = n2361 & ~n2362;
  assign n2364 = x1 | n2363;
  assign n2365 = x2 & n1416;
  assign n2366 = x1 & ~n2365;
  assign n2367 = n2364 & ~n2366;
  assign n2388 = n2359 | n2367;
  assign n2389 = ~x3 & n2388;
  assign n2390 = n2387 | n2389;
  assign n2404 = x0 & n2390;
  assign n2391 = (x6 & x8) | (x6 & n265) | (x8 & n265);
  assign n2392 = (x5 & ~x6) | (x5 & n2391) | (~x6 & n2391);
  assign n2393 = (x5 & x8) | (x5 & ~n2391) | (x8 & ~n2391);
  assign n2394 = n2392 & ~n2393;
  assign n2395 = (~x1 & x4) | (~x1 & x5) | (x4 & x5);
  assign n2396 = (~x1 & x5) | (~x1 & x6) | (x5 & x6);
  assign n2397 = n2395 & ~n2396;
  assign n2398 = x3 & n2397;
  assign n2399 = (x0 & x2) | (x0 & n2398) | (x2 & n2398);
  assign n2400 = ~x0 & n2399;
  assign n2401 = (~n36 & n318) | (~n36 & n2400) | (n318 & n2400);
  assign n2402 = n591 & ~n2401;
  assign n2403 = (n591 & n2400) | (n591 & ~n2402) | (n2400 & ~n2402);
  assign n2405 = n2394 | n2403;
  assign n2406 = (n2390 & ~n2404) | (n2390 & n2405) | (~n2404 & n2405);
  assign n2408 = n2345 | n2406;
  assign n2409 = (n2224 & ~n2407) | (n2224 & n2408) | (~n2407 & n2408);
  assign n2410 = (x3 & x4) | (x3 & x5) | (x4 & x5);
  assign n2411 = ~x5 & n2410;
  assign n2412 = (~x4 & n2410) | (~x4 & n2411) | (n2410 & n2411);
  assign n2413 = n43 & n2412;
  assign n2414 = (x1 & x3) | (x1 & ~x5) | (x3 & ~x5);
  assign n2415 = (x0 & ~x1) | (x0 & n2414) | (~x1 & n2414);
  assign n2416 = (x1 & ~x3) | (x1 & n2415) | (~x3 & n2415);
  assign n2417 = ~n2414 & n2416;
  assign n2418 = (~x0 & n2415) | (~x0 & n2417) | (n2415 & n2417);
  assign n2419 = ~x0 & n1073;
  assign n2420 = n79 & n2419;
  assign n2421 = (~n2413 & n2418) | (~n2413 & n2420) | (n2418 & n2420);
  assign n2422 = x2 & ~n2420;
  assign n2423 = (n2413 & n2421) | (n2413 & ~n2422) | (n2421 & ~n2422);
  assign n2576 = n1564 & n2423;
  assign n2427 = ~x7 & n39;
  assign n2428 = (x4 & x6) | (x4 & n2427) | (x6 & n2427);
  assign n2429 = ~x4 & n2428;
  assign n2430 = (~n15 & n552) | (~n15 & n2429) | (n552 & n2429);
  assign n2431 = x4 & ~n2430;
  assign n2432 = (x4 & n2429) | (x4 & ~n2431) | (n2429 & ~n2431);
  assign n2433 = x3 & ~n2432;
  assign n2424 = (x4 & ~x7) | (x4 & n1061) | (~x7 & n1061);
  assign n2425 = (x2 & ~x7) | (x2 & n1061) | (~x7 & n1061);
  assign n2426 = (n519 & n2424) | (n519 & ~n2425) | (n2424 & ~n2425);
  assign n2434 = x6 & n2426;
  assign n2435 = x3 | n2434;
  assign n2436 = ~n2433 & n2435;
  assign n2509 = x8 & n2436;
  assign n2437 = ~n45 & n60;
  assign n2438 = (x1 & ~n378) | (x1 & n2437) | (~n378 & n2437);
  assign n2439 = ~x1 & n2438;
  assign n2474 = (x6 & x7) | (x6 & n53) | (x7 & n53);
  assign n2475 = n1891 & ~n2474;
  assign n2479 = x1 & n2475;
  assign n2476 = (~x5 & x6) | (~x5 & n2131) | (x6 & n2131);
  assign n2477 = (~x5 & x7) | (~x5 & n2131) | (x7 & n2131);
  assign n2478 = (n552 & n2476) | (n552 & ~n2477) | (n2476 & ~n2477);
  assign n2480 = x1 | n2478;
  assign n2481 = (~x1 & n2479) | (~x1 & n2480) | (n2479 & n2480);
  assign n2482 = x8 & ~n2481;
  assign n2471 = (~x3 & n583) | (~x3 & n1918) | (n583 & n1918);
  assign n2472 = (x6 & n1918) | (x6 & ~n2471) | (n1918 & ~n2471);
  assign n2473 = (x3 & n2471) | (x3 & ~n2472) | (n2471 & ~n2472);
  assign n2483 = x5 & n2473;
  assign n2484 = x8 | n2483;
  assign n2485 = ~n2482 & n2484;
  assign n2502 = x2 & n2485;
  assign n2495 = (x3 & n571) | (x3 & n1861) | (n571 & n1861);
  assign n2496 = ~x3 & n2495;
  assign n2491 = (x1 & x7) | (x1 & n890) | (x7 & n890);
  assign n2492 = (x6 & x7) | (x6 & ~n2491) | (x7 & ~n2491);
  assign n2493 = x5 & n2492;
  assign n2494 = (x1 & ~n2491) | (x1 & n2493) | (~n2491 & n2493);
  assign n2497 = (x3 & n2494) | (x3 & n2496) | (n2494 & n2496);
  assign n2498 = x8 & ~n2497;
  assign n2499 = (x8 & n2496) | (x8 & ~n2498) | (n2496 & ~n2498);
  assign n2486 = (x1 & ~x3) | (x1 & x8) | (~x3 & x8);
  assign n2487 = (x1 & ~x7) | (x1 & n2486) | (~x7 & n2486);
  assign n2488 = x1 & ~n2487;
  assign n2489 = n2487 | n2488;
  assign n2490 = (~x1 & n2488) | (~x1 & n2489) | (n2488 & n2489);
  assign n2500 = (x5 & x6) | (x5 & n2490) | (x6 & n2490);
  assign n2501 = (~n591 & n2499) | (~n591 & n2500) | (n2499 & n2500);
  assign n2503 = x2 | n2501;
  assign n2504 = (~x2 & n2502) | (~x2 & n2503) | (n2502 & n2503);
  assign n2505 = x4 & n2504;
  assign n2440 = (x2 & ~x5) | (x2 & n2414) | (~x5 & n2414);
  assign n2441 = x5 & n2440;
  assign n2442 = n2440 & ~n2441;
  assign n2443 = (x5 & ~n2441) | (x5 & n2442) | (~n2441 & n2442);
  assign n2444 = n571 & ~n2443;
  assign n2445 = (n572 & ~n2443) | (n572 & n2444) | (~n2443 & n2444);
  assign n2455 = (x1 & x8) | (x1 & ~n2292) | (x8 & ~n2292);
  assign n2456 = (~x5 & x6) | (~x5 & n2455) | (x6 & n2455);
  assign n2457 = n2292 & n2456;
  assign n2458 = (~n2455 & n2456) | (~n2455 & n2457) | (n2456 & n2457);
  assign n2459 = ~x1 & n571;
  assign n2460 = ~x5 & n2459;
  assign n2461 = x7 & ~n2460;
  assign n2462 = (n2458 & n2460) | (n2458 & ~n2461) | (n2460 & ~n2461);
  assign n2463 = x3 & ~n2462;
  assign n2464 = x1 & n554;
  assign n2465 = x3 | n2464;
  assign n2466 = ~n2463 & n2465;
  assign n2467 = ~x2 & n2466;
  assign n2450 = (x8 & n96) | (x8 & ~n860) | (n96 & ~n860);
  assign n2446 = (~x6 & x7) | (~x6 & n233) | (x7 & n233);
  assign n2447 = (~x3 & x6) | (~x3 & n233) | (x6 & n233);
  assign n2448 = n2446 | n2447;
  assign n2449 = x1 & ~n2448;
  assign n2451 = x8 & n2449;
  assign n2452 = (n860 & n2450) | (n860 & n2451) | (n2450 & n2451);
  assign n2453 = x1 & n571;
  assign n2454 = n53 & n2453;
  assign n2468 = n2452 | n2454;
  assign n2469 = x2 & n2468;
  assign n2470 = n2467 | n2469;
  assign n2506 = n2445 | n2470;
  assign n2507 = ~x4 & n2506;
  assign n2508 = n2505 | n2507;
  assign n2510 = n2439 | n2508;
  assign n2511 = (n2436 & ~n2509) | (n2436 & n2510) | (~n2509 & n2510);
  assign n2538 = x0 & n2511;
  assign n2526 = n1489 & ~n2022;
  assign n2527 = n1104 & n2526;
  assign n2524 = x4 & n45;
  assign n2525 = (n1308 & n1349) | (n1308 & ~n2524) | (n1349 & ~n2524);
  assign n2528 = (~x8 & n2525) | (~x8 & n2527) | (n2525 & n2527);
  assign n2529 = x7 & ~n2528;
  assign n2530 = (x7 & n2527) | (x7 & ~n2529) | (n2527 & ~n2529);
  assign n2531 = x5 & n2530;
  assign n2522 = (x4 & n184) | (x4 & n618) | (n184 & n618);
  assign n2523 = ~x4 & n2522;
  assign n2532 = n2523 | n2531;
  assign n2533 = (~x0 & n2531) | (~x0 & n2532) | (n2531 & n2532);
  assign n2534 = x1 | n2533;
  assign n2512 = (x3 & x4) | (x3 & n299) | (x4 & n299);
  assign n2513 = (~x2 & x4) | (~x2 & n299) | (x4 & n299);
  assign n2514 = (n45 & ~n2512) | (n45 & n2513) | (~n2512 & n2513);
  assign n2515 = ~x8 & n16;
  assign n2516 = n812 & n2515;
  assign n2517 = x5 & ~n2516;
  assign n2518 = (n2514 & ~n2516) | (n2514 & n2517) | (~n2516 & n2517);
  assign n2519 = n21 & n271;
  assign n2520 = x7 | n2519;
  assign n2521 = (~n2518 & n2519) | (~n2518 & n2520) | (n2519 & n2520);
  assign n2535 = ~x0 & n2521;
  assign n2536 = x1 & ~n2535;
  assign n2537 = n2534 & ~n2536;
  assign n2539 = n883 | n2537;
  assign n2540 = (n2511 & ~n2538) | (n2511 & n2539) | (~n2538 & n2539);
  assign n2559 = (x0 & ~x3) | (x0 & n2515) | (~x3 & n2515);
  assign n2555 = (x4 & ~x8) | (x4 & n594) | (~x8 & n594);
  assign n2556 = x4 & ~n2555;
  assign n2557 = n2555 | n2556;
  assign n2558 = (~x4 & n2556) | (~x4 & n2557) | (n2556 & n2557);
  assign n2560 = (x0 & x3) | (x0 & ~n2558) | (x3 & ~n2558);
  assign n2561 = n2559 & ~n2560;
  assign n2562 = x5 & n684;
  assign n2563 = (x0 & n164) | (x0 & n2562) | (n164 & n2562);
  assign n2564 = ~x0 & n2563;
  assign n2565 = ~x5 & n1596;
  assign n2566 = (n1596 & ~n1856) | (n1596 & n2565) | (~n1856 & n2565);
  assign n2567 = (x1 & n1349) | (x1 & n2566) | (n1349 & n2566);
  assign n2568 = ~n2566 & n2567;
  assign n2569 = (~n2561 & n2564) | (~n2561 & n2568) | (n2564 & n2568);
  assign n2570 = x1 & ~n2568;
  assign n2571 = (n2561 & n2569) | (n2561 & ~n2570) | (n2569 & ~n2570);
  assign n2572 = x2 | n2571;
  assign n2541 = (x3 & x5) | (x3 & ~x8) | (x5 & ~x8);
  assign n2542 = (~x3 & x6) | (~x3 & n2541) | (x6 & n2541);
  assign n2543 = (x5 & x6) | (x5 & ~n2541) | (x6 & ~n2541);
  assign n2544 = n2542 & ~n2543;
  assign n2549 = (x1 & ~x4) | (x1 & n2544) | (~x4 & n2544);
  assign n2545 = (x3 & x5) | (x3 & x8) | (x5 & x8);
  assign n2546 = (x3 & x6) | (x3 & ~n2545) | (x6 & ~n2545);
  assign n2547 = (~x5 & x6) | (~x5 & n2545) | (x6 & n2545);
  assign n2548 = ~n2546 & n2547;
  assign n2550 = (x1 & x4) | (x1 & ~n2548) | (x4 & ~n2548);
  assign n2551 = n2549 & ~n2550;
  assign n2552 = (~x1 & n20) | (~x1 & n2551) | (n20 & n2551);
  assign n2553 = n1021 | n2552;
  assign n2554 = (~n1021 & n2551) | (~n1021 & n2553) | (n2551 & n2553);
  assign n2573 = ~x0 & n2554;
  assign n2574 = x2 & ~n2573;
  assign n2575 = n2572 & ~n2574;
  assign n2577 = n2540 | n2575;
  assign n2578 = (n2423 & ~n2576) | (n2423 & n2577) | (~n2576 & n2577);
  assign n2579 = (x5 & ~x8) | (x5 & n1623) | (~x8 & n1623);
  assign n2580 = (x1 & x4) | (x1 & n2579) | (x4 & n2579);
  assign n2581 = ~n1623 & n2580;
  assign n2582 = (~n2579 & n2580) | (~n2579 & n2581) | (n2580 & n2581);
  assign n2583 = x3 & ~n2582;
  assign n2584 = ~x1 & n1595;
  assign n2585 = x3 | n2584;
  assign n2586 = ~n2583 & n2585;
  assign n2596 = (~x0 & x2) | (~x0 & n2586) | (x2 & n2586);
  assign n2588 = x3 & ~n1483;
  assign n2589 = ~x5 & n2588;
  assign n2590 = (x8 & ~n1483) | (x8 & n2588) | (~n1483 & n2588);
  assign n2591 = (x1 & n2589) | (x1 & n2590) | (n2589 & n2590);
  assign n2592 = x4 | n2591;
  assign n2587 = x8 | n1415;
  assign n2593 = x1 & ~n2587;
  assign n2594 = x4 & ~n2593;
  assign n2595 = n2592 & ~n2594;
  assign n2597 = (x0 & x2) | (x0 & ~n2595) | (x2 & ~n2595);
  assign n2598 = n2596 & ~n2597;
  assign n2599 = (x5 & ~n318) | (x5 & n387) | (~n318 & n387);
  assign n2600 = n318 & n2599;
  assign n2601 = n2598 | n2600;
  assign n2602 = (~x6 & x7) | (~x6 & n2601) | (x7 & n2601);
  assign n2603 = (n552 & n2601) | (n552 & ~n2602) | (n2601 & ~n2602);
  assign n2638 = (~x6 & x8) | (~x6 & n237) | (x8 & n237);
  assign n2639 = x8 & ~n2638;
  assign n2640 = n2638 | n2639;
  assign n2641 = (~x8 & n2639) | (~x8 & n2640) | (n2639 & n2640);
  assign n2642 = x4 & n2641;
  assign n2643 = x1 & ~n2642;
  assign n2644 = ~n77 & n80;
  assign n2645 = x1 | n2644;
  assign n2646 = ~n2643 & n2645;
  assign n2661 = (~x0 & x2) | (~x0 & n2646) | (x2 & n2646);
  assign n2650 = (x6 & ~x7) | (x6 & n1000) | (~x7 & n1000);
  assign n2651 = x6 & ~n2650;
  assign n2652 = n2650 | n2651;
  assign n2653 = (~x6 & n2651) | (~x6 & n2652) | (n2651 & n2652);
  assign n2654 = x1 | n2653;
  assign n2655 = x1 & ~n1254;
  assign n2656 = n2654 & ~n2655;
  assign n2657 = x3 | n2656;
  assign n2647 = (~x4 & x7) | (~x4 & n1515) | (x7 & n1515);
  assign n2648 = (~x7 & x8) | (~x7 & n1515) | (x8 & n1515);
  assign n2649 = n2647 & n2648;
  assign n2658 = x1 & n2649;
  assign n2659 = x3 & ~n2658;
  assign n2660 = n2657 & ~n2659;
  assign n2662 = (x0 & x2) | (x0 & ~n2660) | (x2 & ~n2660);
  assign n2663 = n2661 & ~n2662;
  assign n2664 = (n10 & n46) | (n10 & n2663) | (n46 & n2663);
  assign n2665 = n378 | n2664;
  assign n2666 = (~n378 & n2663) | (~n378 & n2665) | (n2663 & n2665);
  assign n2614 = (x0 & x3) | (x0 & ~x4) | (x3 & ~x4);
  assign n2615 = (x0 & x3) | (x0 & ~x5) | (x3 & ~x5);
  assign n2616 = n2614 & n2615;
  assign n2617 = x5 | n2616;
  assign n2618 = (~n2614 & n2616) | (~n2614 & n2617) | (n2616 & n2617);
  assign n2621 = (~x2 & x6) | (~x2 & n2618) | (x6 & n2618);
  assign n2619 = (x2 & n1105) | (x2 & n1415) | (n1105 & n1415);
  assign n2620 = ~n1415 & n2619;
  assign n2622 = x6 & n2620;
  assign n2623 = (~n2618 & n2621) | (~n2618 & n2622) | (n2621 & n2622);
  assign n2611 = ~x3 & n2137;
  assign n2612 = (x2 & x5) | (x2 & ~n2611) | (x5 & ~n2611);
  assign n2613 = (n2137 & n2611) | (n2137 & ~n2612) | (n2611 & ~n2612);
  assign n2624 = (~x0 & n2613) | (~x0 & n2623) | (n2613 & n2623);
  assign n2625 = x4 & ~n2624;
  assign n2626 = (x4 & n2623) | (x4 & ~n2625) | (n2623 & ~n2625);
  assign n2627 = (x2 & x5) | (x2 & ~x7) | (x5 & ~x7);
  assign n2628 = ~n225 & n2627;
  assign n2629 = ~x4 & n2628;
  assign n2630 = (x0 & ~x6) | (x0 & n2629) | (~x6 & n2629);
  assign n2631 = ~x0 & n2630;
  assign n2632 = x7 | n2631;
  assign n2633 = (n2626 & n2631) | (n2626 & n2632) | (n2631 & n2632);
  assign n2634 = x1 | n2633;
  assign n2604 = (x4 & x5) | (x4 & x7) | (x5 & x7);
  assign n2605 = n2022 & ~n2604;
  assign n2608 = (x2 & ~x6) | (x2 & n2605) | (~x6 & n2605);
  assign n2606 = x4 & n42;
  assign n2607 = n187 & n2606;
  assign n2609 = ~x6 & n2607;
  assign n2610 = (~x2 & n2608) | (~x2 & n2609) | (n2608 & n2609);
  assign n2635 = ~x0 & n2610;
  assign n2636 = x1 & ~n2635;
  assign n2637 = n2634 & ~n2636;
  assign n2707 = (~x3 & x5) | (~x3 & n1480) | (x5 & n1480);
  assign n2708 = (x1 & x7) | (x1 & n2707) | (x7 & n2707);
  assign n2709 = ~n1480 & n2708;
  assign n2710 = (~n2707 & n2708) | (~n2707 & n2709) | (n2708 & n2709);
  assign n2711 = x4 & n2710;
  assign n2712 = ~x0 & n2711;
  assign n2713 = (~x4 & n187) | (~x4 & n2712) | (n187 & n2712);
  assign n2714 = n1355 & ~n2713;
  assign n2715 = (n1355 & n2712) | (n1355 & ~n2714) | (n2712 & ~n2714);
  assign n2743 = ~n337 & n787;
  assign n2741 = (x5 & ~n43) | (x5 & n1803) | (~n43 & n1803);
  assign n2742 = n43 & n2741;
  assign n2744 = (x3 & ~x5) | (x3 & x7) | (~x5 & x7);
  assign n2745 = (x1 & x5) | (x1 & n2744) | (x5 & n2744);
  assign n2746 = (x5 & x7) | (x5 & ~n2745) | (x7 & ~n2745);
  assign n2747 = n2744 | n2746;
  assign n2748 = (x1 & ~n2745) | (x1 & n2747) | (~n2745 & n2747);
  assign n2753 = (x0 & ~x4) | (x0 & n2748) | (~x4 & n2748);
  assign n2749 = (x3 & ~x5) | (x3 & n1480) | (~x5 & n1480);
  assign n2750 = x3 & ~n2749;
  assign n2751 = n2749 | n2750;
  assign n2752 = (~x3 & n2750) | (~x3 & n2751) | (n2750 & n2751);
  assign n2754 = (x0 & x4) | (x0 & ~n2752) | (x4 & ~n2752);
  assign n2755 = n2753 | n2754;
  assign n2756 = ~n2742 & n2755;
  assign n2757 = ~n2743 & n2756;
  assign n2758 = ~x6 & n2757;
  assign n2733 = (x1 & x5) | (x1 & ~x7) | (x5 & ~x7);
  assign n2734 = (~x1 & x7) | (~x1 & n2733) | (x7 & n2733);
  assign n2735 = (~x3 & x7) | (~x3 & n2734) | (x7 & n2734);
  assign n2736 = (~n53 & n2733) | (~n53 & n2735) | (n2733 & n2735);
  assign n2737 = ~x4 & n2736;
  assign n2738 = n96 & n187;
  assign n2739 = x4 & ~n2738;
  assign n2740 = n2737 | n2739;
  assign n2759 = x0 | n2740;
  assign n2760 = x6 & n2759;
  assign n2761 = n2758 | n2760;
  assign n2762 = x8 & n2761;
  assign n2722 = (~x3 & x5) | (~x3 & n437) | (x5 & n437);
  assign n2723 = (x4 & x5) | (x4 & ~n437) | (x5 & ~n437);
  assign n2724 = (~x3 & x7) | (~x3 & n2723) | (x7 & n2723);
  assign n2725 = ~n2722 & n2724;
  assign n2726 = x1 & n2725;
  assign n2718 = (x3 & x5) | (x3 & ~n1571) | (x5 & ~n1571);
  assign n2719 = (x4 & ~x7) | (x4 & n2718) | (~x7 & n2718);
  assign n2720 = n1571 & n2719;
  assign n2721 = (~n2718 & n2719) | (~n2718 & n2720) | (n2719 & n2720);
  assign n2727 = x1 | n2721;
  assign n2728 = (~x1 & n2726) | (~x1 & n2727) | (n2726 & n2727);
  assign n2729 = x6 & ~n2728;
  assign n2716 = x7 & ~n20;
  assign n2717 = (~n755 & n765) | (~n755 & n2716) | (n765 & n2716);
  assign n2730 = x1 & ~n2717;
  assign n2731 = x6 | n2730;
  assign n2732 = ~n2729 & n2731;
  assign n2763 = ~x0 & n2732;
  assign n2764 = x8 | n2763;
  assign n2765 = ~n2762 & n2764;
  assign n2766 = n738 & ~n2765;
  assign n2767 = (n2715 & n2765) | (n2715 & ~n2766) | (n2765 & ~n2766);
  assign n2768 = x2 | n2767;
  assign n2694 = n60 | n78;
  assign n2695 = (n37 & n78) | (n37 & n2694) | (n78 & n2694);
  assign n2696 = x1 & ~n2695;
  assign n2697 = x5 & n572;
  assign n2698 = x1 | n2697;
  assign n2699 = ~n2696 & n2698;
  assign n2689 = (x3 & ~x6) | (x3 & x8) | (~x6 & x8);
  assign n2690 = (~x3 & x6) | (~x3 & n2689) | (x6 & n2689);
  assign n2691 = ~x1 & n2689;
  assign n2692 = (~x8 & n2689) | (~x8 & n2691) | (n2689 & n2691);
  assign n2693 = n2690 | n2692;
  assign n2700 = (x5 & ~n2693) | (x5 & n2699) | (~n2693 & n2699);
  assign n2701 = x7 & ~n2700;
  assign n2702 = (x7 & n2699) | (x7 & ~n2701) | (n2699 & ~n2701);
  assign n2703 = ~x4 & n2702;
  assign n2667 = (x1 & x5) | (x1 & ~n60) | (x5 & ~n60);
  assign n2668 = (~x1 & x7) | (~x1 & n2667) | (x7 & n2667);
  assign n2669 = (~x5 & x8) | (~x5 & n2668) | (x8 & n2668);
  assign n2670 = n2667 & n2669;
  assign n2675 = (~x3 & x6) | (~x3 & n2670) | (x6 & n2670);
  assign n2671 = (x1 & x7) | (x1 & n656) | (x7 & n656);
  assign n2672 = (x3 & ~x7) | (x3 & n2671) | (~x7 & n2671);
  assign n2673 = (x1 & x3) | (x1 & ~n2671) | (x3 & ~n2671);
  assign n2674 = n2672 & ~n2673;
  assign n2676 = ~x6 & n2674;
  assign n2677 = (n2670 & ~n2675) | (n2670 & n2676) | (~n2675 & n2676);
  assign n2678 = (x1 & x7) | (x1 & x8) | (x7 & x8);
  assign n2679 = (~x3 & x8) | (~x3 & n2678) | (x8 & n2678);
  assign n2680 = x8 & ~n2679;
  assign n2681 = n2679 | n2680;
  assign n2682 = (~x8 & n2680) | (~x8 & n2681) | (n2680 & n2681);
  assign n2686 = (x5 & x6) | (x5 & ~n2682) | (x6 & ~n2682);
  assign n2683 = (x1 & x7) | (x1 & ~n1593) | (x7 & ~n1593);
  assign n2684 = x1 & ~n2683;
  assign n2685 = (x7 & ~n2683) | (x7 & n2684) | (~n2683 & n2684);
  assign n2687 = x6 & n2685;
  assign n2688 = (n2682 & n2686) | (n2682 & n2687) | (n2686 & n2687);
  assign n2704 = n2677 | n2688;
  assign n2705 = x4 & n2704;
  assign n2706 = n2703 | n2705;
  assign n2769 = ~x0 & n2706;
  assign n2770 = x2 & ~n2769;
  assign n2771 = n2768 & ~n2770;
  assign n2772 = n2637 | n2771;
  assign n2773 = (~n2603 & n2666) | (~n2603 & n2772) | (n2666 & n2772);
  assign n2774 = n2603 | n2773;
  assign n2786 = ~x3 & n380;
  assign n2800 = n44 & ~n2786;
  assign n2787 = x2 & n43;
  assign n2788 = (x3 & x8) | (x3 & n2787) | (x8 & n2787);
  assign n2789 = ~x8 & n2788;
  assign n2794 = (x2 & x8) | (x2 & ~n1522) | (x8 & ~n1522);
  assign n2795 = (x2 & x5) | (x2 & ~n1522) | (x5 & ~n1522);
  assign n2796 = (n655 & n2794) | (n655 & ~n2795) | (n2794 & ~n2795);
  assign n2797 = (~x0 & x3) | (~x0 & n2796) | (x3 & n2796);
  assign n2790 = (x1 & ~x5) | (x1 & x8) | (~x5 & x8);
  assign n2791 = ~x1 & n2790;
  assign n2792 = (x2 & x8) | (x2 & ~n2791) | (x8 & ~n2791);
  assign n2793 = (n2790 & n2791) | (n2790 & ~n2792) | (n2791 & ~n2792);
  assign n2798 = (x0 & x3) | (x0 & ~n2793) | (x3 & ~n2793);
  assign n2799 = n2797 & ~n2798;
  assign n2801 = n2789 | n2799;
  assign n2802 = (n44 & ~n2800) | (n44 & n2801) | (~n2800 & n2801);
  assign n2803 = x4 & n2802;
  assign n2775 = (x0 & x5) | (x0 & x8) | (x5 & x8);
  assign n2776 = (~x0 & x3) | (~x0 & n2775) | (x3 & n2775);
  assign n2777 = (x5 & x8) | (x5 & n2776) | (x8 & n2776);
  assign n2778 = n2775 & ~n2777;
  assign n2779 = (n2776 & ~n2777) | (n2776 & n2778) | (~n2777 & n2778);
  assign n2781 = (x1 & x2) | (x1 & n2779) | (x2 & n2779);
  assign n2780 = n43 & ~n2587;
  assign n2782 = ~x2 & n2780;
  assign n2783 = (n2779 & ~n2781) | (n2779 & n2782) | (~n2781 & n2782);
  assign n2784 = (x5 & ~n40) | (x5 & n1598) | (~n40 & n1598);
  assign n2785 = n40 & n2784;
  assign n2804 = n2783 | n2785;
  assign n2805 = ~x4 & n2804;
  assign n2806 = n2803 | n2805;
  assign n2807 = (x6 & x7) | (x6 & ~n2806) | (x7 & ~n2806);
  assign n2808 = x6 & ~n2807;
  assign n2809 = (x7 & ~n2807) | (x7 & n2808) | (~n2807 & n2808);
  assign n2907 = x0 & ~x7;
  assign n2908 = x4 & ~n2907;
  assign n2909 = (n60 & n712) | (n60 & ~n2908) | (n712 & ~n2908);
  assign n2910 = x6 & ~n2909;
  assign n2911 = x0 | n811;
  assign n2912 = ~x6 & n2911;
  assign n2913 = n2910 | n2912;
  assign n2914 = ~x3 & n2913;
  assign n2903 = ~x8 & n214;
  assign n2904 = (x6 & x8) | (x6 & ~n214) | (x8 & ~n214);
  assign n2905 = n2903 | n2904;
  assign n2906 = (x8 & n2903) | (x8 & n2905) | (n2903 & n2905);
  assign n2915 = x0 | n2906;
  assign n2916 = x3 & n2915;
  assign n2917 = n2914 | n2916;
  assign n2918 = ~x2 & n2917;
  assign n2896 = (~x7 & x8) | (~x7 & n1561) | (x8 & n1561);
  assign n2897 = (~x4 & x8) | (~x4 & n1561) | (x8 & n1561);
  assign n2898 = (n86 & ~n2896) | (n86 & n2897) | (~n2896 & n2897);
  assign n2899 = x6 | n2898;
  assign n2900 = ~x4 & n29;
  assign n2901 = x6 & ~n2900;
  assign n2902 = n2899 & ~n2901;
  assign n2919 = ~x0 & n2902;
  assign n2920 = x2 & ~n2919;
  assign n2921 = n2918 | n2920;
  assign n2922 = ~x1 & n2921;
  assign n2875 = (x3 & x6) | (x3 & x7) | (x6 & x7);
  assign n2876 = (x3 & x8) | (x3 & ~n2875) | (x8 & ~n2875);
  assign n2877 = (~x3 & x6) | (~x3 & n2876) | (x6 & n2876);
  assign n2878 = n2875 | n2877;
  assign n2879 = (~x8 & n2876) | (~x8 & n2878) | (n2876 & n2878);
  assign n2880 = x4 & ~n2879;
  assign n2874 = (x3 & ~n375) | (x3 & n1506) | (~n375 & n1506);
  assign n2881 = x4 | n2874;
  assign n2882 = (~x4 & n2880) | (~x4 & n2881) | (n2880 & n2881);
  assign n2893 = x2 & n2882;
  assign n2883 = x8 & ~n184;
  assign n2884 = ~x6 & n2883;
  assign n2885 = (x3 & ~n184) | (x3 & n2883) | (~n184 & n2883);
  assign n2886 = (~x7 & n2884) | (~x7 & n2885) | (n2884 & n2885);
  assign n2890 = x4 & ~n2886;
  assign n2887 = (x3 & x7) | (x3 & n738) | (x7 & n738);
  assign n2888 = x3 & ~n2887;
  assign n2889 = (x7 & ~n2887) | (x7 & n2888) | (~n2887 & n2888);
  assign n2891 = ~x4 & n2889;
  assign n2892 = (x4 & ~n2890) | (x4 & n2891) | (~n2890 & n2891);
  assign n2894 = x2 | n2892;
  assign n2895 = (~x2 & n2893) | (~x2 & n2894) | (n2893 & n2894);
  assign n2923 = ~x0 & n2895;
  assign n2924 = x1 & ~n2923;
  assign n2925 = n2922 | n2924;
  assign n2926 = x5 & n2925;
  assign n2851 = (~x1 & x3) | (~x1 & x6) | (x3 & x6);
  assign n2852 = x1 & n2851;
  assign n2853 = (~n1437 & n2851) | (~n1437 & n2852) | (n2851 & n2852);
  assign n2854 = x3 | x6;
  assign n2857 = (~x3 & x7) | (~x3 & n2854) | (x7 & n2854);
  assign n2858 = (x7 & x8) | (x7 & n2854) | (x8 & n2854);
  assign n2859 = (n2242 & n2857) | (n2242 & ~n2858) | (n2857 & ~n2858);
  assign n2860 = x2 & n2859;
  assign n2861 = x3 & n257;
  assign n2862 = x2 | n2861;
  assign n2863 = ~n2860 & n2862;
  assign n2864 = x1 & ~n2863;
  assign n2855 = x7 & ~n812;
  assign n2856 = (~n583 & n2854) | (~n583 & n2855) | (n2854 & n2855);
  assign n2865 = x8 | n2856;
  assign n2866 = ~x1 & n2865;
  assign n2867 = n2864 | n2866;
  assign n2850 = (n10 & n380) | (n10 & ~n1712) | (n380 & ~n1712);
  assign n2868 = ~n2850 & n2867;
  assign n2869 = (~n2853 & n2867) | (~n2853 & n2868) | (n2867 & n2868);
  assign n2870 = x4 & ~n2869;
  assign n2840 = (~x6 & x8) | (~x6 & n1696) | (x8 & n1696);
  assign n2841 = x8 & ~n2840;
  assign n2842 = n2840 | n2841;
  assign n2843 = (~x8 & n2841) | (~x8 & n2842) | (n2841 & n2842);
  assign n2844 = (~x1 & x3) | (~x1 & n2843) | (x3 & n2843);
  assign n2838 = (n184 & n685) | (n184 & ~n2374) | (n685 & ~n2374);
  assign n2839 = (x7 & n184) | (x7 & n2838) | (n184 & n2838);
  assign n2845 = (x1 & x3) | (x1 & n2839) | (x3 & n2839);
  assign n2846 = n2844 & n2845;
  assign n2847 = x3 | n375;
  assign n2848 = (x1 & x2) | (x1 & ~n2847) | (x2 & ~n2847);
  assign n2849 = ~x1 & n2848;
  assign n2871 = n2846 | n2849;
  assign n2872 = ~x4 & n2871;
  assign n2873 = n2870 | n2872;
  assign n2927 = ~x0 & n2873;
  assign n2928 = x5 | n2927;
  assign n2929 = ~n2926 & n2928;
  assign n2819 = (x0 & x4) | (x0 & n129) | (x4 & n129);
  assign n2820 = (x4 & x7) | (x4 & ~n2819) | (x7 & ~n2819);
  assign n2821 = (x0 & ~x5) | (x0 & n2820) | (~x5 & n2820);
  assign n2822 = ~n2819 & n2821;
  assign n2823 = x1 | n2822;
  assign n2824 = ~x0 & n445;
  assign n2825 = x1 & ~n2824;
  assign n2826 = n2823 & ~n2825;
  assign n2827 = x2 | n2826;
  assign n2816 = (~x1 & x4) | (~x1 & n969) | (x4 & n969);
  assign n2817 = (~x4 & x5) | (~x4 & n969) | (x5 & n969);
  assign n2818 = n2816 & n2817;
  assign n2828 = ~x0 & n2818;
  assign n2829 = x2 & ~n2828;
  assign n2830 = n2827 & ~n2829;
  assign n2831 = x3 | n2830;
  assign n2810 = (x1 & ~x2) | (x1 & n750) | (~x2 & n750);
  assign n2811 = (x1 & x2) | (x1 & n1839) | (x2 & n1839);
  assign n2812 = ~n2810 & n2811;
  assign n2813 = (~x4 & n129) | (~x4 & n2812) | (n129 & n2812);
  assign n2814 = n487 & ~n2813;
  assign n2815 = (n487 & n2812) | (n487 & ~n2814) | (n2812 & ~n2814);
  assign n2832 = ~x0 & n2815;
  assign n2833 = x3 & ~n2832;
  assign n2834 = n2831 & ~n2833;
  assign n2835 = (x6 & x8) | (x6 & ~n2834) | (x8 & ~n2834);
  assign n2836 = x6 & ~n2835;
  assign n2837 = (x8 & ~n2835) | (x8 & n2836) | (~n2835 & n2836);
  assign n2946 = (x0 & ~x1) | (x0 & x2) | (~x1 & x2);
  assign n2947 = (x1 & ~x5) | (x1 & n2946) | (~x5 & n2946);
  assign n2948 = (x0 & x2) | (x0 & n2947) | (x2 & n2947);
  assign n2949 = n2946 & ~n2948;
  assign n2950 = (n2947 & ~n2948) | (n2947 & n2949) | (~n2948 & n2949);
  assign n2951 = (~x4 & x7) | (~x4 & n2950) | (x7 & n2950);
  assign n2952 = (x6 & ~x7) | (x6 & n2951) | (~x7 & n2951);
  assign n2953 = (x4 & ~x6) | (x4 & n2951) | (~x6 & n2951);
  assign n2954 = n2952 & n2953;
  assign n2955 = (x2 & x6) | (x2 & ~n755) | (x6 & ~n755);
  assign n2956 = (~x2 & x5) | (~x2 & n2955) | (x5 & n2955);
  assign n2957 = (~x6 & x7) | (~x6 & n2956) | (x7 & n2956);
  assign n2958 = n2955 & n2957;
  assign n2959 = (x4 & ~n43) | (x4 & n2958) | (~n43 & n2958);
  assign n2960 = n2958 & ~n2959;
  assign n2961 = n2954 | n2960;
  assign n2962 = x3 | n2961;
  assign n2937 = x7 & ~n519;
  assign n2938 = (~n583 & n1287) | (~n583 & n2937) | (n1287 & n2937);
  assign n2939 = x1 & ~n2938;
  assign n2933 = (x2 & ~x4) | (x2 & n552) | (~x4 & n552);
  assign n2934 = (x4 & x6) | (x4 & n552) | (x6 & n552);
  assign n2935 = (x2 & x7) | (x2 & ~n2934) | (x7 & ~n2934);
  assign n2936 = ~n2933 & n2935;
  assign n2940 = x1 | n2936;
  assign n2941 = (~x1 & n2939) | (~x1 & n2940) | (n2939 & n2940);
  assign n2942 = x5 | n2941;
  assign n2930 = x1 & x6;
  assign n2931 = x7 | n79;
  assign n2932 = (~n564 & n2930) | (~n564 & n2931) | (n2930 & n2931);
  assign n2943 = ~x4 & n2932;
  assign n2944 = x5 & ~n2943;
  assign n2945 = n2942 & ~n2944;
  assign n2963 = ~x0 & n2945;
  assign n2964 = x3 & ~n2963;
  assign n2965 = n2962 & ~n2964;
  assign n2966 = n2837 | n2965;
  assign n2967 = (~n2809 & n2929) | (~n2809 & n2966) | (n2929 & n2966);
  assign n2968 = n2809 | n2967;
  assign n2972 = (n40 & n1643) | (n40 & ~n1790) | (n1643 & ~n1790);
  assign n2969 = (x1 & ~x3) | (x1 & n1712) | (~x3 & n1712);
  assign n2970 = ~x1 & n2969;
  assign n2971 = x0 & n2970;
  assign n2973 = n1643 & n2971;
  assign n2974 = (n1790 & n2972) | (n1790 & n2973) | (n2972 & n2973);
  assign n3032 = ~x8 & n80;
  assign n3033 = x5 & n3032;
  assign n3034 = (~x1 & x3) | (~x1 & x5) | (x3 & x5);
  assign n3035 = (x5 & x8) | (x5 & ~n3034) | (x8 & ~n3034);
  assign n3036 = (x1 & ~x3) | (x1 & n3035) | (~x3 & n3035);
  assign n3037 = n3034 & n3036;
  assign n3038 = (~n3035 & n3036) | (~n3035 & n3037) | (n3036 & n3037);
  assign n3039 = ~x4 & n3038;
  assign n3040 = ~x0 & n3039;
  assign n3041 = n1595 | n3040;
  assign n3042 = (n1355 & n3040) | (n1355 & n3041) | (n3040 & n3041);
  assign n3043 = ~x2 & n3042;
  assign n3044 = n40 | n3043;
  assign n3045 = (n3033 & n3043) | (n3033 & n3044) | (n3043 & n3044);
  assign n3011 = (x0 & x6) | (x0 & ~x8) | (x6 & ~x8);
  assign n3012 = (x4 & ~x6) | (x4 & n3011) | (~x6 & n3011);
  assign n3013 = (x0 & ~x8) | (x0 & n3012) | (~x8 & n3012);
  assign n3014 = ~n3011 & n3013;
  assign n3015 = (~n3012 & n3013) | (~n3012 & n3014) | (n3013 & n3014);
  assign n3016 = x2 | n3015;
  assign n3010 = x4 & n994;
  assign n3017 = ~x0 & n3010;
  assign n3018 = x2 & ~n3017;
  assign n3019 = n3016 & ~n3018;
  assign n3020 = x1 | n3019;
  assign n3005 = x2 & x8;
  assign n3006 = (x4 & x6) | (x4 & n3005) | (x6 & n3005);
  assign n3007 = (x6 & x8) | (x6 & ~n3006) | (x8 & ~n3006);
  assign n3008 = (x2 & x4) | (x2 & n3007) | (x4 & n3007);
  assign n3009 = ~n3006 & n3008;
  assign n3021 = ~x0 & n3009;
  assign n3022 = x1 & ~n3021;
  assign n3023 = n3020 & ~n3022;
  assign n3024 = x5 | n3023;
  assign n2998 = (x2 & x4) | (x2 & x6) | (x4 & x6);
  assign n2999 = (x4 & x6) | (x4 & ~n2998) | (x6 & ~n2998);
  assign n3000 = (x1 & x4) | (x1 & n2999) | (x4 & n2999);
  assign n3001 = (n487 & n2998) | (n487 & ~n3000) | (n2998 & ~n3000);
  assign n3002 = n39 & n376;
  assign n3003 = x8 | n3002;
  assign n3004 = (n3001 & n3002) | (n3001 & n3003) | (n3002 & n3003);
  assign n3025 = ~x0 & n3004;
  assign n3026 = x5 & ~n3025;
  assign n3027 = n3024 & ~n3026;
  assign n3028 = x3 | n3027;
  assign n2975 = (x6 & ~x8) | (x6 & n634) | (~x8 & n634);
  assign n2976 = (x1 & x6) | (x1 & n634) | (x6 & n634);
  assign n2977 = (n1387 & n2975) | (n1387 & ~n2976) | (n2975 & ~n2976);
  assign n2983 = x4 & n2977;
  assign n2978 = (x1 & ~x6) | (x1 & x8) | (~x6 & x8);
  assign n2979 = (~x5 & x8) | (~x5 & n2978) | (x8 & n2978);
  assign n2980 = x8 & ~n2979;
  assign n2981 = n2979 | n2980;
  assign n2982 = (~x8 & n2980) | (~x8 & n2981) | (n2980 & n2981);
  assign n2984 = x4 | n2982;
  assign n2985 = (~x4 & n2983) | (~x4 & n2984) | (n2983 & n2984);
  assign n2995 = x2 & n2985;
  assign n2987 = (x1 & x6) | (x1 & ~n2790) | (x6 & ~n2790);
  assign n2988 = (x5 & ~x8) | (x5 & n2987) | (~x8 & n2987);
  assign n2989 = n2790 & n2988;
  assign n2990 = (~n2987 & n2988) | (~n2987 & n2989) | (n2988 & n2989);
  assign n2991 = x4 & ~n2990;
  assign n2986 = n1223 | n1541;
  assign n2992 = ~x1 & n2986;
  assign n2993 = x4 | n2992;
  assign n2994 = ~n2991 & n2993;
  assign n2996 = x2 | n2994;
  assign n2997 = (~x2 & n2995) | (~x2 & n2996) | (n2995 & n2996);
  assign n3029 = ~x0 & n2997;
  assign n3030 = x3 & ~n3029;
  assign n3031 = n3028 & ~n3030;
  assign n3054 = n318 & n684;
  assign n3055 = n53 & n3054;
  assign n3046 = (~x1 & x6) | (~x1 & n634) | (x6 & n634);
  assign n3047 = (x6 & x8) | (x6 & ~n634) | (x8 & ~n634);
  assign n3048 = (~x1 & x5) | (~x1 & n3047) | (x5 & n3047);
  assign n3049 = ~n3046 & n3048;
  assign n3050 = x3 | n3049;
  assign n3051 = x1 | n1021;
  assign n3052 = x3 & n3051;
  assign n3053 = n3050 & ~n3052;
  assign n3056 = (~x0 & n3053) | (~x0 & n3055) | (n3053 & n3055);
  assign n3057 = x2 & ~n3056;
  assign n3058 = (x2 & n3055) | (x2 & ~n3057) | (n3055 & ~n3057);
  assign n3158 = n215 & n3058;
  assign n3079 = n1582 & ~n2689;
  assign n3080 = x6 & n118;
  assign n3081 = (x6 & n851) | (x6 & ~n3080) | (n851 & ~n3080);
  assign n3082 = (x3 & ~x8) | (x3 & n3081) | (~x8 & n3081);
  assign n3083 = (~x7 & x8) | (~x7 & n3082) | (x8 & n3082);
  assign n3084 = (~x3 & x7) | (~x3 & n3082) | (x7 & n3082);
  assign n3085 = n3083 | n3084;
  assign n3086 = (x4 & x5) | (x4 & n3085) | (x5 & n3085);
  assign n3087 = n3079 & n3086;
  assign n3088 = (~n3079 & n3085) | (~n3079 & n3087) | (n3085 & n3087);
  assign n3089 = x2 & ~n3088;
  assign n3059 = (x5 & x6) | (x5 & ~x7) | (x6 & ~x7);
  assign n3060 = x8 | n3059;
  assign n3061 = ~n658 & n3060;
  assign n3066 = (x3 & ~x4) | (x3 & n3061) | (~x4 & n3061);
  assign n3062 = (x5 & n70) | (x5 & n184) | (n70 & n184);
  assign n3063 = (~x5 & x7) | (~x5 & n3062) | (x7 & n3062);
  assign n3064 = (~x8 & n70) | (~x8 & n3063) | (n70 & n3063);
  assign n3065 = (~n70 & n3062) | (~n70 & n3064) | (n3062 & n3064);
  assign n3067 = (x3 & x4) | (x3 & ~n3065) | (x4 & ~n3065);
  assign n3068 = n3066 & ~n3067;
  assign n3069 = (x6 & x8) | (x6 & n337) | (x8 & n337);
  assign n3070 = (x5 & x6) | (x5 & ~n3069) | (x6 & ~n3069);
  assign n3071 = (x7 & x8) | (x7 & n3070) | (x8 & n3070);
  assign n3072 = n3069 & ~n3071;
  assign n3076 = (~x3 & x4) | (~x3 & n3072) | (x4 & n3072);
  assign n3073 = (x7 & x8) | (x7 & n640) | (x8 & n640);
  assign n3074 = (x5 & x8) | (x5 & n640) | (x8 & n640);
  assign n3075 = (n187 & n3073) | (n187 & ~n3074) | (n3073 & ~n3074);
  assign n3077 = (x3 & x4) | (x3 & n3075) | (x4 & n3075);
  assign n3078 = n3076 & n3077;
  assign n3090 = n3068 | n3078;
  assign n3091 = ~x2 & n3090;
  assign n3092 = n3089 | n3091;
  assign n3129 = (~x0 & x1) | (~x0 & n3092) | (x1 & n3092);
  assign n3116 = n20 & n571;
  assign n3113 = x6 | n1494;
  assign n3114 = (x6 & ~x8) | (x6 & n1494) | (~x8 & n1494);
  assign n3115 = (x8 & ~n3113) | (x8 & n3114) | (~n3113 & n3114);
  assign n3117 = n3115 | n3116;
  assign n3118 = (~x7 & n3116) | (~x7 & n3117) | (n3116 & n3117);
  assign n3119 = x2 | n3118;
  assign n3110 = ~x8 & n237;
  assign n3111 = (x3 & x4) | (x3 & ~n3110) | (x4 & ~n3110);
  assign n3112 = (n237 & n3110) | (n237 & ~n3111) | (n3110 & ~n3111);
  assign n3120 = x6 & n3112;
  assign n3121 = x2 & ~n3120;
  assign n3122 = n3119 & ~n3121;
  assign n3106 = (x4 & ~x6) | (x4 & n1494) | (~x6 & n1494);
  assign n3107 = x4 & ~n3106;
  assign n3108 = n3106 | n3107;
  assign n3109 = (~x4 & n3107) | (~x4 & n3108) | (n3107 & n3108);
  assign n3123 = (~x2 & x7) | (~x2 & n3109) | (x7 & n3109);
  assign n3124 = (~n1712 & n3122) | (~n1712 & n3123) | (n3122 & n3123);
  assign n3125 = ~x5 & n3124;
  assign n3095 = (x3 & ~x7) | (x3 & n1927) | (~x7 & n1927);
  assign n3096 = x2 & ~n1927;
  assign n3097 = (x8 & ~n1927) | (x8 & n3096) | (~n1927 & n3096);
  assign n3098 = n3095 & ~n3097;
  assign n3099 = x6 | n3098;
  assign n3093 = x7 | n1696;
  assign n3094 = (~x2 & n1696) | (~x2 & n3093) | (n1696 & n3093);
  assign n3100 = x3 & ~n3094;
  assign n3101 = x6 & ~n3100;
  assign n3102 = n3099 & ~n3101;
  assign n3103 = x4 & n3102;
  assign n3104 = x6 & n260;
  assign n3105 = n60 & n3104;
  assign n3126 = n3103 | n3105;
  assign n3127 = x5 & n3126;
  assign n3128 = n3125 | n3127;
  assign n3130 = (x0 & x1) | (x0 & ~n3128) | (x1 & ~n3128);
  assign n3131 = n3129 & ~n3130;
  assign n3132 = (~x6 & x7) | (~x6 & n2998) | (x7 & n2998);
  assign n3133 = (x2 & x4) | (x2 & n3132) | (x4 & n3132);
  assign n3134 = n2998 & ~n3133;
  assign n3135 = (n3132 & ~n3133) | (n3132 & n3134) | (~n3133 & n3134);
  assign n3136 = (x3 & n1522) | (x3 & n3135) | (n1522 & n3135);
  assign n3137 = n3135 & ~n3136;
  assign n3138 = (x3 & x4) | (x3 & x6) | (x4 & x6);
  assign n3139 = (x3 & x8) | (x3 & ~n3138) | (x8 & ~n3138);
  assign n3140 = (~x6 & x8) | (~x6 & n3138) | (x8 & n3138);
  assign n3141 = ~n3139 & n3140;
  assign n3142 = x2 & ~n3141;
  assign n3143 = ~x3 & n1416;
  assign n3144 = x2 | n3143;
  assign n3145 = ~n3142 & n3144;
  assign n3149 = (~x1 & x7) | (~x1 & n3145) | (x7 & n3145);
  assign n3146 = ~x4 & n10;
  assign n3147 = (x2 & x3) | (x2 & n3146) | (x3 & n3146);
  assign n3148 = ~x2 & n3147;
  assign n3150 = x1 & n3148;
  assign n3151 = (n3145 & ~n3149) | (n3145 & n3150) | (~n3149 & n3150);
  assign n3152 = n10 & n46;
  assign n3153 = (x4 & x6) | (x4 & n3152) | (x6 & n3152);
  assign n3154 = ~x6 & n3153;
  assign n3155 = (~n3137 & n3151) | (~n3137 & n3154) | (n3151 & n3154);
  assign n3156 = x0 & ~n3154;
  assign n3157 = (n3137 & n3155) | (n3137 & ~n3156) | (n3155 & ~n3156);
  assign n3159 = n3131 | n3157;
  assign n3160 = (n3058 & ~n3158) | (n3058 & n3159) | (~n3158 & n3159);
  assign n3161 = n3031 | n3160;
  assign n3162 = (~n2974 & n3045) | (~n2974 & n3161) | (n3045 & n3161);
  assign n3163 = n2974 | n3162;
  assign n3173 = ~x5 & n530;
  assign n3174 = (x2 & ~x3) | (x2 & n3173) | (~x3 & n3173);
  assign n3175 = (n530 & n3173) | (n530 & n3174) | (n3173 & n3174);
  assign n3179 = x1 & n3175;
  assign n3176 = (~x2 & x4) | (~x2 & n1448) | (x4 & n1448);
  assign n3177 = (x2 & x5) | (x2 & ~n3176) | (x5 & ~n3176);
  assign n3178 = (n53 & n1448) | (n53 & ~n3177) | (n1448 & ~n3177);
  assign n3180 = x1 | n3178;
  assign n3181 = (~x1 & n3179) | (~x1 & n3180) | (n3179 & n3180);
  assign n3182 = x8 & ~n3181;
  assign n3169 = x1 | x5;
  assign n3170 = (x3 & x5) | (x3 & ~n3169) | (x5 & ~n3169);
  assign n3171 = (x2 & x3) | (x2 & ~n3169) | (x3 & ~n3169);
  assign n3172 = (n178 & n3170) | (n178 & ~n3171) | (n3170 & ~n3171);
  assign n3183 = ~x4 & n3172;
  assign n3184 = x8 | n3183;
  assign n3185 = ~n3182 & n3184;
  assign n3186 = (x0 & ~n2247) | (x0 & n3185) | (~n2247 & n3185);
  assign n3164 = x4 & n2541;
  assign n3165 = (~x3 & x4) | (~x3 & n2541) | (x4 & n2541);
  assign n3166 = (x3 & ~n3164) | (x3 & n3165) | (~n3164 & n3165);
  assign n3167 = x1 | n3166;
  assign n3168 = x2 | n3167;
  assign n3187 = (x0 & n2247) | (x0 & n3168) | (n2247 & n3168);
  assign n3188 = n3186 & ~n3187;
  assign n3203 = (x1 & n750) | (x1 & n812) | (n750 & n812);
  assign n3204 = ~n750 & n3203;
  assign n3205 = ~x3 & n1839;
  assign n3206 = (x1 & x2) | (x1 & n3205) | (x2 & n3205);
  assign n3207 = ~x1 & n3206;
  assign n3208 = n318 & ~n337;
  assign n3209 = n20 & n3208;
  assign n3210 = (~n3204 & n3207) | (~n3204 & n3209) | (n3207 & n3209);
  assign n3211 = x0 & ~n3209;
  assign n3212 = (n3204 & n3210) | (n3204 & ~n3211) | (n3210 & ~n3211);
  assign n3294 = n738 & n3212;
  assign n3213 = (~n46 & n118) | (~n46 & n2287) | (n118 & n2287);
  assign n3214 = n46 & n3213;
  assign n3279 = (x2 & x6) | (x2 & x7) | (x6 & x7);
  assign n3280 = (x2 & x8) | (x2 & ~n3279) | (x8 & ~n3279);
  assign n3281 = (~x7 & x8) | (~x7 & n3279) | (x8 & n3279);
  assign n3282 = ~n3280 & n3281;
  assign n3283 = x1 | n3282;
  assign n3284 = x2 & n571;
  assign n3285 = x1 & ~n3284;
  assign n3286 = n3283 & ~n3285;
  assign n3287 = x4 & n3286;
  assign n3277 = (x6 & n29) | (x6 & ~n519) | (n29 & ~n519);
  assign n3278 = n29 & ~n3277;
  assign n3288 = n3278 | n3287;
  assign n3289 = (x1 & n3287) | (x1 & n3288) | (n3287 & n3288);
  assign n3290 = ~n1415 & n3289;
  assign n3234 = x5 & ~n1017;
  assign n3235 = (~x3 & x4) | (~x3 & n3234) | (x4 & n3234);
  assign n3236 = (~n1017 & n3234) | (~n1017 & n3235) | (n3234 & n3235);
  assign n3240 = x7 & n3236;
  assign n3237 = (x3 & ~x4) | (x3 & n153) | (~x4 & n153);
  assign n3238 = (~x5 & n20) | (~x5 & n3237) | (n20 & n3237);
  assign n3239 = (x5 & ~n1595) | (x5 & n3238) | (~n1595 & n3238);
  assign n3241 = ~x7 & n3239;
  assign n3242 = (x7 & ~n3240) | (x7 & n3241) | (~n3240 & n3241);
  assign n3243 = x2 | n3242;
  assign n3231 = ~x5 & n184;
  assign n3232 = n80 & n3231;
  assign n3233 = n20 & n231;
  assign n3244 = n3232 | n3233;
  assign n3245 = x2 & n3244;
  assign n3246 = n3243 & ~n3245;
  assign n3247 = (x1 & ~x6) | (x1 & n3246) | (~x6 & n3246);
  assign n3228 = n21 & ~n231;
  assign n3215 = (x3 & x8) | (x3 & n500) | (x8 & n500);
  assign n3216 = (x7 & x8) | (x7 & ~n3215) | (x8 & ~n3215);
  assign n3217 = n500 & n3216;
  assign n3218 = (x3 & ~n3215) | (x3 & n3217) | (~n3215 & n3217);
  assign n3221 = (x4 & x5) | (x4 & n3218) | (x5 & n3218);
  assign n3219 = (x3 & ~n29) | (x3 & n147) | (~n29 & n147);
  assign n3220 = n29 & n3219;
  assign n3222 = ~x5 & n3220;
  assign n3223 = (n3218 & ~n3221) | (n3218 & n3222) | (~n3221 & n3222);
  assign n3224 = x2 & ~n42;
  assign n3225 = n271 & n3224;
  assign n3226 = (n11 & ~n42) | (n11 & n3224) | (~n42 & n3224);
  assign n3227 = (x3 & n3225) | (x3 & n3226) | (n3225 & n3226);
  assign n3229 = n3223 | n3227;
  assign n3230 = (n21 & ~n3228) | (n21 & n3229) | (~n3228 & n3229);
  assign n3248 = (x1 & x6) | (x1 & n3230) | (x6 & n3230);
  assign n3249 = ~n3247 & n3248;
  assign n3253 = x1 & ~n241;
  assign n3254 = x1 | n330;
  assign n3255 = ~n3253 & n3254;
  assign n3256 = x4 & ~n3255;
  assign n3250 = (x3 & x5) | (x3 & n227) | (x5 & n227);
  assign n3251 = n225 & ~n3250;
  assign n3252 = (n227 & ~n3250) | (n227 & n3251) | (~n3250 & n3251);
  assign n3257 = ~x1 & n3252;
  assign n3258 = x4 | n3257;
  assign n3259 = ~n3256 & n3258;
  assign n3274 = (x2 & ~x6) | (x2 & n3259) | (~x6 & n3259);
  assign n3262 = (x4 & ~x8) | (x4 & n547) | (~x8 & n547);
  assign n3263 = x4 & ~n3262;
  assign n3264 = n3262 | n3263;
  assign n3265 = (~x4 & n3263) | (~x4 & n3264) | (n3263 & n3264);
  assign n3266 = x1 & ~n3265;
  assign n3267 = ~x4 & n213;
  assign n3268 = x1 | n3267;
  assign n3269 = ~n3266 & n3268;
  assign n3270 = x3 | n3269;
  assign n3260 = (~x1 & x4) | (~x1 & x8) | (x4 & x8);
  assign n3261 = n2678 & n3260;
  assign n3271 = ~x5 & n3261;
  assign n3272 = x3 & ~n3271;
  assign n3273 = n3270 & ~n3272;
  assign n3275 = (x2 & x6) | (x2 & ~n3273) | (x6 & ~n3273);
  assign n3276 = n3274 & ~n3275;
  assign n3291 = (~x0 & n3249) | (~x0 & n3276) | (n3249 & n3276);
  assign n3292 = ~n3290 & n3291;
  assign n3293 = (~x0 & n3290) | (~x0 & n3292) | (n3290 & n3292);
  assign n3295 = n3214 | n3293;
  assign n3296 = (n3212 & ~n3294) | (n3212 & n3295) | (~n3294 & n3295);
  assign n3193 = (x1 & ~n45) | (x1 & n1369) | (~n45 & n1369);
  assign n3194 = ~x1 & n3193;
  assign n3189 = (~x3 & x5) | (~x3 & n1709) | (x5 & n1709);
  assign n3190 = (x1 & ~x5) | (x1 & n1709) | (~x5 & n1709);
  assign n3191 = (x3 & ~x6) | (x3 & n3190) | (~x6 & n3190);
  assign n3192 = n3189 | n3191;
  assign n3195 = (x2 & ~n3192) | (x2 & n3194) | (~n3192 & n3194);
  assign n3196 = x4 & ~n3195;
  assign n3197 = (x4 & n3194) | (x4 & ~n3196) | (n3194 & ~n3196);
  assign n3200 = (x0 & n29) | (x0 & n3197) | (n29 & n3197);
  assign n3198 = (x5 & x6) | (x5 & n319) | (x6 & n319);
  assign n3199 = ~x6 & n3198;
  assign n3201 = ~n29 & n3199;
  assign n3202 = (n3197 & ~n3200) | (n3197 & n3201) | (~n3200 & n3201);
  assign n3323 = (~x4 & x7) | (~x4 & x8) | (x7 & x8);
  assign n3324 = (x0 & x8) | (x0 & ~n3323) | (x8 & ~n3323);
  assign n3325 = (x4 & ~x7) | (x4 & n3324) | (~x7 & n3324);
  assign n3326 = n3323 & n3325;
  assign n3327 = (~n3324 & n3325) | (~n3324 & n3326) | (n3325 & n3326);
  assign n3328 = x1 | n3327;
  assign n3321 = x4 & ~n266;
  assign n3322 = (x7 & ~n266) | (x7 & n3321) | (~n266 & n3321);
  assign n3329 = ~x0 & n3322;
  assign n3330 = x1 & ~n3329;
  assign n3331 = n3328 & ~n3330;
  assign n3332 = x2 | n3331;
  assign n3318 = (x4 & x7) | (x4 & ~x8) | (x7 & ~x8);
  assign n3319 = (~x1 & x7) | (~x1 & x8) | (x7 & x8);
  assign n3320 = n3318 | n3319;
  assign n3333 = x0 | n3320;
  assign n3334 = x2 & n3333;
  assign n3335 = n3332 & ~n3334;
  assign n3336 = x3 | n3335;
  assign n3310 = (x4 & x7) | (x4 & ~n1336) | (x7 & ~n1336);
  assign n3311 = (x1 & x2) | (x1 & ~n3310) | (x2 & ~n3310);
  assign n3312 = ~n1336 & n3311;
  assign n3313 = (n3310 & n3311) | (n3310 & n3312) | (n3311 & n3312);
  assign n3314 = x4 & n184;
  assign n3315 = ~n15 & n3314;
  assign n3316 = x8 & ~n3315;
  assign n3317 = (n3313 & n3315) | (n3313 & ~n3316) | (n3315 & ~n3316);
  assign n3337 = ~x0 & n3317;
  assign n3338 = x3 & ~n3337;
  assign n3339 = n3336 & ~n3338;
  assign n3340 = x6 & n3339;
  assign n3297 = ~n28 & n80;
  assign n3298 = (x0 & x1) | (x0 & ~x4) | (x1 & ~x4);
  assign n3299 = x0 & ~n3298;
  assign n3300 = (x1 & ~x8) | (x1 & n3299) | (~x8 & n3299);
  assign n3301 = (~n3298 & n3299) | (~n3298 & n3300) | (n3299 & n3300);
  assign n3304 = (x3 & x7) | (x3 & n3301) | (x7 & n3301);
  assign n3302 = (x4 & n43) | (x4 & n1598) | (n43 & n1598);
  assign n3303 = ~x4 & n3302;
  assign n3305 = x7 & n3303;
  assign n3306 = (~x3 & n3304) | (~x3 & n3305) | (n3304 & n3305);
  assign n3307 = ~x2 & n3306;
  assign n3308 = n40 | n3307;
  assign n3309 = (n3297 & n3307) | (n3297 & n3308) | (n3307 & n3308);
  assign n3341 = x6 | n3309;
  assign n3342 = (~x6 & n3340) | (~x6 & n3341) | (n3340 & n3341);
  assign n3343 = n3202 | n3342;
  assign n3344 = (~n3188 & n3296) | (~n3188 & n3343) | (n3296 & n3343);
  assign n3345 = n3188 | n3344;
  assign n3350 = x0 & ~x2;
  assign n3351 = (~x0 & x2) | (~x0 & n1668) | (x2 & n1668);
  assign n3352 = x1 & n1668;
  assign n3353 = (n3350 & n3351) | (n3350 & ~n3352) | (n3351 & ~n3352);
  assign n3354 = ~x8 & n3353;
  assign n3349 = n1233 & n1668;
  assign n3355 = n3349 | n3354;
  assign n3356 = (~x0 & n3354) | (~x0 & n3355) | (n3354 & n3355);
  assign n3357 = x3 | n3356;
  assign n3346 = ~x8 & n1233;
  assign n3347 = (x1 & ~x2) | (x1 & n3346) | (~x2 & n3346);
  assign n3348 = (n1233 & n3346) | (n1233 & n3347) | (n3346 & n3347);
  assign n3358 = ~x0 & n3348;
  assign n3359 = x3 & ~n3358;
  assign n3360 = n3357 & ~n3359;
  assign n3484 = n750 & n3360;
  assign n3363 = (x8 & n1392) | (x8 & ~n2131) | (n1392 & ~n2131);
  assign n3364 = x2 & ~n3363;
  assign n3361 = x3 & ~n2978;
  assign n3362 = n2851 & ~n3361;
  assign n3365 = x2 | n3362;
  assign n3366 = (~x2 & n3364) | (~x2 & n3365) | (n3364 & n3365);
  assign n3367 = x0 | n3366;
  assign n3368 = x1 | n45;
  assign n3369 = x0 & n3368;
  assign n3370 = n3367 & ~n3369;
  assign n3371 = (x5 & x7) | (x5 & n3370) | (x7 & n3370);
  assign n3372 = (x4 & ~x5) | (x4 & n3371) | (~x5 & n3371);
  assign n3373 = (x4 & x7) | (x4 & ~n3371) | (x7 & ~n3371);
  assign n3374 = n3372 & ~n3373;
  assign n3375 = ~x6 & n184;
  assign n3376 = n61 & n3375;
  assign n3481 = n46 & ~n3376;
  assign n3411 = (x1 & x6) | (x1 & n129) | (x6 & n129);
  assign n3412 = (x6 & x7) | (x6 & ~n3411) | (x7 & ~n3411);
  assign n3413 = (x1 & ~x5) | (x1 & n3412) | (~x5 & n3412);
  assign n3414 = ~n3411 & n3413;
  assign n3415 = x3 | n3414;
  assign n3416 = x1 & n553;
  assign n3417 = x3 & ~n3416;
  assign n3418 = n3415 & ~n3417;
  assign n3419 = x2 & n3418;
  assign n3399 = (x3 & x6) | (x3 & n129) | (x6 & n129);
  assign n3400 = (x5 & ~x6) | (x5 & n129) | (~x6 & n129);
  assign n3401 = (x3 & x7) | (x3 & ~n3400) | (x7 & ~n3400);
  assign n3402 = ~n3399 & n3401;
  assign n3403 = x1 | n3402;
  assign n3404 = ~x3 & n860;
  assign n3405 = x1 & ~n3404;
  assign n3406 = n3403 & ~n3405;
  assign n3407 = (x1 & ~x3) | (x1 & n583) | (~x3 & n583);
  assign n3408 = (x3 & ~x6) | (x3 & n583) | (~x6 & n583);
  assign n3409 = (x1 & x7) | (x1 & ~n3408) | (x7 & ~n3408);
  assign n3410 = ~n3407 & n3409;
  assign n3420 = n3406 | n3410;
  assign n3421 = ~x2 & n3420;
  assign n3422 = n3419 | n3421;
  assign n3423 = ~x4 & n3422;
  assign n3377 = ~x7 & n1881;
  assign n3378 = (x1 & x2) | (x1 & ~n1881) | (x2 & ~n1881);
  assign n3379 = (x7 & n39) | (x7 & ~n3378) | (n39 & ~n3378);
  assign n3380 = (x7 & n3377) | (x7 & ~n3379) | (n3377 & ~n3379);
  assign n3383 = (x3 & x6) | (x3 & n3380) | (x6 & n3380);
  assign n3381 = (x5 & ~n39) | (x5 & n1803) | (~n39 & n1803);
  assign n3382 = n39 & n3381;
  assign n3384 = ~x6 & n3382;
  assign n3385 = (n3380 & ~n3383) | (n3380 & n3384) | (~n3383 & n3384);
  assign n3386 = (x1 & ~x2) | (x1 & x7) | (~x2 & x7);
  assign n3387 = (x3 & ~x7) | (x3 & n3386) | (~x7 & n3386);
  assign n3388 = (x1 & ~x2) | (x1 & n3387) | (~x2 & n3387);
  assign n3389 = ~n3386 & n3388;
  assign n3390 = (~n3387 & n3388) | (~n3387 & n3389) | (n3388 & n3389);
  assign n3396 = (x5 & x6) | (x5 & ~n3390) | (x6 & ~n3390);
  assign n3391 = (x2 & ~x3) | (x2 & x5) | (~x3 & x5);
  assign n3392 = (~x5 & x7) | (~x5 & n3391) | (x7 & n3391);
  assign n3393 = (x2 & ~x3) | (x2 & n3392) | (~x3 & n3392);
  assign n3394 = ~n3391 & n3393;
  assign n3395 = (~n3392 & n3393) | (~n3392 & n3394) | (n3393 & n3394);
  assign n3397 = x6 & n3395;
  assign n3398 = (n3390 & n3396) | (n3390 & n3397) | (n3396 & n3397);
  assign n3424 = n3385 | n3398;
  assign n3425 = x4 & n3424;
  assign n3426 = n3423 | n3425;
  assign n3430 = (x0 & ~x8) | (x0 & n3426) | (~x8 & n3426);
  assign n3427 = n15 | n632;
  assign n3428 = (n10 & n36) | (n10 & n3427) | (n36 & n3427);
  assign n3429 = n10 & ~n3428;
  assign n3431 = ~x0 & n3429;
  assign n3432 = (n3426 & ~n3430) | (n3426 & n3431) | (~n3430 & n3431);
  assign n3444 = (x4 & ~n39) | (x4 & n1437) | (~n39 & n1437);
  assign n3445 = n39 & n3444;
  assign n3447 = ~x8 & n3445;
  assign n3454 = (x1 & x2) | (x1 & ~x6) | (x2 & ~x6);
  assign n3455 = (~x2 & x6) | (~x2 & n3454) | (x6 & n3454);
  assign n3456 = (x2 & x4) | (x2 & ~n3455) | (x4 & ~n3455);
  assign n3457 = (n338 & n3454) | (n338 & ~n3456) | (n3454 & ~n3456);
  assign n3458 = (x3 & x8) | (x3 & n3457) | (x8 & n3457);
  assign n3459 = (n3447 & n3457) | (n3447 & ~n3458) | (n3457 & ~n3458);
  assign n3460 = ~x5 & n3459;
  assign n3440 = x4 & n1392;
  assign n3441 = (~x1 & x4) | (~x1 & n1437) | (x4 & n1437);
  assign n3442 = x1 & ~n1437;
  assign n3443 = (~n3440 & n3441) | (~n3440 & n3442) | (n3441 & n3442);
  assign n3446 = (x2 & x8) | (x2 & ~n3443) | (x8 & ~n3443);
  assign n3448 = (n3443 & n3446) | (n3443 & ~n3447) | (n3446 & ~n3447);
  assign n3449 = (n311 & n684) | (n311 & ~n2374) | (n684 & ~n2374);
  assign n3450 = (x1 & x4) | (x1 & ~n3449) | (x4 & ~n3449);
  assign n3451 = (x3 & ~x4) | (x3 & n3450) | (~x4 & n3450);
  assign n3452 = (x1 & x3) | (x1 & ~n3450) | (x3 & ~n3450);
  assign n3453 = n3451 & ~n3452;
  assign n3461 = n3448 & ~n3453;
  assign n3462 = x5 & ~n3461;
  assign n3463 = n3460 | n3462;
  assign n3433 = x1 | x6;
  assign n3434 = (n61 & n573) | (n61 & n3433) | (n573 & n3433);
  assign n3435 = (~x4 & n61) | (~x4 & n3434) | (n61 & n3434);
  assign n3436 = ~x4 & n1541;
  assign n3437 = x1 & n3436;
  assign n3438 = x8 | n3437;
  assign n3439 = (n3435 & n3437) | (n3435 & n3438) | (n3437 & n3438);
  assign n3464 = (x2 & x3) | (x2 & n3439) | (x3 & n3439);
  assign n3465 = (~n42 & n3463) | (~n42 & n3464) | (n3463 & n3464);
  assign n3467 = (x1 & x2) | (x1 & x6) | (x2 & x6);
  assign n3468 = (x1 & x3) | (x1 & ~n3467) | (x3 & ~n3467);
  assign n3469 = (~x2 & x3) | (~x2 & n3467) | (x3 & n3467);
  assign n3470 = ~n3468 & n3469;
  assign n3471 = x0 | n3470;
  assign n3466 = x3 | n1287;
  assign n3472 = x1 | n3466;
  assign n3473 = x0 & n3472;
  assign n3474 = n3471 & ~n3473;
  assign n3475 = (x4 & x8) | (x4 & n3474) | (x8 & n3474);
  assign n3476 = (x5 & ~x8) | (x5 & n3475) | (~x8 & n3475);
  assign n3477 = (x4 & x5) | (x4 & ~n3475) | (x5 & ~n3475);
  assign n3478 = n3476 & ~n3477;
  assign n3479 = x0 & ~n3478;
  assign n3480 = (n3465 & n3478) | (n3465 & ~n3479) | (n3478 & ~n3479);
  assign n3482 = n3432 | n3480;
  assign n3483 = (n46 & ~n3481) | (n46 & n3482) | (~n3481 & n3482);
  assign n3485 = n3374 | n3483;
  assign n3486 = (n3360 & ~n3484) | (n3360 & n3485) | (~n3484 & n3485);
  assign y0 = n35;
  assign y1 = n110;
  assign y2 = n212;
  assign y3 = n329;
  assign y4 = n518;
  assign y5 = n737;
  assign y6 = n919;
  assign y7 = n1094;
  assign y8 = n1286;
  assign y9 = n1479;
  assign y10 = n1665;
  assign y11 = n1855;
  assign y12 = n2045;
  assign y13 = n2211;
  assign y14 = n2409;
  assign y15 = n2578;
  assign y16 = n2774;
  assign y17 = n2968;
  assign y18 = n3163;
  assign y19 = n3345;
  assign y20 = n3486;
endmodule
