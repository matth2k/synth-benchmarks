module s420 (
  CK,
  C_0,
  C_1,
  C_10,
  C_11,
  C_12,
  C_13,
  C_14,
  C_15,
  C_16,
  C_2,
  C_3,
  C_4,
  C_5,
  C_6,
  C_7,
  C_8,
  C_9,
  P_0,
  Z
);
  input CK;
  wire CK;
  input C_0;
  wire C_0;
  input C_1;
  wire C_1;
  input C_10;
  wire C_10;
  input C_11;
  wire C_11;
  input C_12;
  wire C_12;
  input C_13;
  wire C_13;
  input C_14;
  wire C_14;
  input C_15;
  wire C_15;
  input C_16;
  wire C_16;
  input C_2;
  wire C_2;
  input C_3;
  wire C_3;
  input C_4;
  wire C_4;
  input C_5;
  wire C_5;
  input C_6;
  wire C_6;
  input C_7;
  wire C_7;
  input C_8;
  wire C_8;
  input C_9;
  wire C_9;
  input P_0;
  wire P_0;
  output Z;
  wire Z;
  wire __0__;
  wire __1__;
  wire __2__;
  wire __3__;
  wire __4__;
  wire __5__;
  wire __6__;
  wire __7__;
  wire __8__;
  wire __9__;
  wire __10__;
  wire __11__;
  wire __12__;
  wire __13__;
  wire __14__;
  wire __15__;
  wire __17__;
  wire __18__;
  wire __19__;
  wire __21__;
  wire __22__;
  wire __23__;
  wire __24__;
  wire __25__;
  wire __26__;
  wire __27__;
  wire __28__;
  wire __29__;
  wire __30__;
  wire __31__;
  wire __32__;
  wire __33__;
  wire __34__;
  wire __35__;
  wire __36__;
  wire __37__;
  wire __38__;
  wire __39__;
  wire __40__;
  wire __41__;
  wire __42__;
  wire __43__;
  wire __44__;
  wire __45__;
  wire __46__;
  wire __47__;
  wire __48__;
  wire __49__;
  wire __50__;
  wire __51__;
  wire __52__;
  wire __53__;
  wire __54__;
  FDRE #(
    .INIT(1'bx)
  ) __55__ (
    .D(__19__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__0__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __56__ (
    .D(__17__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __57__ (
    .D(__18__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__2__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __58__ (
    .D(__53__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__3__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __59__ (
    .D(__47__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__4__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __60__ (
    .D(__45__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__5__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __61__ (
    .D(__52__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__6__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __62__ (
    .D(__51__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__7__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __63__ (
    .D(__54__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__8__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __64__ (
    .D(__48__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__9__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __65__ (
    .D(__50__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__10__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __66__ (
    .D(__46__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__11__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __67__ (
    .D(__44__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__12__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __68__ (
    .D(__42__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__13__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __69__ (
    .D(__41__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__14__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __70__ (
    .D(__49__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__15__)
  );
  LUT4 #(
    .INIT(16'h7f80)
  ) __72__ (
    .I3(__1__),
    .I2(P_0),
    .I1(__3__),
    .I0(__0__),
    .O(__17__)
  );
  LUT5 #(
    .INIT(32'h7fff8000)
  ) __73__ (
    .I4(__2__),
    .I3(P_0),
    .I2(__3__),
    .I1(__0__),
    .I0(__1__),
    .O(__18__)
  );
  LUT3 #(
    .INIT(8'h78)
  ) __74__ (
    .I2(__0__),
    .I1(P_0),
    .I0(__3__),
    .O(__19__)
  );
  LUT4 #(
    .INIT(16'h0001)
  ) __76__ (
    .I3(__4__),
    .I2(__6__),
    .I1(__5__),
    .I0(__7__),
    .O(__21__)
  );
  LUT4 #(
    .INIT(16'h0001)
  ) __77__ (
    .I3(__8__),
    .I2(__9__),
    .I1(__11__),
    .I0(__10__),
    .O(__22__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __78__ (
    .I1(__13__),
    .I0(C_15),
    .O(__23__)
  );
  LUT6 #(
    .INIT(64'h0f0f5533ffffffff)
  ) __79__ (
    .I5(P_0),
    .I4(__15__),
    .I3(__14__),
    .I2(C_13),
    .I1(__23__),
    .I0(C_14),
    .O(__24__)
  );
  LUT3 #(
    .INIT(8'h07)
  ) __80__ (
    .I2(__9__),
    .I1(__8__),
    .I0(C_12),
    .O(__25__)
  );
  LUT6 #(
    .INIT(64'h00000f0f0000ff44)
  ) __81__ (
    .I5(__10__),
    .I4(__11__),
    .I3(__25__),
    .I2(C_10),
    .I1(__9__),
    .I0(C_11),
    .O(__26__)
  );
  LUT6 #(
    .INIT(64'hff0f4404ff0fff0f)
  ) __82__ (
    .I5(P_0),
    .I4(__26__),
    .I3(__24__),
    .I2(__22__),
    .I1(__11__),
    .I0(C_9),
    .O(__27__)
  );
  LUT4 #(
    .INIT(16'h0001)
  ) __83__ (
    .I3(__2__),
    .I2(__3__),
    .I1(__0__),
    .I0(__1__),
    .O(__28__)
  );
  LUT5 #(
    .INIT(32'h00f00088)
  ) __84__ (
    .I4(__5__),
    .I3(__6__),
    .I2(C_7),
    .I1(__4__),
    .I0(C_8),
    .O(__29__)
  );
  LUT6 #(
    .INIT(64'hf0f0ff8800000000)
  ) __85__ (
    .I5(P_0),
    .I4(__7__),
    .I3(__29__),
    .I2(C_5),
    .I1(__6__),
    .I0(C_6),
    .O(__30__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __86__ (
    .I1(P_0),
    .I0(__15__),
    .O(__31__)
  );
  LUT3 #(
    .INIT(8'h08)
  ) __87__ (
    .I2(__13__),
    .I1(__12__),
    .I0(C_16),
    .O(__32__)
  );
  LUT6 #(
    .INIT(64'h4000000000000000)
  ) __88__ (
    .I5(__28__),
    .I4(__32__),
    .I3(__31__),
    .I2(__22__),
    .I1(__21__),
    .I0(__14__),
    .O(__33__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __89__ (
    .I1(__2__),
    .I0(C_4),
    .O(__34__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __90__ (
    .I1(P_0),
    .I0(__3__),
    .O(__35__)
  );
  LUT6 #(
    .INIT(64'hf0f0aacc00000000)
  ) __91__ (
    .I5(__35__),
    .I4(__0__),
    .I3(__1__),
    .I2(C_2),
    .I1(__34__),
    .I0(C_3),
    .O(__36__)
  );
  LUT5 #(
    .INIT(32'h00000f7f)
  ) __92__ (
    .I4(__36__),
    .I3(C_0),
    .I2(P_0),
    .I1(__3__),
    .I0(C_1),
    .O(__37__)
  );
  LUT6 #(
    .INIT(64'hfffff020ffffffff)
  ) __93__ (
    .I5(__37__),
    .I4(__33__),
    .I3(__30__),
    .I2(__28__),
    .I1(__27__),
    .I0(__21__),
    .O(__38__)
  );
  LUT6 #(
    .INIT(64'h8000000000000000)
  ) __94__ (
    .I5(__7__),
    .I4(__2__),
    .I3(P_0),
    .I2(__3__),
    .I1(__0__),
    .I0(__1__),
    .O(__39__)
  );
  LUT6 #(
    .INIT(64'h8000000000000000)
  ) __95__ (
    .I5(__11__),
    .I4(__10__),
    .I3(__4__),
    .I2(__6__),
    .I1(__5__),
    .I0(__39__),
    .O(__40__)
  );
  LUT5 #(
    .INIT(32'h7fff8000)
  ) __96__ (
    .I4(__14__),
    .I3(__8__),
    .I2(__9__),
    .I1(__40__),
    .I0(__15__),
    .O(__41__)
  );
  LUT6 #(
    .INIT(64'h7fffffff80000000)
  ) __97__ (
    .I5(__13__),
    .I4(__8__),
    .I3(__9__),
    .I2(__40__),
    .I1(__15__),
    .I0(__14__),
    .O(__42__)
  );
  LUT6 #(
    .INIT(64'h8000000000000000)
  ) __98__ (
    .I5(__8__),
    .I4(__9__),
    .I3(__40__),
    .I2(__15__),
    .I1(__13__),
    .I0(__14__),
    .O(__43__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __99__ (
    .I1(__12__),
    .I0(__43__),
    .O(__44__)
  );
  LUT3 #(
    .INIT(8'h78)
  ) __100__ (
    .I2(__5__),
    .I1(__6__),
    .I0(__39__),
    .O(__45__)
  );
  LUT5 #(
    .INIT(32'h7fff8000)
  ) __101__ (
    .I4(__11__),
    .I3(__4__),
    .I2(__6__),
    .I1(__5__),
    .I0(__39__),
    .O(__46__)
  );
  LUT4 #(
    .INIT(16'h7f80)
  ) __102__ (
    .I3(__4__),
    .I2(__6__),
    .I1(__5__),
    .I0(__39__),
    .O(__47__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __103__ (
    .I1(__9__),
    .I0(__40__),
    .O(__48__)
  );
  LUT4 #(
    .INIT(16'h7f80)
  ) __104__ (
    .I3(__15__),
    .I2(__8__),
    .I1(__9__),
    .I0(__40__),
    .O(__49__)
  );
  LUT6 #(
    .INIT(64'h7fffffff80000000)
  ) __105__ (
    .I5(__10__),
    .I4(__11__),
    .I3(__4__),
    .I2(__6__),
    .I1(__5__),
    .I0(__39__),
    .O(__50__)
  );
  LUT6 #(
    .INIT(64'h7fffffff80000000)
  ) __106__ (
    .I5(__7__),
    .I4(__2__),
    .I3(P_0),
    .I2(__3__),
    .I1(__0__),
    .I0(__1__),
    .O(__51__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __107__ (
    .I1(__6__),
    .I0(__39__),
    .O(__52__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __108__ (
    .I1(P_0),
    .I0(__3__),
    .O(__53__)
  );
  LUT3 #(
    .INIT(8'h78)
  ) __109__ (
    .I2(__8__),
    .I1(__9__),
    .I0(__40__),
    .O(__54__)
  );
  assign Z = __38__;
endmodule
