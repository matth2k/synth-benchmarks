// IWLS benchmark module "b9" printed on Wed May 29 16:27:40 2002
module b9(a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, \xx , y, z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0, o0, p0, q0, r0, s0, t0, u0, v0, w0, x0, y0, z0, a1, b1, c1, d1, e1, f1, g1, h1, i1, j1);
input
  a,
  b,
  c,
  d,
  e,
  f,
  g,
  h,
  i,
  j,
  k,
  l,
  m,
  n,
  o,
  p,
  q,
  r,
  s,
  t,
  u,
  v,
  w,
  \xx ,
  y,
  z,
  a0,
  b0,
  c0,
  d0,
  e0,
  f0,
  g0,
  h0,
  i0,
  j0,
  k0,
  l0,
  m0,
  n0,
  o0;
output
  a1,
  b1,
  c1,
  d1,
  e1,
  f1,
  g1,
  h1,
  i1,
  j1,
  p0,
  q0,
  r0,
  s0,
  t0,
  u0,
  v0,
  w0,
  x0,
  y0,
  z0;
wire
  \[15] ,
  \[16] ,
  \[17] ,
  \[18] ,
  \[19] ,
  \[0] ,
  \[1] ,
  \[20] ,
  \[2] ,
  \[3] ,
  \[4] ,
  \[5] ,
  \[6] ,
  \[7] ,
  \[8] ,
  \[9] ,
  a3,
  a4,
  a5,
  b3,
  b4,
  b5,
  c3,
  c4,
  c5,
  d3,
  d4,
  d5,
  e3,
  e4,
  e5,
  f2,
  f3,
  f4,
  f5,
  g2,
  g3,
  g4,
  g5,
  h2,
  h3,
  h4,
  h5,
  i2,
  i3,
  i4,
  i5,
  j2,
  j3,
  j4,
  j5,
  k2,
  k3,
  k4,
  k5,
  l2,
  l3,
  l4,
  l5,
  m2,
  m3,
  m4,
  m5,
  n2,
  n3,
  n4,
  n5,
  o2,
  o3,
  o4,
  o5,
  p2,
  p3,
  p4,
  p5,
  q2,
  q3,
  q4,
  q5,
  r2,
  r3,
  r4,
  r5,
  s2,
  s3,
  s4,
  s5,
  t2,
  t3,
  t4,
  t5,
  u2,
  u3,
  u4,
  u5,
  v2,
  v3,
  v4,
  v5,
  w2,
  w3,
  w4,
  w5,
  x2,
  x3,
  x4,
  y2,
  y3,
  y4,
  z2,
  z3,
  z4,
  \[10] ,
  \[11] ,
  \[12] ,
  \[13] ,
  \[14] ;
assign
  \[15]  = ~i3,
  \[16]  = ~d4,
  \[17]  = ~e4,
  \[18]  = ~\[11] ,
  \[19]  = ~\[18] ,
  \[0]  = (~p & ~o2) | ~q,
  \[1]  = ~z3,
  \[20]  = (~t2 & ~s2) | (~n0 & ~s2),
  \[2]  = ~o0 | (~n0 | ~l3),
  \[3]  = ~f3,
  \[4]  = ~g3,
  \[5]  = ~\[6] ,
  \[6]  = ~j4,
  \[7]  = (~m0 & ~u2) | (~v2 & ~u2),
  \[8]  = ~a5,
  \[9]  = ~x2,
  a1 = \[11] ,
  a3 = ~o0,
  a4 = ~j0,
  a5 = ~n0 | ~o0,
  b1 = \[12] ,
  b3 = ~\xx ,
  b4 = ~g0,
  b5 = ~n4 | ~u3,
  c1 = \[13] ,
  c3 = ~y,
  c4 = ~e,
  c5 = ~o0 | ~c4,
  d1 = \[14] ,
  d3 = ~v,
  d4 = ~b | (~w | ~b3),
  d5 = (~t5 & ~b5) | (~b0 & ~b5),
  e1 = \[15] ,
  e3 = ~o0,
  e4 = ~b | (~w | (~\xx  | ~c3)),
  e5 = ~d5 & (~c5 & ~n),
  f1 = \[16] ,
  f2 = ~o,
  f3 = ~d3 & ~k3,
  f4 = (~j0 & ~k0) | (~r3 & ~k0),
  f5 = ~w5,
  g1 = \[17] ,
  g2 = ~m2 | (~l2 | ~k2),
  g3 = ~k3 & ~v,
  g4 = ~f4,
  g5 = ~r3 | ~j0,
  h1 = \[18] ,
  h2 = ~j2 & ~i2,
  h3 = ~b0,
  h4 = ~g4 | (~b0 | (~c4 | ~h)),
  h5 = ~r,
  i1 = \[19] ,
  i2 = ~d0 | ~i,
  i3 = ~f5 | (~b0 | ~m),
  i4 = ~a3 & ~f4,
  i5 = ~l0 | (~g | ~b0),
  j1 = \[20] ,
  j2 = ~o0,
  j3 = ~a4 & ~r3,
  j4 = (~h3 & ~r3) | ~k4,
  j5 = ~f | (~m5 | (~c4 | ~n0)),
  k2 = ~e0 & ~j,
  k3 = (~j3 & ~l0) | ((~j3 & ~h3) | ((~b0 & ~l0) | (~b0 & ~h3))),
  k4 = ~l0,
  k5 = ~n5,
  l2 = ~c4 | (~b0 | (~r3 | ~j0)),
  l3 = ~m3,
  l4 = ~h5 & ~p,
  l5 = ~e0,
  m2 = ~n3 | ~h3,
  m3 = (~v5 & ~c4) | ~q3,
  m4 = ~h0 & (~f0 & ~l4),
  m5 = ~p5 | ~o5,
  n2 = ~\[12] ,
  n3 = ~c0 & (~y4 & ~a4),
  n4 = ~g0,
  n5 = (~n0 & ~h4) | (~o0 & ~h4),
  o2 = ~n2,
  o3 = ~d0 | ~i,
  o4 = ~k0,
  o5 = ~b0 | ~i4,
  p0 = \[0] ,
  p2 = ~j0,
  p3 = ~c,
  p4 = ~t,
  p5 = ~o0 | ~q5,
  q0 = \[1] ,
  q2 = ~p2 & ~r3,
  q3 = ~p3 | ~o3,
  q4 = ~s,
  q5 = ~b4 | ~l5,
  r0 = \[2] ,
  r2 = ~q2 & ~l0,
  r3 = ~c0,
  r4 = ~q4 | (~u | ~p4),
  r5 = (~j0 & ~l0) | (~c0 & ~l0),
  s0 = \[3] ,
  s2 = ~v3 | (~u3 | (~s3 | ~t3)),
  s3 = ~j0 | (~i | ~r3),
  s4 = (~v4 & ~x4) | (~b0 & ~x4),
  s5 = ~r4 & (~r5 & ~h3),
  t0 = \[4] ,
  t2 = ~z4 & (~y4 & ~y2),
  t3 = ~b0 | ~j0,
  t4 = ~e3 & ~s4,
  t5 = (~a4 & ~o4) | ~c0,
  u0 = \[5] ,
  u2 = (~f2 & ~m4) | ~d,
  u3 = ~e0,
  u4 = (~r3 & ~k0) | (~j0 & ~k0),
  u5 = ~h3 & ~r2,
  v0 = \[6] ,
  v2 = (~a & ~f2) | ((~a & ~z) | ((~z2 & ~f2) | (~z2 & ~z))),
  v3 = ~j,
  v4 = ~e & ~u4,
  v5 = (~h3 & ~g5) | (~y4 & ~g5),
  w0 = \[7] ,
  w2 = (~e5 & ~s5) | (~n0 & ~s5),
  w3 = ~k0 | (~b0 | ~e),
  w4 = ~k,
  w5 = ~a0 | ~i0,
  x0 = \[8] ,
  x2 = ~f5 | (~b0 | ~l),
  x3 = ~r3 | (~e | (~b0 | ~j0)),
  x4 = ~e & ~w4,
  y0 = \[9] ,
  y2 = ~o0,
  y3 = (~g0 & ~e0) | ~e,
  y4 = ~i,
  z0 = \[10] ,
  z2 = ~z,
  z3 = ~y3 | (~x3 | ~w3),
  z4 = ~d0,
  \[10]  = ~k5 | (~j5 | ~i5),
  \[11]  = (~h2 & ~g2) | (~n0 & ~g2),
  \[12]  = (~n0 & ~u5) | (~t4 & ~u5),
  \[13]  = ~w2,
  \[14]  = ~\[13] ;
endmodule

