module alu_2048(
  input wire a0, input wire b0,
  input wire a1, input wire b1,
  input wire a2, input wire b2,
  input wire a3, input wire b3,
  input wire a4, input wire b4,
  input wire a5, input wire b5,
  input wire a6, input wire b6,
  input wire a7, input wire b7,
  input wire a8, input wire b8,
  input wire a9, input wire b9,
  input wire a10, input wire b10,
  input wire a11, input wire b11,
  input wire a12, input wire b12,
  input wire a13, input wire b13,
  input wire a14, input wire b14,
  input wire a15, input wire b15,
  input wire a16, input wire b16,
  input wire a17, input wire b17,
  input wire a18, input wire b18,
  input wire a19, input wire b19,
  input wire a20, input wire b20,
  input wire a21, input wire b21,
  input wire a22, input wire b22,
  input wire a23, input wire b23,
  input wire a24, input wire b24,
  input wire a25, input wire b25,
  input wire a26, input wire b26,
  input wire a27, input wire b27,
  input wire a28, input wire b28,
  input wire a29, input wire b29,
  input wire a30, input wire b30,
  input wire a31, input wire b31,
  input wire a32, input wire b32,
  input wire a33, input wire b33,
  input wire a34, input wire b34,
  input wire a35, input wire b35,
  input wire a36, input wire b36,
  input wire a37, input wire b37,
  input wire a38, input wire b38,
  input wire a39, input wire b39,
  input wire a40, input wire b40,
  input wire a41, input wire b41,
  input wire a42, input wire b42,
  input wire a43, input wire b43,
  input wire a44, input wire b44,
  input wire a45, input wire b45,
  input wire a46, input wire b46,
  input wire a47, input wire b47,
  input wire a48, input wire b48,
  input wire a49, input wire b49,
  input wire a50, input wire b50,
  input wire a51, input wire b51,
  input wire a52, input wire b52,
  input wire a53, input wire b53,
  input wire a54, input wire b54,
  input wire a55, input wire b55,
  input wire a56, input wire b56,
  input wire a57, input wire b57,
  input wire a58, input wire b58,
  input wire a59, input wire b59,
  input wire a60, input wire b60,
  input wire a61, input wire b61,
  input wire a62, input wire b62,
  input wire a63, input wire b63,
  input wire a64, input wire b64,
  input wire a65, input wire b65,
  input wire a66, input wire b66,
  input wire a67, input wire b67,
  input wire a68, input wire b68,
  input wire a69, input wire b69,
  input wire a70, input wire b70,
  input wire a71, input wire b71,
  input wire a72, input wire b72,
  input wire a73, input wire b73,
  input wire a74, input wire b74,
  input wire a75, input wire b75,
  input wire a76, input wire b76,
  input wire a77, input wire b77,
  input wire a78, input wire b78,
  input wire a79, input wire b79,
  input wire a80, input wire b80,
  input wire a81, input wire b81,
  input wire a82, input wire b82,
  input wire a83, input wire b83,
  input wire a84, input wire b84,
  input wire a85, input wire b85,
  input wire a86, input wire b86,
  input wire a87, input wire b87,
  input wire a88, input wire b88,
  input wire a89, input wire b89,
  input wire a90, input wire b90,
  input wire a91, input wire b91,
  input wire a92, input wire b92,
  input wire a93, input wire b93,
  input wire a94, input wire b94,
  input wire a95, input wire b95,
  input wire a96, input wire b96,
  input wire a97, input wire b97,
  input wire a98, input wire b98,
  input wire a99, input wire b99,
  input wire a100, input wire b100,
  input wire a101, input wire b101,
  input wire a102, input wire b102,
  input wire a103, input wire b103,
  input wire a104, input wire b104,
  input wire a105, input wire b105,
  input wire a106, input wire b106,
  input wire a107, input wire b107,
  input wire a108, input wire b108,
  input wire a109, input wire b109,
  input wire a110, input wire b110,
  input wire a111, input wire b111,
  input wire a112, input wire b112,
  input wire a113, input wire b113,
  input wire a114, input wire b114,
  input wire a115, input wire b115,
  input wire a116, input wire b116,
  input wire a117, input wire b117,
  input wire a118, input wire b118,
  input wire a119, input wire b119,
  input wire a120, input wire b120,
  input wire a121, input wire b121,
  input wire a122, input wire b122,
  input wire a123, input wire b123,
  input wire a124, input wire b124,
  input wire a125, input wire b125,
  input wire a126, input wire b126,
  input wire a127, input wire b127,
  input wire a128, input wire b128,
  input wire a129, input wire b129,
  input wire a130, input wire b130,
  input wire a131, input wire b131,
  input wire a132, input wire b132,
  input wire a133, input wire b133,
  input wire a134, input wire b134,
  input wire a135, input wire b135,
  input wire a136, input wire b136,
  input wire a137, input wire b137,
  input wire a138, input wire b138,
  input wire a139, input wire b139,
  input wire a140, input wire b140,
  input wire a141, input wire b141,
  input wire a142, input wire b142,
  input wire a143, input wire b143,
  input wire a144, input wire b144,
  input wire a145, input wire b145,
  input wire a146, input wire b146,
  input wire a147, input wire b147,
  input wire a148, input wire b148,
  input wire a149, input wire b149,
  input wire a150, input wire b150,
  input wire a151, input wire b151,
  input wire a152, input wire b152,
  input wire a153, input wire b153,
  input wire a154, input wire b154,
  input wire a155, input wire b155,
  input wire a156, input wire b156,
  input wire a157, input wire b157,
  input wire a158, input wire b158,
  input wire a159, input wire b159,
  input wire a160, input wire b160,
  input wire a161, input wire b161,
  input wire a162, input wire b162,
  input wire a163, input wire b163,
  input wire a164, input wire b164,
  input wire a165, input wire b165,
  input wire a166, input wire b166,
  input wire a167, input wire b167,
  input wire a168, input wire b168,
  input wire a169, input wire b169,
  input wire a170, input wire b170,
  input wire a171, input wire b171,
  input wire a172, input wire b172,
  input wire a173, input wire b173,
  input wire a174, input wire b174,
  input wire a175, input wire b175,
  input wire a176, input wire b176,
  input wire a177, input wire b177,
  input wire a178, input wire b178,
  input wire a179, input wire b179,
  input wire a180, input wire b180,
  input wire a181, input wire b181,
  input wire a182, input wire b182,
  input wire a183, input wire b183,
  input wire a184, input wire b184,
  input wire a185, input wire b185,
  input wire a186, input wire b186,
  input wire a187, input wire b187,
  input wire a188, input wire b188,
  input wire a189, input wire b189,
  input wire a190, input wire b190,
  input wire a191, input wire b191,
  input wire a192, input wire b192,
  input wire a193, input wire b193,
  input wire a194, input wire b194,
  input wire a195, input wire b195,
  input wire a196, input wire b196,
  input wire a197, input wire b197,
  input wire a198, input wire b198,
  input wire a199, input wire b199,
  input wire a200, input wire b200,
  input wire a201, input wire b201,
  input wire a202, input wire b202,
  input wire a203, input wire b203,
  input wire a204, input wire b204,
  input wire a205, input wire b205,
  input wire a206, input wire b206,
  input wire a207, input wire b207,
  input wire a208, input wire b208,
  input wire a209, input wire b209,
  input wire a210, input wire b210,
  input wire a211, input wire b211,
  input wire a212, input wire b212,
  input wire a213, input wire b213,
  input wire a214, input wire b214,
  input wire a215, input wire b215,
  input wire a216, input wire b216,
  input wire a217, input wire b217,
  input wire a218, input wire b218,
  input wire a219, input wire b219,
  input wire a220, input wire b220,
  input wire a221, input wire b221,
  input wire a222, input wire b222,
  input wire a223, input wire b223,
  input wire a224, input wire b224,
  input wire a225, input wire b225,
  input wire a226, input wire b226,
  input wire a227, input wire b227,
  input wire a228, input wire b228,
  input wire a229, input wire b229,
  input wire a230, input wire b230,
  input wire a231, input wire b231,
  input wire a232, input wire b232,
  input wire a233, input wire b233,
  input wire a234, input wire b234,
  input wire a235, input wire b235,
  input wire a236, input wire b236,
  input wire a237, input wire b237,
  input wire a238, input wire b238,
  input wire a239, input wire b239,
  input wire a240, input wire b240,
  input wire a241, input wire b241,
  input wire a242, input wire b242,
  input wire a243, input wire b243,
  input wire a244, input wire b244,
  input wire a245, input wire b245,
  input wire a246, input wire b246,
  input wire a247, input wire b247,
  input wire a248, input wire b248,
  input wire a249, input wire b249,
  input wire a250, input wire b250,
  input wire a251, input wire b251,
  input wire a252, input wire b252,
  input wire a253, input wire b253,
  input wire a254, input wire b254,
  input wire a255, input wire b255,
  input wire a256, input wire b256,
  input wire a257, input wire b257,
  input wire a258, input wire b258,
  input wire a259, input wire b259,
  input wire a260, input wire b260,
  input wire a261, input wire b261,
  input wire a262, input wire b262,
  input wire a263, input wire b263,
  input wire a264, input wire b264,
  input wire a265, input wire b265,
  input wire a266, input wire b266,
  input wire a267, input wire b267,
  input wire a268, input wire b268,
  input wire a269, input wire b269,
  input wire a270, input wire b270,
  input wire a271, input wire b271,
  input wire a272, input wire b272,
  input wire a273, input wire b273,
  input wire a274, input wire b274,
  input wire a275, input wire b275,
  input wire a276, input wire b276,
  input wire a277, input wire b277,
  input wire a278, input wire b278,
  input wire a279, input wire b279,
  input wire a280, input wire b280,
  input wire a281, input wire b281,
  input wire a282, input wire b282,
  input wire a283, input wire b283,
  input wire a284, input wire b284,
  input wire a285, input wire b285,
  input wire a286, input wire b286,
  input wire a287, input wire b287,
  input wire a288, input wire b288,
  input wire a289, input wire b289,
  input wire a290, input wire b290,
  input wire a291, input wire b291,
  input wire a292, input wire b292,
  input wire a293, input wire b293,
  input wire a294, input wire b294,
  input wire a295, input wire b295,
  input wire a296, input wire b296,
  input wire a297, input wire b297,
  input wire a298, input wire b298,
  input wire a299, input wire b299,
  input wire a300, input wire b300,
  input wire a301, input wire b301,
  input wire a302, input wire b302,
  input wire a303, input wire b303,
  input wire a304, input wire b304,
  input wire a305, input wire b305,
  input wire a306, input wire b306,
  input wire a307, input wire b307,
  input wire a308, input wire b308,
  input wire a309, input wire b309,
  input wire a310, input wire b310,
  input wire a311, input wire b311,
  input wire a312, input wire b312,
  input wire a313, input wire b313,
  input wire a314, input wire b314,
  input wire a315, input wire b315,
  input wire a316, input wire b316,
  input wire a317, input wire b317,
  input wire a318, input wire b318,
  input wire a319, input wire b319,
  input wire a320, input wire b320,
  input wire a321, input wire b321,
  input wire a322, input wire b322,
  input wire a323, input wire b323,
  input wire a324, input wire b324,
  input wire a325, input wire b325,
  input wire a326, input wire b326,
  input wire a327, input wire b327,
  input wire a328, input wire b328,
  input wire a329, input wire b329,
  input wire a330, input wire b330,
  input wire a331, input wire b331,
  input wire a332, input wire b332,
  input wire a333, input wire b333,
  input wire a334, input wire b334,
  input wire a335, input wire b335,
  input wire a336, input wire b336,
  input wire a337, input wire b337,
  input wire a338, input wire b338,
  input wire a339, input wire b339,
  input wire a340, input wire b340,
  input wire a341, input wire b341,
  input wire a342, input wire b342,
  input wire a343, input wire b343,
  input wire a344, input wire b344,
  input wire a345, input wire b345,
  input wire a346, input wire b346,
  input wire a347, input wire b347,
  input wire a348, input wire b348,
  input wire a349, input wire b349,
  input wire a350, input wire b350,
  input wire a351, input wire b351,
  input wire a352, input wire b352,
  input wire a353, input wire b353,
  input wire a354, input wire b354,
  input wire a355, input wire b355,
  input wire a356, input wire b356,
  input wire a357, input wire b357,
  input wire a358, input wire b358,
  input wire a359, input wire b359,
  input wire a360, input wire b360,
  input wire a361, input wire b361,
  input wire a362, input wire b362,
  input wire a363, input wire b363,
  input wire a364, input wire b364,
  input wire a365, input wire b365,
  input wire a366, input wire b366,
  input wire a367, input wire b367,
  input wire a368, input wire b368,
  input wire a369, input wire b369,
  input wire a370, input wire b370,
  input wire a371, input wire b371,
  input wire a372, input wire b372,
  input wire a373, input wire b373,
  input wire a374, input wire b374,
  input wire a375, input wire b375,
  input wire a376, input wire b376,
  input wire a377, input wire b377,
  input wire a378, input wire b378,
  input wire a379, input wire b379,
  input wire a380, input wire b380,
  input wire a381, input wire b381,
  input wire a382, input wire b382,
  input wire a383, input wire b383,
  input wire a384, input wire b384,
  input wire a385, input wire b385,
  input wire a386, input wire b386,
  input wire a387, input wire b387,
  input wire a388, input wire b388,
  input wire a389, input wire b389,
  input wire a390, input wire b390,
  input wire a391, input wire b391,
  input wire a392, input wire b392,
  input wire a393, input wire b393,
  input wire a394, input wire b394,
  input wire a395, input wire b395,
  input wire a396, input wire b396,
  input wire a397, input wire b397,
  input wire a398, input wire b398,
  input wire a399, input wire b399,
  input wire a400, input wire b400,
  input wire a401, input wire b401,
  input wire a402, input wire b402,
  input wire a403, input wire b403,
  input wire a404, input wire b404,
  input wire a405, input wire b405,
  input wire a406, input wire b406,
  input wire a407, input wire b407,
  input wire a408, input wire b408,
  input wire a409, input wire b409,
  input wire a410, input wire b410,
  input wire a411, input wire b411,
  input wire a412, input wire b412,
  input wire a413, input wire b413,
  input wire a414, input wire b414,
  input wire a415, input wire b415,
  input wire a416, input wire b416,
  input wire a417, input wire b417,
  input wire a418, input wire b418,
  input wire a419, input wire b419,
  input wire a420, input wire b420,
  input wire a421, input wire b421,
  input wire a422, input wire b422,
  input wire a423, input wire b423,
  input wire a424, input wire b424,
  input wire a425, input wire b425,
  input wire a426, input wire b426,
  input wire a427, input wire b427,
  input wire a428, input wire b428,
  input wire a429, input wire b429,
  input wire a430, input wire b430,
  input wire a431, input wire b431,
  input wire a432, input wire b432,
  input wire a433, input wire b433,
  input wire a434, input wire b434,
  input wire a435, input wire b435,
  input wire a436, input wire b436,
  input wire a437, input wire b437,
  input wire a438, input wire b438,
  input wire a439, input wire b439,
  input wire a440, input wire b440,
  input wire a441, input wire b441,
  input wire a442, input wire b442,
  input wire a443, input wire b443,
  input wire a444, input wire b444,
  input wire a445, input wire b445,
  input wire a446, input wire b446,
  input wire a447, input wire b447,
  input wire a448, input wire b448,
  input wire a449, input wire b449,
  input wire a450, input wire b450,
  input wire a451, input wire b451,
  input wire a452, input wire b452,
  input wire a453, input wire b453,
  input wire a454, input wire b454,
  input wire a455, input wire b455,
  input wire a456, input wire b456,
  input wire a457, input wire b457,
  input wire a458, input wire b458,
  input wire a459, input wire b459,
  input wire a460, input wire b460,
  input wire a461, input wire b461,
  input wire a462, input wire b462,
  input wire a463, input wire b463,
  input wire a464, input wire b464,
  input wire a465, input wire b465,
  input wire a466, input wire b466,
  input wire a467, input wire b467,
  input wire a468, input wire b468,
  input wire a469, input wire b469,
  input wire a470, input wire b470,
  input wire a471, input wire b471,
  input wire a472, input wire b472,
  input wire a473, input wire b473,
  input wire a474, input wire b474,
  input wire a475, input wire b475,
  input wire a476, input wire b476,
  input wire a477, input wire b477,
  input wire a478, input wire b478,
  input wire a479, input wire b479,
  input wire a480, input wire b480,
  input wire a481, input wire b481,
  input wire a482, input wire b482,
  input wire a483, input wire b483,
  input wire a484, input wire b484,
  input wire a485, input wire b485,
  input wire a486, input wire b486,
  input wire a487, input wire b487,
  input wire a488, input wire b488,
  input wire a489, input wire b489,
  input wire a490, input wire b490,
  input wire a491, input wire b491,
  input wire a492, input wire b492,
  input wire a493, input wire b493,
  input wire a494, input wire b494,
  input wire a495, input wire b495,
  input wire a496, input wire b496,
  input wire a497, input wire b497,
  input wire a498, input wire b498,
  input wire a499, input wire b499,
  input wire a500, input wire b500,
  input wire a501, input wire b501,
  input wire a502, input wire b502,
  input wire a503, input wire b503,
  input wire a504, input wire b504,
  input wire a505, input wire b505,
  input wire a506, input wire b506,
  input wire a507, input wire b507,
  input wire a508, input wire b508,
  input wire a509, input wire b509,
  input wire a510, input wire b510,
  input wire a511, input wire b511,
  input wire a512, input wire b512,
  input wire a513, input wire b513,
  input wire a514, input wire b514,
  input wire a515, input wire b515,
  input wire a516, input wire b516,
  input wire a517, input wire b517,
  input wire a518, input wire b518,
  input wire a519, input wire b519,
  input wire a520, input wire b520,
  input wire a521, input wire b521,
  input wire a522, input wire b522,
  input wire a523, input wire b523,
  input wire a524, input wire b524,
  input wire a525, input wire b525,
  input wire a526, input wire b526,
  input wire a527, input wire b527,
  input wire a528, input wire b528,
  input wire a529, input wire b529,
  input wire a530, input wire b530,
  input wire a531, input wire b531,
  input wire a532, input wire b532,
  input wire a533, input wire b533,
  input wire a534, input wire b534,
  input wire a535, input wire b535,
  input wire a536, input wire b536,
  input wire a537, input wire b537,
  input wire a538, input wire b538,
  input wire a539, input wire b539,
  input wire a540, input wire b540,
  input wire a541, input wire b541,
  input wire a542, input wire b542,
  input wire a543, input wire b543,
  input wire a544, input wire b544,
  input wire a545, input wire b545,
  input wire a546, input wire b546,
  input wire a547, input wire b547,
  input wire a548, input wire b548,
  input wire a549, input wire b549,
  input wire a550, input wire b550,
  input wire a551, input wire b551,
  input wire a552, input wire b552,
  input wire a553, input wire b553,
  input wire a554, input wire b554,
  input wire a555, input wire b555,
  input wire a556, input wire b556,
  input wire a557, input wire b557,
  input wire a558, input wire b558,
  input wire a559, input wire b559,
  input wire a560, input wire b560,
  input wire a561, input wire b561,
  input wire a562, input wire b562,
  input wire a563, input wire b563,
  input wire a564, input wire b564,
  input wire a565, input wire b565,
  input wire a566, input wire b566,
  input wire a567, input wire b567,
  input wire a568, input wire b568,
  input wire a569, input wire b569,
  input wire a570, input wire b570,
  input wire a571, input wire b571,
  input wire a572, input wire b572,
  input wire a573, input wire b573,
  input wire a574, input wire b574,
  input wire a575, input wire b575,
  input wire a576, input wire b576,
  input wire a577, input wire b577,
  input wire a578, input wire b578,
  input wire a579, input wire b579,
  input wire a580, input wire b580,
  input wire a581, input wire b581,
  input wire a582, input wire b582,
  input wire a583, input wire b583,
  input wire a584, input wire b584,
  input wire a585, input wire b585,
  input wire a586, input wire b586,
  input wire a587, input wire b587,
  input wire a588, input wire b588,
  input wire a589, input wire b589,
  input wire a590, input wire b590,
  input wire a591, input wire b591,
  input wire a592, input wire b592,
  input wire a593, input wire b593,
  input wire a594, input wire b594,
  input wire a595, input wire b595,
  input wire a596, input wire b596,
  input wire a597, input wire b597,
  input wire a598, input wire b598,
  input wire a599, input wire b599,
  input wire a600, input wire b600,
  input wire a601, input wire b601,
  input wire a602, input wire b602,
  input wire a603, input wire b603,
  input wire a604, input wire b604,
  input wire a605, input wire b605,
  input wire a606, input wire b606,
  input wire a607, input wire b607,
  input wire a608, input wire b608,
  input wire a609, input wire b609,
  input wire a610, input wire b610,
  input wire a611, input wire b611,
  input wire a612, input wire b612,
  input wire a613, input wire b613,
  input wire a614, input wire b614,
  input wire a615, input wire b615,
  input wire a616, input wire b616,
  input wire a617, input wire b617,
  input wire a618, input wire b618,
  input wire a619, input wire b619,
  input wire a620, input wire b620,
  input wire a621, input wire b621,
  input wire a622, input wire b622,
  input wire a623, input wire b623,
  input wire a624, input wire b624,
  input wire a625, input wire b625,
  input wire a626, input wire b626,
  input wire a627, input wire b627,
  input wire a628, input wire b628,
  input wire a629, input wire b629,
  input wire a630, input wire b630,
  input wire a631, input wire b631,
  input wire a632, input wire b632,
  input wire a633, input wire b633,
  input wire a634, input wire b634,
  input wire a635, input wire b635,
  input wire a636, input wire b636,
  input wire a637, input wire b637,
  input wire a638, input wire b638,
  input wire a639, input wire b639,
  input wire a640, input wire b640,
  input wire a641, input wire b641,
  input wire a642, input wire b642,
  input wire a643, input wire b643,
  input wire a644, input wire b644,
  input wire a645, input wire b645,
  input wire a646, input wire b646,
  input wire a647, input wire b647,
  input wire a648, input wire b648,
  input wire a649, input wire b649,
  input wire a650, input wire b650,
  input wire a651, input wire b651,
  input wire a652, input wire b652,
  input wire a653, input wire b653,
  input wire a654, input wire b654,
  input wire a655, input wire b655,
  input wire a656, input wire b656,
  input wire a657, input wire b657,
  input wire a658, input wire b658,
  input wire a659, input wire b659,
  input wire a660, input wire b660,
  input wire a661, input wire b661,
  input wire a662, input wire b662,
  input wire a663, input wire b663,
  input wire a664, input wire b664,
  input wire a665, input wire b665,
  input wire a666, input wire b666,
  input wire a667, input wire b667,
  input wire a668, input wire b668,
  input wire a669, input wire b669,
  input wire a670, input wire b670,
  input wire a671, input wire b671,
  input wire a672, input wire b672,
  input wire a673, input wire b673,
  input wire a674, input wire b674,
  input wire a675, input wire b675,
  input wire a676, input wire b676,
  input wire a677, input wire b677,
  input wire a678, input wire b678,
  input wire a679, input wire b679,
  input wire a680, input wire b680,
  input wire a681, input wire b681,
  input wire a682, input wire b682,
  input wire a683, input wire b683,
  input wire a684, input wire b684,
  input wire a685, input wire b685,
  input wire a686, input wire b686,
  input wire a687, input wire b687,
  input wire a688, input wire b688,
  input wire a689, input wire b689,
  input wire a690, input wire b690,
  input wire a691, input wire b691,
  input wire a692, input wire b692,
  input wire a693, input wire b693,
  input wire a694, input wire b694,
  input wire a695, input wire b695,
  input wire a696, input wire b696,
  input wire a697, input wire b697,
  input wire a698, input wire b698,
  input wire a699, input wire b699,
  input wire a700, input wire b700,
  input wire a701, input wire b701,
  input wire a702, input wire b702,
  input wire a703, input wire b703,
  input wire a704, input wire b704,
  input wire a705, input wire b705,
  input wire a706, input wire b706,
  input wire a707, input wire b707,
  input wire a708, input wire b708,
  input wire a709, input wire b709,
  input wire a710, input wire b710,
  input wire a711, input wire b711,
  input wire a712, input wire b712,
  input wire a713, input wire b713,
  input wire a714, input wire b714,
  input wire a715, input wire b715,
  input wire a716, input wire b716,
  input wire a717, input wire b717,
  input wire a718, input wire b718,
  input wire a719, input wire b719,
  input wire a720, input wire b720,
  input wire a721, input wire b721,
  input wire a722, input wire b722,
  input wire a723, input wire b723,
  input wire a724, input wire b724,
  input wire a725, input wire b725,
  input wire a726, input wire b726,
  input wire a727, input wire b727,
  input wire a728, input wire b728,
  input wire a729, input wire b729,
  input wire a730, input wire b730,
  input wire a731, input wire b731,
  input wire a732, input wire b732,
  input wire a733, input wire b733,
  input wire a734, input wire b734,
  input wire a735, input wire b735,
  input wire a736, input wire b736,
  input wire a737, input wire b737,
  input wire a738, input wire b738,
  input wire a739, input wire b739,
  input wire a740, input wire b740,
  input wire a741, input wire b741,
  input wire a742, input wire b742,
  input wire a743, input wire b743,
  input wire a744, input wire b744,
  input wire a745, input wire b745,
  input wire a746, input wire b746,
  input wire a747, input wire b747,
  input wire a748, input wire b748,
  input wire a749, input wire b749,
  input wire a750, input wire b750,
  input wire a751, input wire b751,
  input wire a752, input wire b752,
  input wire a753, input wire b753,
  input wire a754, input wire b754,
  input wire a755, input wire b755,
  input wire a756, input wire b756,
  input wire a757, input wire b757,
  input wire a758, input wire b758,
  input wire a759, input wire b759,
  input wire a760, input wire b760,
  input wire a761, input wire b761,
  input wire a762, input wire b762,
  input wire a763, input wire b763,
  input wire a764, input wire b764,
  input wire a765, input wire b765,
  input wire a766, input wire b766,
  input wire a767, input wire b767,
  input wire a768, input wire b768,
  input wire a769, input wire b769,
  input wire a770, input wire b770,
  input wire a771, input wire b771,
  input wire a772, input wire b772,
  input wire a773, input wire b773,
  input wire a774, input wire b774,
  input wire a775, input wire b775,
  input wire a776, input wire b776,
  input wire a777, input wire b777,
  input wire a778, input wire b778,
  input wire a779, input wire b779,
  input wire a780, input wire b780,
  input wire a781, input wire b781,
  input wire a782, input wire b782,
  input wire a783, input wire b783,
  input wire a784, input wire b784,
  input wire a785, input wire b785,
  input wire a786, input wire b786,
  input wire a787, input wire b787,
  input wire a788, input wire b788,
  input wire a789, input wire b789,
  input wire a790, input wire b790,
  input wire a791, input wire b791,
  input wire a792, input wire b792,
  input wire a793, input wire b793,
  input wire a794, input wire b794,
  input wire a795, input wire b795,
  input wire a796, input wire b796,
  input wire a797, input wire b797,
  input wire a798, input wire b798,
  input wire a799, input wire b799,
  input wire a800, input wire b800,
  input wire a801, input wire b801,
  input wire a802, input wire b802,
  input wire a803, input wire b803,
  input wire a804, input wire b804,
  input wire a805, input wire b805,
  input wire a806, input wire b806,
  input wire a807, input wire b807,
  input wire a808, input wire b808,
  input wire a809, input wire b809,
  input wire a810, input wire b810,
  input wire a811, input wire b811,
  input wire a812, input wire b812,
  input wire a813, input wire b813,
  input wire a814, input wire b814,
  input wire a815, input wire b815,
  input wire a816, input wire b816,
  input wire a817, input wire b817,
  input wire a818, input wire b818,
  input wire a819, input wire b819,
  input wire a820, input wire b820,
  input wire a821, input wire b821,
  input wire a822, input wire b822,
  input wire a823, input wire b823,
  input wire a824, input wire b824,
  input wire a825, input wire b825,
  input wire a826, input wire b826,
  input wire a827, input wire b827,
  input wire a828, input wire b828,
  input wire a829, input wire b829,
  input wire a830, input wire b830,
  input wire a831, input wire b831,
  input wire a832, input wire b832,
  input wire a833, input wire b833,
  input wire a834, input wire b834,
  input wire a835, input wire b835,
  input wire a836, input wire b836,
  input wire a837, input wire b837,
  input wire a838, input wire b838,
  input wire a839, input wire b839,
  input wire a840, input wire b840,
  input wire a841, input wire b841,
  input wire a842, input wire b842,
  input wire a843, input wire b843,
  input wire a844, input wire b844,
  input wire a845, input wire b845,
  input wire a846, input wire b846,
  input wire a847, input wire b847,
  input wire a848, input wire b848,
  input wire a849, input wire b849,
  input wire a850, input wire b850,
  input wire a851, input wire b851,
  input wire a852, input wire b852,
  input wire a853, input wire b853,
  input wire a854, input wire b854,
  input wire a855, input wire b855,
  input wire a856, input wire b856,
  input wire a857, input wire b857,
  input wire a858, input wire b858,
  input wire a859, input wire b859,
  input wire a860, input wire b860,
  input wire a861, input wire b861,
  input wire a862, input wire b862,
  input wire a863, input wire b863,
  input wire a864, input wire b864,
  input wire a865, input wire b865,
  input wire a866, input wire b866,
  input wire a867, input wire b867,
  input wire a868, input wire b868,
  input wire a869, input wire b869,
  input wire a870, input wire b870,
  input wire a871, input wire b871,
  input wire a872, input wire b872,
  input wire a873, input wire b873,
  input wire a874, input wire b874,
  input wire a875, input wire b875,
  input wire a876, input wire b876,
  input wire a877, input wire b877,
  input wire a878, input wire b878,
  input wire a879, input wire b879,
  input wire a880, input wire b880,
  input wire a881, input wire b881,
  input wire a882, input wire b882,
  input wire a883, input wire b883,
  input wire a884, input wire b884,
  input wire a885, input wire b885,
  input wire a886, input wire b886,
  input wire a887, input wire b887,
  input wire a888, input wire b888,
  input wire a889, input wire b889,
  input wire a890, input wire b890,
  input wire a891, input wire b891,
  input wire a892, input wire b892,
  input wire a893, input wire b893,
  input wire a894, input wire b894,
  input wire a895, input wire b895,
  input wire a896, input wire b896,
  input wire a897, input wire b897,
  input wire a898, input wire b898,
  input wire a899, input wire b899,
  input wire a900, input wire b900,
  input wire a901, input wire b901,
  input wire a902, input wire b902,
  input wire a903, input wire b903,
  input wire a904, input wire b904,
  input wire a905, input wire b905,
  input wire a906, input wire b906,
  input wire a907, input wire b907,
  input wire a908, input wire b908,
  input wire a909, input wire b909,
  input wire a910, input wire b910,
  input wire a911, input wire b911,
  input wire a912, input wire b912,
  input wire a913, input wire b913,
  input wire a914, input wire b914,
  input wire a915, input wire b915,
  input wire a916, input wire b916,
  input wire a917, input wire b917,
  input wire a918, input wire b918,
  input wire a919, input wire b919,
  input wire a920, input wire b920,
  input wire a921, input wire b921,
  input wire a922, input wire b922,
  input wire a923, input wire b923,
  input wire a924, input wire b924,
  input wire a925, input wire b925,
  input wire a926, input wire b926,
  input wire a927, input wire b927,
  input wire a928, input wire b928,
  input wire a929, input wire b929,
  input wire a930, input wire b930,
  input wire a931, input wire b931,
  input wire a932, input wire b932,
  input wire a933, input wire b933,
  input wire a934, input wire b934,
  input wire a935, input wire b935,
  input wire a936, input wire b936,
  input wire a937, input wire b937,
  input wire a938, input wire b938,
  input wire a939, input wire b939,
  input wire a940, input wire b940,
  input wire a941, input wire b941,
  input wire a942, input wire b942,
  input wire a943, input wire b943,
  input wire a944, input wire b944,
  input wire a945, input wire b945,
  input wire a946, input wire b946,
  input wire a947, input wire b947,
  input wire a948, input wire b948,
  input wire a949, input wire b949,
  input wire a950, input wire b950,
  input wire a951, input wire b951,
  input wire a952, input wire b952,
  input wire a953, input wire b953,
  input wire a954, input wire b954,
  input wire a955, input wire b955,
  input wire a956, input wire b956,
  input wire a957, input wire b957,
  input wire a958, input wire b958,
  input wire a959, input wire b959,
  input wire a960, input wire b960,
  input wire a961, input wire b961,
  input wire a962, input wire b962,
  input wire a963, input wire b963,
  input wire a964, input wire b964,
  input wire a965, input wire b965,
  input wire a966, input wire b966,
  input wire a967, input wire b967,
  input wire a968, input wire b968,
  input wire a969, input wire b969,
  input wire a970, input wire b970,
  input wire a971, input wire b971,
  input wire a972, input wire b972,
  input wire a973, input wire b973,
  input wire a974, input wire b974,
  input wire a975, input wire b975,
  input wire a976, input wire b976,
  input wire a977, input wire b977,
  input wire a978, input wire b978,
  input wire a979, input wire b979,
  input wire a980, input wire b980,
  input wire a981, input wire b981,
  input wire a982, input wire b982,
  input wire a983, input wire b983,
  input wire a984, input wire b984,
  input wire a985, input wire b985,
  input wire a986, input wire b986,
  input wire a987, input wire b987,
  input wire a988, input wire b988,
  input wire a989, input wire b989,
  input wire a990, input wire b990,
  input wire a991, input wire b991,
  input wire a992, input wire b992,
  input wire a993, input wire b993,
  input wire a994, input wire b994,
  input wire a995, input wire b995,
  input wire a996, input wire b996,
  input wire a997, input wire b997,
  input wire a998, input wire b998,
  input wire a999, input wire b999,
  input wire a1000, input wire b1000,
  input wire a1001, input wire b1001,
  input wire a1002, input wire b1002,
  input wire a1003, input wire b1003,
  input wire a1004, input wire b1004,
  input wire a1005, input wire b1005,
  input wire a1006, input wire b1006,
  input wire a1007, input wire b1007,
  input wire a1008, input wire b1008,
  input wire a1009, input wire b1009,
  input wire a1010, input wire b1010,
  input wire a1011, input wire b1011,
  input wire a1012, input wire b1012,
  input wire a1013, input wire b1013,
  input wire a1014, input wire b1014,
  input wire a1015, input wire b1015,
  input wire a1016, input wire b1016,
  input wire a1017, input wire b1017,
  input wire a1018, input wire b1018,
  input wire a1019, input wire b1019,
  input wire a1020, input wire b1020,
  input wire a1021, input wire b1021,
  input wire a1022, input wire b1022,
  input wire a1023, input wire b1023,
  input wire a1024, input wire b1024,
  input wire a1025, input wire b1025,
  input wire a1026, input wire b1026,
  input wire a1027, input wire b1027,
  input wire a1028, input wire b1028,
  input wire a1029, input wire b1029,
  input wire a1030, input wire b1030,
  input wire a1031, input wire b1031,
  input wire a1032, input wire b1032,
  input wire a1033, input wire b1033,
  input wire a1034, input wire b1034,
  input wire a1035, input wire b1035,
  input wire a1036, input wire b1036,
  input wire a1037, input wire b1037,
  input wire a1038, input wire b1038,
  input wire a1039, input wire b1039,
  input wire a1040, input wire b1040,
  input wire a1041, input wire b1041,
  input wire a1042, input wire b1042,
  input wire a1043, input wire b1043,
  input wire a1044, input wire b1044,
  input wire a1045, input wire b1045,
  input wire a1046, input wire b1046,
  input wire a1047, input wire b1047,
  input wire a1048, input wire b1048,
  input wire a1049, input wire b1049,
  input wire a1050, input wire b1050,
  input wire a1051, input wire b1051,
  input wire a1052, input wire b1052,
  input wire a1053, input wire b1053,
  input wire a1054, input wire b1054,
  input wire a1055, input wire b1055,
  input wire a1056, input wire b1056,
  input wire a1057, input wire b1057,
  input wire a1058, input wire b1058,
  input wire a1059, input wire b1059,
  input wire a1060, input wire b1060,
  input wire a1061, input wire b1061,
  input wire a1062, input wire b1062,
  input wire a1063, input wire b1063,
  input wire a1064, input wire b1064,
  input wire a1065, input wire b1065,
  input wire a1066, input wire b1066,
  input wire a1067, input wire b1067,
  input wire a1068, input wire b1068,
  input wire a1069, input wire b1069,
  input wire a1070, input wire b1070,
  input wire a1071, input wire b1071,
  input wire a1072, input wire b1072,
  input wire a1073, input wire b1073,
  input wire a1074, input wire b1074,
  input wire a1075, input wire b1075,
  input wire a1076, input wire b1076,
  input wire a1077, input wire b1077,
  input wire a1078, input wire b1078,
  input wire a1079, input wire b1079,
  input wire a1080, input wire b1080,
  input wire a1081, input wire b1081,
  input wire a1082, input wire b1082,
  input wire a1083, input wire b1083,
  input wire a1084, input wire b1084,
  input wire a1085, input wire b1085,
  input wire a1086, input wire b1086,
  input wire a1087, input wire b1087,
  input wire a1088, input wire b1088,
  input wire a1089, input wire b1089,
  input wire a1090, input wire b1090,
  input wire a1091, input wire b1091,
  input wire a1092, input wire b1092,
  input wire a1093, input wire b1093,
  input wire a1094, input wire b1094,
  input wire a1095, input wire b1095,
  input wire a1096, input wire b1096,
  input wire a1097, input wire b1097,
  input wire a1098, input wire b1098,
  input wire a1099, input wire b1099,
  input wire a1100, input wire b1100,
  input wire a1101, input wire b1101,
  input wire a1102, input wire b1102,
  input wire a1103, input wire b1103,
  input wire a1104, input wire b1104,
  input wire a1105, input wire b1105,
  input wire a1106, input wire b1106,
  input wire a1107, input wire b1107,
  input wire a1108, input wire b1108,
  input wire a1109, input wire b1109,
  input wire a1110, input wire b1110,
  input wire a1111, input wire b1111,
  input wire a1112, input wire b1112,
  input wire a1113, input wire b1113,
  input wire a1114, input wire b1114,
  input wire a1115, input wire b1115,
  input wire a1116, input wire b1116,
  input wire a1117, input wire b1117,
  input wire a1118, input wire b1118,
  input wire a1119, input wire b1119,
  input wire a1120, input wire b1120,
  input wire a1121, input wire b1121,
  input wire a1122, input wire b1122,
  input wire a1123, input wire b1123,
  input wire a1124, input wire b1124,
  input wire a1125, input wire b1125,
  input wire a1126, input wire b1126,
  input wire a1127, input wire b1127,
  input wire a1128, input wire b1128,
  input wire a1129, input wire b1129,
  input wire a1130, input wire b1130,
  input wire a1131, input wire b1131,
  input wire a1132, input wire b1132,
  input wire a1133, input wire b1133,
  input wire a1134, input wire b1134,
  input wire a1135, input wire b1135,
  input wire a1136, input wire b1136,
  input wire a1137, input wire b1137,
  input wire a1138, input wire b1138,
  input wire a1139, input wire b1139,
  input wire a1140, input wire b1140,
  input wire a1141, input wire b1141,
  input wire a1142, input wire b1142,
  input wire a1143, input wire b1143,
  input wire a1144, input wire b1144,
  input wire a1145, input wire b1145,
  input wire a1146, input wire b1146,
  input wire a1147, input wire b1147,
  input wire a1148, input wire b1148,
  input wire a1149, input wire b1149,
  input wire a1150, input wire b1150,
  input wire a1151, input wire b1151,
  input wire a1152, input wire b1152,
  input wire a1153, input wire b1153,
  input wire a1154, input wire b1154,
  input wire a1155, input wire b1155,
  input wire a1156, input wire b1156,
  input wire a1157, input wire b1157,
  input wire a1158, input wire b1158,
  input wire a1159, input wire b1159,
  input wire a1160, input wire b1160,
  input wire a1161, input wire b1161,
  input wire a1162, input wire b1162,
  input wire a1163, input wire b1163,
  input wire a1164, input wire b1164,
  input wire a1165, input wire b1165,
  input wire a1166, input wire b1166,
  input wire a1167, input wire b1167,
  input wire a1168, input wire b1168,
  input wire a1169, input wire b1169,
  input wire a1170, input wire b1170,
  input wire a1171, input wire b1171,
  input wire a1172, input wire b1172,
  input wire a1173, input wire b1173,
  input wire a1174, input wire b1174,
  input wire a1175, input wire b1175,
  input wire a1176, input wire b1176,
  input wire a1177, input wire b1177,
  input wire a1178, input wire b1178,
  input wire a1179, input wire b1179,
  input wire a1180, input wire b1180,
  input wire a1181, input wire b1181,
  input wire a1182, input wire b1182,
  input wire a1183, input wire b1183,
  input wire a1184, input wire b1184,
  input wire a1185, input wire b1185,
  input wire a1186, input wire b1186,
  input wire a1187, input wire b1187,
  input wire a1188, input wire b1188,
  input wire a1189, input wire b1189,
  input wire a1190, input wire b1190,
  input wire a1191, input wire b1191,
  input wire a1192, input wire b1192,
  input wire a1193, input wire b1193,
  input wire a1194, input wire b1194,
  input wire a1195, input wire b1195,
  input wire a1196, input wire b1196,
  input wire a1197, input wire b1197,
  input wire a1198, input wire b1198,
  input wire a1199, input wire b1199,
  input wire a1200, input wire b1200,
  input wire a1201, input wire b1201,
  input wire a1202, input wire b1202,
  input wire a1203, input wire b1203,
  input wire a1204, input wire b1204,
  input wire a1205, input wire b1205,
  input wire a1206, input wire b1206,
  input wire a1207, input wire b1207,
  input wire a1208, input wire b1208,
  input wire a1209, input wire b1209,
  input wire a1210, input wire b1210,
  input wire a1211, input wire b1211,
  input wire a1212, input wire b1212,
  input wire a1213, input wire b1213,
  input wire a1214, input wire b1214,
  input wire a1215, input wire b1215,
  input wire a1216, input wire b1216,
  input wire a1217, input wire b1217,
  input wire a1218, input wire b1218,
  input wire a1219, input wire b1219,
  input wire a1220, input wire b1220,
  input wire a1221, input wire b1221,
  input wire a1222, input wire b1222,
  input wire a1223, input wire b1223,
  input wire a1224, input wire b1224,
  input wire a1225, input wire b1225,
  input wire a1226, input wire b1226,
  input wire a1227, input wire b1227,
  input wire a1228, input wire b1228,
  input wire a1229, input wire b1229,
  input wire a1230, input wire b1230,
  input wire a1231, input wire b1231,
  input wire a1232, input wire b1232,
  input wire a1233, input wire b1233,
  input wire a1234, input wire b1234,
  input wire a1235, input wire b1235,
  input wire a1236, input wire b1236,
  input wire a1237, input wire b1237,
  input wire a1238, input wire b1238,
  input wire a1239, input wire b1239,
  input wire a1240, input wire b1240,
  input wire a1241, input wire b1241,
  input wire a1242, input wire b1242,
  input wire a1243, input wire b1243,
  input wire a1244, input wire b1244,
  input wire a1245, input wire b1245,
  input wire a1246, input wire b1246,
  input wire a1247, input wire b1247,
  input wire a1248, input wire b1248,
  input wire a1249, input wire b1249,
  input wire a1250, input wire b1250,
  input wire a1251, input wire b1251,
  input wire a1252, input wire b1252,
  input wire a1253, input wire b1253,
  input wire a1254, input wire b1254,
  input wire a1255, input wire b1255,
  input wire a1256, input wire b1256,
  input wire a1257, input wire b1257,
  input wire a1258, input wire b1258,
  input wire a1259, input wire b1259,
  input wire a1260, input wire b1260,
  input wire a1261, input wire b1261,
  input wire a1262, input wire b1262,
  input wire a1263, input wire b1263,
  input wire a1264, input wire b1264,
  input wire a1265, input wire b1265,
  input wire a1266, input wire b1266,
  input wire a1267, input wire b1267,
  input wire a1268, input wire b1268,
  input wire a1269, input wire b1269,
  input wire a1270, input wire b1270,
  input wire a1271, input wire b1271,
  input wire a1272, input wire b1272,
  input wire a1273, input wire b1273,
  input wire a1274, input wire b1274,
  input wire a1275, input wire b1275,
  input wire a1276, input wire b1276,
  input wire a1277, input wire b1277,
  input wire a1278, input wire b1278,
  input wire a1279, input wire b1279,
  input wire a1280, input wire b1280,
  input wire a1281, input wire b1281,
  input wire a1282, input wire b1282,
  input wire a1283, input wire b1283,
  input wire a1284, input wire b1284,
  input wire a1285, input wire b1285,
  input wire a1286, input wire b1286,
  input wire a1287, input wire b1287,
  input wire a1288, input wire b1288,
  input wire a1289, input wire b1289,
  input wire a1290, input wire b1290,
  input wire a1291, input wire b1291,
  input wire a1292, input wire b1292,
  input wire a1293, input wire b1293,
  input wire a1294, input wire b1294,
  input wire a1295, input wire b1295,
  input wire a1296, input wire b1296,
  input wire a1297, input wire b1297,
  input wire a1298, input wire b1298,
  input wire a1299, input wire b1299,
  input wire a1300, input wire b1300,
  input wire a1301, input wire b1301,
  input wire a1302, input wire b1302,
  input wire a1303, input wire b1303,
  input wire a1304, input wire b1304,
  input wire a1305, input wire b1305,
  input wire a1306, input wire b1306,
  input wire a1307, input wire b1307,
  input wire a1308, input wire b1308,
  input wire a1309, input wire b1309,
  input wire a1310, input wire b1310,
  input wire a1311, input wire b1311,
  input wire a1312, input wire b1312,
  input wire a1313, input wire b1313,
  input wire a1314, input wire b1314,
  input wire a1315, input wire b1315,
  input wire a1316, input wire b1316,
  input wire a1317, input wire b1317,
  input wire a1318, input wire b1318,
  input wire a1319, input wire b1319,
  input wire a1320, input wire b1320,
  input wire a1321, input wire b1321,
  input wire a1322, input wire b1322,
  input wire a1323, input wire b1323,
  input wire a1324, input wire b1324,
  input wire a1325, input wire b1325,
  input wire a1326, input wire b1326,
  input wire a1327, input wire b1327,
  input wire a1328, input wire b1328,
  input wire a1329, input wire b1329,
  input wire a1330, input wire b1330,
  input wire a1331, input wire b1331,
  input wire a1332, input wire b1332,
  input wire a1333, input wire b1333,
  input wire a1334, input wire b1334,
  input wire a1335, input wire b1335,
  input wire a1336, input wire b1336,
  input wire a1337, input wire b1337,
  input wire a1338, input wire b1338,
  input wire a1339, input wire b1339,
  input wire a1340, input wire b1340,
  input wire a1341, input wire b1341,
  input wire a1342, input wire b1342,
  input wire a1343, input wire b1343,
  input wire a1344, input wire b1344,
  input wire a1345, input wire b1345,
  input wire a1346, input wire b1346,
  input wire a1347, input wire b1347,
  input wire a1348, input wire b1348,
  input wire a1349, input wire b1349,
  input wire a1350, input wire b1350,
  input wire a1351, input wire b1351,
  input wire a1352, input wire b1352,
  input wire a1353, input wire b1353,
  input wire a1354, input wire b1354,
  input wire a1355, input wire b1355,
  input wire a1356, input wire b1356,
  input wire a1357, input wire b1357,
  input wire a1358, input wire b1358,
  input wire a1359, input wire b1359,
  input wire a1360, input wire b1360,
  input wire a1361, input wire b1361,
  input wire a1362, input wire b1362,
  input wire a1363, input wire b1363,
  input wire a1364, input wire b1364,
  input wire a1365, input wire b1365,
  input wire a1366, input wire b1366,
  input wire a1367, input wire b1367,
  input wire a1368, input wire b1368,
  input wire a1369, input wire b1369,
  input wire a1370, input wire b1370,
  input wire a1371, input wire b1371,
  input wire a1372, input wire b1372,
  input wire a1373, input wire b1373,
  input wire a1374, input wire b1374,
  input wire a1375, input wire b1375,
  input wire a1376, input wire b1376,
  input wire a1377, input wire b1377,
  input wire a1378, input wire b1378,
  input wire a1379, input wire b1379,
  input wire a1380, input wire b1380,
  input wire a1381, input wire b1381,
  input wire a1382, input wire b1382,
  input wire a1383, input wire b1383,
  input wire a1384, input wire b1384,
  input wire a1385, input wire b1385,
  input wire a1386, input wire b1386,
  input wire a1387, input wire b1387,
  input wire a1388, input wire b1388,
  input wire a1389, input wire b1389,
  input wire a1390, input wire b1390,
  input wire a1391, input wire b1391,
  input wire a1392, input wire b1392,
  input wire a1393, input wire b1393,
  input wire a1394, input wire b1394,
  input wire a1395, input wire b1395,
  input wire a1396, input wire b1396,
  input wire a1397, input wire b1397,
  input wire a1398, input wire b1398,
  input wire a1399, input wire b1399,
  input wire a1400, input wire b1400,
  input wire a1401, input wire b1401,
  input wire a1402, input wire b1402,
  input wire a1403, input wire b1403,
  input wire a1404, input wire b1404,
  input wire a1405, input wire b1405,
  input wire a1406, input wire b1406,
  input wire a1407, input wire b1407,
  input wire a1408, input wire b1408,
  input wire a1409, input wire b1409,
  input wire a1410, input wire b1410,
  input wire a1411, input wire b1411,
  input wire a1412, input wire b1412,
  input wire a1413, input wire b1413,
  input wire a1414, input wire b1414,
  input wire a1415, input wire b1415,
  input wire a1416, input wire b1416,
  input wire a1417, input wire b1417,
  input wire a1418, input wire b1418,
  input wire a1419, input wire b1419,
  input wire a1420, input wire b1420,
  input wire a1421, input wire b1421,
  input wire a1422, input wire b1422,
  input wire a1423, input wire b1423,
  input wire a1424, input wire b1424,
  input wire a1425, input wire b1425,
  input wire a1426, input wire b1426,
  input wire a1427, input wire b1427,
  input wire a1428, input wire b1428,
  input wire a1429, input wire b1429,
  input wire a1430, input wire b1430,
  input wire a1431, input wire b1431,
  input wire a1432, input wire b1432,
  input wire a1433, input wire b1433,
  input wire a1434, input wire b1434,
  input wire a1435, input wire b1435,
  input wire a1436, input wire b1436,
  input wire a1437, input wire b1437,
  input wire a1438, input wire b1438,
  input wire a1439, input wire b1439,
  input wire a1440, input wire b1440,
  input wire a1441, input wire b1441,
  input wire a1442, input wire b1442,
  input wire a1443, input wire b1443,
  input wire a1444, input wire b1444,
  input wire a1445, input wire b1445,
  input wire a1446, input wire b1446,
  input wire a1447, input wire b1447,
  input wire a1448, input wire b1448,
  input wire a1449, input wire b1449,
  input wire a1450, input wire b1450,
  input wire a1451, input wire b1451,
  input wire a1452, input wire b1452,
  input wire a1453, input wire b1453,
  input wire a1454, input wire b1454,
  input wire a1455, input wire b1455,
  input wire a1456, input wire b1456,
  input wire a1457, input wire b1457,
  input wire a1458, input wire b1458,
  input wire a1459, input wire b1459,
  input wire a1460, input wire b1460,
  input wire a1461, input wire b1461,
  input wire a1462, input wire b1462,
  input wire a1463, input wire b1463,
  input wire a1464, input wire b1464,
  input wire a1465, input wire b1465,
  input wire a1466, input wire b1466,
  input wire a1467, input wire b1467,
  input wire a1468, input wire b1468,
  input wire a1469, input wire b1469,
  input wire a1470, input wire b1470,
  input wire a1471, input wire b1471,
  input wire a1472, input wire b1472,
  input wire a1473, input wire b1473,
  input wire a1474, input wire b1474,
  input wire a1475, input wire b1475,
  input wire a1476, input wire b1476,
  input wire a1477, input wire b1477,
  input wire a1478, input wire b1478,
  input wire a1479, input wire b1479,
  input wire a1480, input wire b1480,
  input wire a1481, input wire b1481,
  input wire a1482, input wire b1482,
  input wire a1483, input wire b1483,
  input wire a1484, input wire b1484,
  input wire a1485, input wire b1485,
  input wire a1486, input wire b1486,
  input wire a1487, input wire b1487,
  input wire a1488, input wire b1488,
  input wire a1489, input wire b1489,
  input wire a1490, input wire b1490,
  input wire a1491, input wire b1491,
  input wire a1492, input wire b1492,
  input wire a1493, input wire b1493,
  input wire a1494, input wire b1494,
  input wire a1495, input wire b1495,
  input wire a1496, input wire b1496,
  input wire a1497, input wire b1497,
  input wire a1498, input wire b1498,
  input wire a1499, input wire b1499,
  input wire a1500, input wire b1500,
  input wire a1501, input wire b1501,
  input wire a1502, input wire b1502,
  input wire a1503, input wire b1503,
  input wire a1504, input wire b1504,
  input wire a1505, input wire b1505,
  input wire a1506, input wire b1506,
  input wire a1507, input wire b1507,
  input wire a1508, input wire b1508,
  input wire a1509, input wire b1509,
  input wire a1510, input wire b1510,
  input wire a1511, input wire b1511,
  input wire a1512, input wire b1512,
  input wire a1513, input wire b1513,
  input wire a1514, input wire b1514,
  input wire a1515, input wire b1515,
  input wire a1516, input wire b1516,
  input wire a1517, input wire b1517,
  input wire a1518, input wire b1518,
  input wire a1519, input wire b1519,
  input wire a1520, input wire b1520,
  input wire a1521, input wire b1521,
  input wire a1522, input wire b1522,
  input wire a1523, input wire b1523,
  input wire a1524, input wire b1524,
  input wire a1525, input wire b1525,
  input wire a1526, input wire b1526,
  input wire a1527, input wire b1527,
  input wire a1528, input wire b1528,
  input wire a1529, input wire b1529,
  input wire a1530, input wire b1530,
  input wire a1531, input wire b1531,
  input wire a1532, input wire b1532,
  input wire a1533, input wire b1533,
  input wire a1534, input wire b1534,
  input wire a1535, input wire b1535,
  input wire a1536, input wire b1536,
  input wire a1537, input wire b1537,
  input wire a1538, input wire b1538,
  input wire a1539, input wire b1539,
  input wire a1540, input wire b1540,
  input wire a1541, input wire b1541,
  input wire a1542, input wire b1542,
  input wire a1543, input wire b1543,
  input wire a1544, input wire b1544,
  input wire a1545, input wire b1545,
  input wire a1546, input wire b1546,
  input wire a1547, input wire b1547,
  input wire a1548, input wire b1548,
  input wire a1549, input wire b1549,
  input wire a1550, input wire b1550,
  input wire a1551, input wire b1551,
  input wire a1552, input wire b1552,
  input wire a1553, input wire b1553,
  input wire a1554, input wire b1554,
  input wire a1555, input wire b1555,
  input wire a1556, input wire b1556,
  input wire a1557, input wire b1557,
  input wire a1558, input wire b1558,
  input wire a1559, input wire b1559,
  input wire a1560, input wire b1560,
  input wire a1561, input wire b1561,
  input wire a1562, input wire b1562,
  input wire a1563, input wire b1563,
  input wire a1564, input wire b1564,
  input wire a1565, input wire b1565,
  input wire a1566, input wire b1566,
  input wire a1567, input wire b1567,
  input wire a1568, input wire b1568,
  input wire a1569, input wire b1569,
  input wire a1570, input wire b1570,
  input wire a1571, input wire b1571,
  input wire a1572, input wire b1572,
  input wire a1573, input wire b1573,
  input wire a1574, input wire b1574,
  input wire a1575, input wire b1575,
  input wire a1576, input wire b1576,
  input wire a1577, input wire b1577,
  input wire a1578, input wire b1578,
  input wire a1579, input wire b1579,
  input wire a1580, input wire b1580,
  input wire a1581, input wire b1581,
  input wire a1582, input wire b1582,
  input wire a1583, input wire b1583,
  input wire a1584, input wire b1584,
  input wire a1585, input wire b1585,
  input wire a1586, input wire b1586,
  input wire a1587, input wire b1587,
  input wire a1588, input wire b1588,
  input wire a1589, input wire b1589,
  input wire a1590, input wire b1590,
  input wire a1591, input wire b1591,
  input wire a1592, input wire b1592,
  input wire a1593, input wire b1593,
  input wire a1594, input wire b1594,
  input wire a1595, input wire b1595,
  input wire a1596, input wire b1596,
  input wire a1597, input wire b1597,
  input wire a1598, input wire b1598,
  input wire a1599, input wire b1599,
  input wire a1600, input wire b1600,
  input wire a1601, input wire b1601,
  input wire a1602, input wire b1602,
  input wire a1603, input wire b1603,
  input wire a1604, input wire b1604,
  input wire a1605, input wire b1605,
  input wire a1606, input wire b1606,
  input wire a1607, input wire b1607,
  input wire a1608, input wire b1608,
  input wire a1609, input wire b1609,
  input wire a1610, input wire b1610,
  input wire a1611, input wire b1611,
  input wire a1612, input wire b1612,
  input wire a1613, input wire b1613,
  input wire a1614, input wire b1614,
  input wire a1615, input wire b1615,
  input wire a1616, input wire b1616,
  input wire a1617, input wire b1617,
  input wire a1618, input wire b1618,
  input wire a1619, input wire b1619,
  input wire a1620, input wire b1620,
  input wire a1621, input wire b1621,
  input wire a1622, input wire b1622,
  input wire a1623, input wire b1623,
  input wire a1624, input wire b1624,
  input wire a1625, input wire b1625,
  input wire a1626, input wire b1626,
  input wire a1627, input wire b1627,
  input wire a1628, input wire b1628,
  input wire a1629, input wire b1629,
  input wire a1630, input wire b1630,
  input wire a1631, input wire b1631,
  input wire a1632, input wire b1632,
  input wire a1633, input wire b1633,
  input wire a1634, input wire b1634,
  input wire a1635, input wire b1635,
  input wire a1636, input wire b1636,
  input wire a1637, input wire b1637,
  input wire a1638, input wire b1638,
  input wire a1639, input wire b1639,
  input wire a1640, input wire b1640,
  input wire a1641, input wire b1641,
  input wire a1642, input wire b1642,
  input wire a1643, input wire b1643,
  input wire a1644, input wire b1644,
  input wire a1645, input wire b1645,
  input wire a1646, input wire b1646,
  input wire a1647, input wire b1647,
  input wire a1648, input wire b1648,
  input wire a1649, input wire b1649,
  input wire a1650, input wire b1650,
  input wire a1651, input wire b1651,
  input wire a1652, input wire b1652,
  input wire a1653, input wire b1653,
  input wire a1654, input wire b1654,
  input wire a1655, input wire b1655,
  input wire a1656, input wire b1656,
  input wire a1657, input wire b1657,
  input wire a1658, input wire b1658,
  input wire a1659, input wire b1659,
  input wire a1660, input wire b1660,
  input wire a1661, input wire b1661,
  input wire a1662, input wire b1662,
  input wire a1663, input wire b1663,
  input wire a1664, input wire b1664,
  input wire a1665, input wire b1665,
  input wire a1666, input wire b1666,
  input wire a1667, input wire b1667,
  input wire a1668, input wire b1668,
  input wire a1669, input wire b1669,
  input wire a1670, input wire b1670,
  input wire a1671, input wire b1671,
  input wire a1672, input wire b1672,
  input wire a1673, input wire b1673,
  input wire a1674, input wire b1674,
  input wire a1675, input wire b1675,
  input wire a1676, input wire b1676,
  input wire a1677, input wire b1677,
  input wire a1678, input wire b1678,
  input wire a1679, input wire b1679,
  input wire a1680, input wire b1680,
  input wire a1681, input wire b1681,
  input wire a1682, input wire b1682,
  input wire a1683, input wire b1683,
  input wire a1684, input wire b1684,
  input wire a1685, input wire b1685,
  input wire a1686, input wire b1686,
  input wire a1687, input wire b1687,
  input wire a1688, input wire b1688,
  input wire a1689, input wire b1689,
  input wire a1690, input wire b1690,
  input wire a1691, input wire b1691,
  input wire a1692, input wire b1692,
  input wire a1693, input wire b1693,
  input wire a1694, input wire b1694,
  input wire a1695, input wire b1695,
  input wire a1696, input wire b1696,
  input wire a1697, input wire b1697,
  input wire a1698, input wire b1698,
  input wire a1699, input wire b1699,
  input wire a1700, input wire b1700,
  input wire a1701, input wire b1701,
  input wire a1702, input wire b1702,
  input wire a1703, input wire b1703,
  input wire a1704, input wire b1704,
  input wire a1705, input wire b1705,
  input wire a1706, input wire b1706,
  input wire a1707, input wire b1707,
  input wire a1708, input wire b1708,
  input wire a1709, input wire b1709,
  input wire a1710, input wire b1710,
  input wire a1711, input wire b1711,
  input wire a1712, input wire b1712,
  input wire a1713, input wire b1713,
  input wire a1714, input wire b1714,
  input wire a1715, input wire b1715,
  input wire a1716, input wire b1716,
  input wire a1717, input wire b1717,
  input wire a1718, input wire b1718,
  input wire a1719, input wire b1719,
  input wire a1720, input wire b1720,
  input wire a1721, input wire b1721,
  input wire a1722, input wire b1722,
  input wire a1723, input wire b1723,
  input wire a1724, input wire b1724,
  input wire a1725, input wire b1725,
  input wire a1726, input wire b1726,
  input wire a1727, input wire b1727,
  input wire a1728, input wire b1728,
  input wire a1729, input wire b1729,
  input wire a1730, input wire b1730,
  input wire a1731, input wire b1731,
  input wire a1732, input wire b1732,
  input wire a1733, input wire b1733,
  input wire a1734, input wire b1734,
  input wire a1735, input wire b1735,
  input wire a1736, input wire b1736,
  input wire a1737, input wire b1737,
  input wire a1738, input wire b1738,
  input wire a1739, input wire b1739,
  input wire a1740, input wire b1740,
  input wire a1741, input wire b1741,
  input wire a1742, input wire b1742,
  input wire a1743, input wire b1743,
  input wire a1744, input wire b1744,
  input wire a1745, input wire b1745,
  input wire a1746, input wire b1746,
  input wire a1747, input wire b1747,
  input wire a1748, input wire b1748,
  input wire a1749, input wire b1749,
  input wire a1750, input wire b1750,
  input wire a1751, input wire b1751,
  input wire a1752, input wire b1752,
  input wire a1753, input wire b1753,
  input wire a1754, input wire b1754,
  input wire a1755, input wire b1755,
  input wire a1756, input wire b1756,
  input wire a1757, input wire b1757,
  input wire a1758, input wire b1758,
  input wire a1759, input wire b1759,
  input wire a1760, input wire b1760,
  input wire a1761, input wire b1761,
  input wire a1762, input wire b1762,
  input wire a1763, input wire b1763,
  input wire a1764, input wire b1764,
  input wire a1765, input wire b1765,
  input wire a1766, input wire b1766,
  input wire a1767, input wire b1767,
  input wire a1768, input wire b1768,
  input wire a1769, input wire b1769,
  input wire a1770, input wire b1770,
  input wire a1771, input wire b1771,
  input wire a1772, input wire b1772,
  input wire a1773, input wire b1773,
  input wire a1774, input wire b1774,
  input wire a1775, input wire b1775,
  input wire a1776, input wire b1776,
  input wire a1777, input wire b1777,
  input wire a1778, input wire b1778,
  input wire a1779, input wire b1779,
  input wire a1780, input wire b1780,
  input wire a1781, input wire b1781,
  input wire a1782, input wire b1782,
  input wire a1783, input wire b1783,
  input wire a1784, input wire b1784,
  input wire a1785, input wire b1785,
  input wire a1786, input wire b1786,
  input wire a1787, input wire b1787,
  input wire a1788, input wire b1788,
  input wire a1789, input wire b1789,
  input wire a1790, input wire b1790,
  input wire a1791, input wire b1791,
  input wire a1792, input wire b1792,
  input wire a1793, input wire b1793,
  input wire a1794, input wire b1794,
  input wire a1795, input wire b1795,
  input wire a1796, input wire b1796,
  input wire a1797, input wire b1797,
  input wire a1798, input wire b1798,
  input wire a1799, input wire b1799,
  input wire a1800, input wire b1800,
  input wire a1801, input wire b1801,
  input wire a1802, input wire b1802,
  input wire a1803, input wire b1803,
  input wire a1804, input wire b1804,
  input wire a1805, input wire b1805,
  input wire a1806, input wire b1806,
  input wire a1807, input wire b1807,
  input wire a1808, input wire b1808,
  input wire a1809, input wire b1809,
  input wire a1810, input wire b1810,
  input wire a1811, input wire b1811,
  input wire a1812, input wire b1812,
  input wire a1813, input wire b1813,
  input wire a1814, input wire b1814,
  input wire a1815, input wire b1815,
  input wire a1816, input wire b1816,
  input wire a1817, input wire b1817,
  input wire a1818, input wire b1818,
  input wire a1819, input wire b1819,
  input wire a1820, input wire b1820,
  input wire a1821, input wire b1821,
  input wire a1822, input wire b1822,
  input wire a1823, input wire b1823,
  input wire a1824, input wire b1824,
  input wire a1825, input wire b1825,
  input wire a1826, input wire b1826,
  input wire a1827, input wire b1827,
  input wire a1828, input wire b1828,
  input wire a1829, input wire b1829,
  input wire a1830, input wire b1830,
  input wire a1831, input wire b1831,
  input wire a1832, input wire b1832,
  input wire a1833, input wire b1833,
  input wire a1834, input wire b1834,
  input wire a1835, input wire b1835,
  input wire a1836, input wire b1836,
  input wire a1837, input wire b1837,
  input wire a1838, input wire b1838,
  input wire a1839, input wire b1839,
  input wire a1840, input wire b1840,
  input wire a1841, input wire b1841,
  input wire a1842, input wire b1842,
  input wire a1843, input wire b1843,
  input wire a1844, input wire b1844,
  input wire a1845, input wire b1845,
  input wire a1846, input wire b1846,
  input wire a1847, input wire b1847,
  input wire a1848, input wire b1848,
  input wire a1849, input wire b1849,
  input wire a1850, input wire b1850,
  input wire a1851, input wire b1851,
  input wire a1852, input wire b1852,
  input wire a1853, input wire b1853,
  input wire a1854, input wire b1854,
  input wire a1855, input wire b1855,
  input wire a1856, input wire b1856,
  input wire a1857, input wire b1857,
  input wire a1858, input wire b1858,
  input wire a1859, input wire b1859,
  input wire a1860, input wire b1860,
  input wire a1861, input wire b1861,
  input wire a1862, input wire b1862,
  input wire a1863, input wire b1863,
  input wire a1864, input wire b1864,
  input wire a1865, input wire b1865,
  input wire a1866, input wire b1866,
  input wire a1867, input wire b1867,
  input wire a1868, input wire b1868,
  input wire a1869, input wire b1869,
  input wire a1870, input wire b1870,
  input wire a1871, input wire b1871,
  input wire a1872, input wire b1872,
  input wire a1873, input wire b1873,
  input wire a1874, input wire b1874,
  input wire a1875, input wire b1875,
  input wire a1876, input wire b1876,
  input wire a1877, input wire b1877,
  input wire a1878, input wire b1878,
  input wire a1879, input wire b1879,
  input wire a1880, input wire b1880,
  input wire a1881, input wire b1881,
  input wire a1882, input wire b1882,
  input wire a1883, input wire b1883,
  input wire a1884, input wire b1884,
  input wire a1885, input wire b1885,
  input wire a1886, input wire b1886,
  input wire a1887, input wire b1887,
  input wire a1888, input wire b1888,
  input wire a1889, input wire b1889,
  input wire a1890, input wire b1890,
  input wire a1891, input wire b1891,
  input wire a1892, input wire b1892,
  input wire a1893, input wire b1893,
  input wire a1894, input wire b1894,
  input wire a1895, input wire b1895,
  input wire a1896, input wire b1896,
  input wire a1897, input wire b1897,
  input wire a1898, input wire b1898,
  input wire a1899, input wire b1899,
  input wire a1900, input wire b1900,
  input wire a1901, input wire b1901,
  input wire a1902, input wire b1902,
  input wire a1903, input wire b1903,
  input wire a1904, input wire b1904,
  input wire a1905, input wire b1905,
  input wire a1906, input wire b1906,
  input wire a1907, input wire b1907,
  input wire a1908, input wire b1908,
  input wire a1909, input wire b1909,
  input wire a1910, input wire b1910,
  input wire a1911, input wire b1911,
  input wire a1912, input wire b1912,
  input wire a1913, input wire b1913,
  input wire a1914, input wire b1914,
  input wire a1915, input wire b1915,
  input wire a1916, input wire b1916,
  input wire a1917, input wire b1917,
  input wire a1918, input wire b1918,
  input wire a1919, input wire b1919,
  input wire a1920, input wire b1920,
  input wire a1921, input wire b1921,
  input wire a1922, input wire b1922,
  input wire a1923, input wire b1923,
  input wire a1924, input wire b1924,
  input wire a1925, input wire b1925,
  input wire a1926, input wire b1926,
  input wire a1927, input wire b1927,
  input wire a1928, input wire b1928,
  input wire a1929, input wire b1929,
  input wire a1930, input wire b1930,
  input wire a1931, input wire b1931,
  input wire a1932, input wire b1932,
  input wire a1933, input wire b1933,
  input wire a1934, input wire b1934,
  input wire a1935, input wire b1935,
  input wire a1936, input wire b1936,
  input wire a1937, input wire b1937,
  input wire a1938, input wire b1938,
  input wire a1939, input wire b1939,
  input wire a1940, input wire b1940,
  input wire a1941, input wire b1941,
  input wire a1942, input wire b1942,
  input wire a1943, input wire b1943,
  input wire a1944, input wire b1944,
  input wire a1945, input wire b1945,
  input wire a1946, input wire b1946,
  input wire a1947, input wire b1947,
  input wire a1948, input wire b1948,
  input wire a1949, input wire b1949,
  input wire a1950, input wire b1950,
  input wire a1951, input wire b1951,
  input wire a1952, input wire b1952,
  input wire a1953, input wire b1953,
  input wire a1954, input wire b1954,
  input wire a1955, input wire b1955,
  input wire a1956, input wire b1956,
  input wire a1957, input wire b1957,
  input wire a1958, input wire b1958,
  input wire a1959, input wire b1959,
  input wire a1960, input wire b1960,
  input wire a1961, input wire b1961,
  input wire a1962, input wire b1962,
  input wire a1963, input wire b1963,
  input wire a1964, input wire b1964,
  input wire a1965, input wire b1965,
  input wire a1966, input wire b1966,
  input wire a1967, input wire b1967,
  input wire a1968, input wire b1968,
  input wire a1969, input wire b1969,
  input wire a1970, input wire b1970,
  input wire a1971, input wire b1971,
  input wire a1972, input wire b1972,
  input wire a1973, input wire b1973,
  input wire a1974, input wire b1974,
  input wire a1975, input wire b1975,
  input wire a1976, input wire b1976,
  input wire a1977, input wire b1977,
  input wire a1978, input wire b1978,
  input wire a1979, input wire b1979,
  input wire a1980, input wire b1980,
  input wire a1981, input wire b1981,
  input wire a1982, input wire b1982,
  input wire a1983, input wire b1983,
  input wire a1984, input wire b1984,
  input wire a1985, input wire b1985,
  input wire a1986, input wire b1986,
  input wire a1987, input wire b1987,
  input wire a1988, input wire b1988,
  input wire a1989, input wire b1989,
  input wire a1990, input wire b1990,
  input wire a1991, input wire b1991,
  input wire a1992, input wire b1992,
  input wire a1993, input wire b1993,
  input wire a1994, input wire b1994,
  input wire a1995, input wire b1995,
  input wire a1996, input wire b1996,
  input wire a1997, input wire b1997,
  input wire a1998, input wire b1998,
  input wire a1999, input wire b1999,
  input wire a2000, input wire b2000,
  input wire a2001, input wire b2001,
  input wire a2002, input wire b2002,
  input wire a2003, input wire b2003,
  input wire a2004, input wire b2004,
  input wire a2005, input wire b2005,
  input wire a2006, input wire b2006,
  input wire a2007, input wire b2007,
  input wire a2008, input wire b2008,
  input wire a2009, input wire b2009,
  input wire a2010, input wire b2010,
  input wire a2011, input wire b2011,
  input wire a2012, input wire b2012,
  input wire a2013, input wire b2013,
  input wire a2014, input wire b2014,
  input wire a2015, input wire b2015,
  input wire a2016, input wire b2016,
  input wire a2017, input wire b2017,
  input wire a2018, input wire b2018,
  input wire a2019, input wire b2019,
  input wire a2020, input wire b2020,
  input wire a2021, input wire b2021,
  input wire a2022, input wire b2022,
  input wire a2023, input wire b2023,
  input wire a2024, input wire b2024,
  input wire a2025, input wire b2025,
  input wire a2026, input wire b2026,
  input wire a2027, input wire b2027,
  input wire a2028, input wire b2028,
  input wire a2029, input wire b2029,
  input wire a2030, input wire b2030,
  input wire a2031, input wire b2031,
  input wire a2032, input wire b2032,
  input wire a2033, input wire b2033,
  input wire a2034, input wire b2034,
  input wire a2035, input wire b2035,
  input wire a2036, input wire b2036,
  input wire a2037, input wire b2037,
  input wire a2038, input wire b2038,
  input wire a2039, input wire b2039,
  input wire a2040, input wire b2040,
  input wire a2041, input wire b2041,
  input wire a2042, input wire b2042,
  input wire a2043, input wire b2043,
  input wire a2044, input wire b2044,
  input wire a2045, input wire b2045,
  input wire a2046, input wire b2046,
  input wire a2047, input wire b2047,
  input wire op0,
  input wire op1,
  output wire y0,
  output wire y1,
  output wire y2,
  output wire y3,
  output wire y4,
  output wire y5,
  output wire y6,
  output wire y7,
  output wire y8,
  output wire y9,
  output wire y10,
  output wire y11,
  output wire y12,
  output wire y13,
  output wire y14,
  output wire y15,
  output wire y16,
  output wire y17,
  output wire y18,
  output wire y19,
  output wire y20,
  output wire y21,
  output wire y22,
  output wire y23,
  output wire y24,
  output wire y25,
  output wire y26,
  output wire y27,
  output wire y28,
  output wire y29,
  output wire y30,
  output wire y31,
  output wire y32,
  output wire y33,
  output wire y34,
  output wire y35,
  output wire y36,
  output wire y37,
  output wire y38,
  output wire y39,
  output wire y40,
  output wire y41,
  output wire y42,
  output wire y43,
  output wire y44,
  output wire y45,
  output wire y46,
  output wire y47,
  output wire y48,
  output wire y49,
  output wire y50,
  output wire y51,
  output wire y52,
  output wire y53,
  output wire y54,
  output wire y55,
  output wire y56,
  output wire y57,
  output wire y58,
  output wire y59,
  output wire y60,
  output wire y61,
  output wire y62,
  output wire y63,
  output wire y64,
  output wire y65,
  output wire y66,
  output wire y67,
  output wire y68,
  output wire y69,
  output wire y70,
  output wire y71,
  output wire y72,
  output wire y73,
  output wire y74,
  output wire y75,
  output wire y76,
  output wire y77,
  output wire y78,
  output wire y79,
  output wire y80,
  output wire y81,
  output wire y82,
  output wire y83,
  output wire y84,
  output wire y85,
  output wire y86,
  output wire y87,
  output wire y88,
  output wire y89,
  output wire y90,
  output wire y91,
  output wire y92,
  output wire y93,
  output wire y94,
  output wire y95,
  output wire y96,
  output wire y97,
  output wire y98,
  output wire y99,
  output wire y100,
  output wire y101,
  output wire y102,
  output wire y103,
  output wire y104,
  output wire y105,
  output wire y106,
  output wire y107,
  output wire y108,
  output wire y109,
  output wire y110,
  output wire y111,
  output wire y112,
  output wire y113,
  output wire y114,
  output wire y115,
  output wire y116,
  output wire y117,
  output wire y118,
  output wire y119,
  output wire y120,
  output wire y121,
  output wire y122,
  output wire y123,
  output wire y124,
  output wire y125,
  output wire y126,
  output wire y127,
  output wire y128,
  output wire y129,
  output wire y130,
  output wire y131,
  output wire y132,
  output wire y133,
  output wire y134,
  output wire y135,
  output wire y136,
  output wire y137,
  output wire y138,
  output wire y139,
  output wire y140,
  output wire y141,
  output wire y142,
  output wire y143,
  output wire y144,
  output wire y145,
  output wire y146,
  output wire y147,
  output wire y148,
  output wire y149,
  output wire y150,
  output wire y151,
  output wire y152,
  output wire y153,
  output wire y154,
  output wire y155,
  output wire y156,
  output wire y157,
  output wire y158,
  output wire y159,
  output wire y160,
  output wire y161,
  output wire y162,
  output wire y163,
  output wire y164,
  output wire y165,
  output wire y166,
  output wire y167,
  output wire y168,
  output wire y169,
  output wire y170,
  output wire y171,
  output wire y172,
  output wire y173,
  output wire y174,
  output wire y175,
  output wire y176,
  output wire y177,
  output wire y178,
  output wire y179,
  output wire y180,
  output wire y181,
  output wire y182,
  output wire y183,
  output wire y184,
  output wire y185,
  output wire y186,
  output wire y187,
  output wire y188,
  output wire y189,
  output wire y190,
  output wire y191,
  output wire y192,
  output wire y193,
  output wire y194,
  output wire y195,
  output wire y196,
  output wire y197,
  output wire y198,
  output wire y199,
  output wire y200,
  output wire y201,
  output wire y202,
  output wire y203,
  output wire y204,
  output wire y205,
  output wire y206,
  output wire y207,
  output wire y208,
  output wire y209,
  output wire y210,
  output wire y211,
  output wire y212,
  output wire y213,
  output wire y214,
  output wire y215,
  output wire y216,
  output wire y217,
  output wire y218,
  output wire y219,
  output wire y220,
  output wire y221,
  output wire y222,
  output wire y223,
  output wire y224,
  output wire y225,
  output wire y226,
  output wire y227,
  output wire y228,
  output wire y229,
  output wire y230,
  output wire y231,
  output wire y232,
  output wire y233,
  output wire y234,
  output wire y235,
  output wire y236,
  output wire y237,
  output wire y238,
  output wire y239,
  output wire y240,
  output wire y241,
  output wire y242,
  output wire y243,
  output wire y244,
  output wire y245,
  output wire y246,
  output wire y247,
  output wire y248,
  output wire y249,
  output wire y250,
  output wire y251,
  output wire y252,
  output wire y253,
  output wire y254,
  output wire y255,
  output wire y256,
  output wire y257,
  output wire y258,
  output wire y259,
  output wire y260,
  output wire y261,
  output wire y262,
  output wire y263,
  output wire y264,
  output wire y265,
  output wire y266,
  output wire y267,
  output wire y268,
  output wire y269,
  output wire y270,
  output wire y271,
  output wire y272,
  output wire y273,
  output wire y274,
  output wire y275,
  output wire y276,
  output wire y277,
  output wire y278,
  output wire y279,
  output wire y280,
  output wire y281,
  output wire y282,
  output wire y283,
  output wire y284,
  output wire y285,
  output wire y286,
  output wire y287,
  output wire y288,
  output wire y289,
  output wire y290,
  output wire y291,
  output wire y292,
  output wire y293,
  output wire y294,
  output wire y295,
  output wire y296,
  output wire y297,
  output wire y298,
  output wire y299,
  output wire y300,
  output wire y301,
  output wire y302,
  output wire y303,
  output wire y304,
  output wire y305,
  output wire y306,
  output wire y307,
  output wire y308,
  output wire y309,
  output wire y310,
  output wire y311,
  output wire y312,
  output wire y313,
  output wire y314,
  output wire y315,
  output wire y316,
  output wire y317,
  output wire y318,
  output wire y319,
  output wire y320,
  output wire y321,
  output wire y322,
  output wire y323,
  output wire y324,
  output wire y325,
  output wire y326,
  output wire y327,
  output wire y328,
  output wire y329,
  output wire y330,
  output wire y331,
  output wire y332,
  output wire y333,
  output wire y334,
  output wire y335,
  output wire y336,
  output wire y337,
  output wire y338,
  output wire y339,
  output wire y340,
  output wire y341,
  output wire y342,
  output wire y343,
  output wire y344,
  output wire y345,
  output wire y346,
  output wire y347,
  output wire y348,
  output wire y349,
  output wire y350,
  output wire y351,
  output wire y352,
  output wire y353,
  output wire y354,
  output wire y355,
  output wire y356,
  output wire y357,
  output wire y358,
  output wire y359,
  output wire y360,
  output wire y361,
  output wire y362,
  output wire y363,
  output wire y364,
  output wire y365,
  output wire y366,
  output wire y367,
  output wire y368,
  output wire y369,
  output wire y370,
  output wire y371,
  output wire y372,
  output wire y373,
  output wire y374,
  output wire y375,
  output wire y376,
  output wire y377,
  output wire y378,
  output wire y379,
  output wire y380,
  output wire y381,
  output wire y382,
  output wire y383,
  output wire y384,
  output wire y385,
  output wire y386,
  output wire y387,
  output wire y388,
  output wire y389,
  output wire y390,
  output wire y391,
  output wire y392,
  output wire y393,
  output wire y394,
  output wire y395,
  output wire y396,
  output wire y397,
  output wire y398,
  output wire y399,
  output wire y400,
  output wire y401,
  output wire y402,
  output wire y403,
  output wire y404,
  output wire y405,
  output wire y406,
  output wire y407,
  output wire y408,
  output wire y409,
  output wire y410,
  output wire y411,
  output wire y412,
  output wire y413,
  output wire y414,
  output wire y415,
  output wire y416,
  output wire y417,
  output wire y418,
  output wire y419,
  output wire y420,
  output wire y421,
  output wire y422,
  output wire y423,
  output wire y424,
  output wire y425,
  output wire y426,
  output wire y427,
  output wire y428,
  output wire y429,
  output wire y430,
  output wire y431,
  output wire y432,
  output wire y433,
  output wire y434,
  output wire y435,
  output wire y436,
  output wire y437,
  output wire y438,
  output wire y439,
  output wire y440,
  output wire y441,
  output wire y442,
  output wire y443,
  output wire y444,
  output wire y445,
  output wire y446,
  output wire y447,
  output wire y448,
  output wire y449,
  output wire y450,
  output wire y451,
  output wire y452,
  output wire y453,
  output wire y454,
  output wire y455,
  output wire y456,
  output wire y457,
  output wire y458,
  output wire y459,
  output wire y460,
  output wire y461,
  output wire y462,
  output wire y463,
  output wire y464,
  output wire y465,
  output wire y466,
  output wire y467,
  output wire y468,
  output wire y469,
  output wire y470,
  output wire y471,
  output wire y472,
  output wire y473,
  output wire y474,
  output wire y475,
  output wire y476,
  output wire y477,
  output wire y478,
  output wire y479,
  output wire y480,
  output wire y481,
  output wire y482,
  output wire y483,
  output wire y484,
  output wire y485,
  output wire y486,
  output wire y487,
  output wire y488,
  output wire y489,
  output wire y490,
  output wire y491,
  output wire y492,
  output wire y493,
  output wire y494,
  output wire y495,
  output wire y496,
  output wire y497,
  output wire y498,
  output wire y499,
  output wire y500,
  output wire y501,
  output wire y502,
  output wire y503,
  output wire y504,
  output wire y505,
  output wire y506,
  output wire y507,
  output wire y508,
  output wire y509,
  output wire y510,
  output wire y511,
  output wire y512,
  output wire y513,
  output wire y514,
  output wire y515,
  output wire y516,
  output wire y517,
  output wire y518,
  output wire y519,
  output wire y520,
  output wire y521,
  output wire y522,
  output wire y523,
  output wire y524,
  output wire y525,
  output wire y526,
  output wire y527,
  output wire y528,
  output wire y529,
  output wire y530,
  output wire y531,
  output wire y532,
  output wire y533,
  output wire y534,
  output wire y535,
  output wire y536,
  output wire y537,
  output wire y538,
  output wire y539,
  output wire y540,
  output wire y541,
  output wire y542,
  output wire y543,
  output wire y544,
  output wire y545,
  output wire y546,
  output wire y547,
  output wire y548,
  output wire y549,
  output wire y550,
  output wire y551,
  output wire y552,
  output wire y553,
  output wire y554,
  output wire y555,
  output wire y556,
  output wire y557,
  output wire y558,
  output wire y559,
  output wire y560,
  output wire y561,
  output wire y562,
  output wire y563,
  output wire y564,
  output wire y565,
  output wire y566,
  output wire y567,
  output wire y568,
  output wire y569,
  output wire y570,
  output wire y571,
  output wire y572,
  output wire y573,
  output wire y574,
  output wire y575,
  output wire y576,
  output wire y577,
  output wire y578,
  output wire y579,
  output wire y580,
  output wire y581,
  output wire y582,
  output wire y583,
  output wire y584,
  output wire y585,
  output wire y586,
  output wire y587,
  output wire y588,
  output wire y589,
  output wire y590,
  output wire y591,
  output wire y592,
  output wire y593,
  output wire y594,
  output wire y595,
  output wire y596,
  output wire y597,
  output wire y598,
  output wire y599,
  output wire y600,
  output wire y601,
  output wire y602,
  output wire y603,
  output wire y604,
  output wire y605,
  output wire y606,
  output wire y607,
  output wire y608,
  output wire y609,
  output wire y610,
  output wire y611,
  output wire y612,
  output wire y613,
  output wire y614,
  output wire y615,
  output wire y616,
  output wire y617,
  output wire y618,
  output wire y619,
  output wire y620,
  output wire y621,
  output wire y622,
  output wire y623,
  output wire y624,
  output wire y625,
  output wire y626,
  output wire y627,
  output wire y628,
  output wire y629,
  output wire y630,
  output wire y631,
  output wire y632,
  output wire y633,
  output wire y634,
  output wire y635,
  output wire y636,
  output wire y637,
  output wire y638,
  output wire y639,
  output wire y640,
  output wire y641,
  output wire y642,
  output wire y643,
  output wire y644,
  output wire y645,
  output wire y646,
  output wire y647,
  output wire y648,
  output wire y649,
  output wire y650,
  output wire y651,
  output wire y652,
  output wire y653,
  output wire y654,
  output wire y655,
  output wire y656,
  output wire y657,
  output wire y658,
  output wire y659,
  output wire y660,
  output wire y661,
  output wire y662,
  output wire y663,
  output wire y664,
  output wire y665,
  output wire y666,
  output wire y667,
  output wire y668,
  output wire y669,
  output wire y670,
  output wire y671,
  output wire y672,
  output wire y673,
  output wire y674,
  output wire y675,
  output wire y676,
  output wire y677,
  output wire y678,
  output wire y679,
  output wire y680,
  output wire y681,
  output wire y682,
  output wire y683,
  output wire y684,
  output wire y685,
  output wire y686,
  output wire y687,
  output wire y688,
  output wire y689,
  output wire y690,
  output wire y691,
  output wire y692,
  output wire y693,
  output wire y694,
  output wire y695,
  output wire y696,
  output wire y697,
  output wire y698,
  output wire y699,
  output wire y700,
  output wire y701,
  output wire y702,
  output wire y703,
  output wire y704,
  output wire y705,
  output wire y706,
  output wire y707,
  output wire y708,
  output wire y709,
  output wire y710,
  output wire y711,
  output wire y712,
  output wire y713,
  output wire y714,
  output wire y715,
  output wire y716,
  output wire y717,
  output wire y718,
  output wire y719,
  output wire y720,
  output wire y721,
  output wire y722,
  output wire y723,
  output wire y724,
  output wire y725,
  output wire y726,
  output wire y727,
  output wire y728,
  output wire y729,
  output wire y730,
  output wire y731,
  output wire y732,
  output wire y733,
  output wire y734,
  output wire y735,
  output wire y736,
  output wire y737,
  output wire y738,
  output wire y739,
  output wire y740,
  output wire y741,
  output wire y742,
  output wire y743,
  output wire y744,
  output wire y745,
  output wire y746,
  output wire y747,
  output wire y748,
  output wire y749,
  output wire y750,
  output wire y751,
  output wire y752,
  output wire y753,
  output wire y754,
  output wire y755,
  output wire y756,
  output wire y757,
  output wire y758,
  output wire y759,
  output wire y760,
  output wire y761,
  output wire y762,
  output wire y763,
  output wire y764,
  output wire y765,
  output wire y766,
  output wire y767,
  output wire y768,
  output wire y769,
  output wire y770,
  output wire y771,
  output wire y772,
  output wire y773,
  output wire y774,
  output wire y775,
  output wire y776,
  output wire y777,
  output wire y778,
  output wire y779,
  output wire y780,
  output wire y781,
  output wire y782,
  output wire y783,
  output wire y784,
  output wire y785,
  output wire y786,
  output wire y787,
  output wire y788,
  output wire y789,
  output wire y790,
  output wire y791,
  output wire y792,
  output wire y793,
  output wire y794,
  output wire y795,
  output wire y796,
  output wire y797,
  output wire y798,
  output wire y799,
  output wire y800,
  output wire y801,
  output wire y802,
  output wire y803,
  output wire y804,
  output wire y805,
  output wire y806,
  output wire y807,
  output wire y808,
  output wire y809,
  output wire y810,
  output wire y811,
  output wire y812,
  output wire y813,
  output wire y814,
  output wire y815,
  output wire y816,
  output wire y817,
  output wire y818,
  output wire y819,
  output wire y820,
  output wire y821,
  output wire y822,
  output wire y823,
  output wire y824,
  output wire y825,
  output wire y826,
  output wire y827,
  output wire y828,
  output wire y829,
  output wire y830,
  output wire y831,
  output wire y832,
  output wire y833,
  output wire y834,
  output wire y835,
  output wire y836,
  output wire y837,
  output wire y838,
  output wire y839,
  output wire y840,
  output wire y841,
  output wire y842,
  output wire y843,
  output wire y844,
  output wire y845,
  output wire y846,
  output wire y847,
  output wire y848,
  output wire y849,
  output wire y850,
  output wire y851,
  output wire y852,
  output wire y853,
  output wire y854,
  output wire y855,
  output wire y856,
  output wire y857,
  output wire y858,
  output wire y859,
  output wire y860,
  output wire y861,
  output wire y862,
  output wire y863,
  output wire y864,
  output wire y865,
  output wire y866,
  output wire y867,
  output wire y868,
  output wire y869,
  output wire y870,
  output wire y871,
  output wire y872,
  output wire y873,
  output wire y874,
  output wire y875,
  output wire y876,
  output wire y877,
  output wire y878,
  output wire y879,
  output wire y880,
  output wire y881,
  output wire y882,
  output wire y883,
  output wire y884,
  output wire y885,
  output wire y886,
  output wire y887,
  output wire y888,
  output wire y889,
  output wire y890,
  output wire y891,
  output wire y892,
  output wire y893,
  output wire y894,
  output wire y895,
  output wire y896,
  output wire y897,
  output wire y898,
  output wire y899,
  output wire y900,
  output wire y901,
  output wire y902,
  output wire y903,
  output wire y904,
  output wire y905,
  output wire y906,
  output wire y907,
  output wire y908,
  output wire y909,
  output wire y910,
  output wire y911,
  output wire y912,
  output wire y913,
  output wire y914,
  output wire y915,
  output wire y916,
  output wire y917,
  output wire y918,
  output wire y919,
  output wire y920,
  output wire y921,
  output wire y922,
  output wire y923,
  output wire y924,
  output wire y925,
  output wire y926,
  output wire y927,
  output wire y928,
  output wire y929,
  output wire y930,
  output wire y931,
  output wire y932,
  output wire y933,
  output wire y934,
  output wire y935,
  output wire y936,
  output wire y937,
  output wire y938,
  output wire y939,
  output wire y940,
  output wire y941,
  output wire y942,
  output wire y943,
  output wire y944,
  output wire y945,
  output wire y946,
  output wire y947,
  output wire y948,
  output wire y949,
  output wire y950,
  output wire y951,
  output wire y952,
  output wire y953,
  output wire y954,
  output wire y955,
  output wire y956,
  output wire y957,
  output wire y958,
  output wire y959,
  output wire y960,
  output wire y961,
  output wire y962,
  output wire y963,
  output wire y964,
  output wire y965,
  output wire y966,
  output wire y967,
  output wire y968,
  output wire y969,
  output wire y970,
  output wire y971,
  output wire y972,
  output wire y973,
  output wire y974,
  output wire y975,
  output wire y976,
  output wire y977,
  output wire y978,
  output wire y979,
  output wire y980,
  output wire y981,
  output wire y982,
  output wire y983,
  output wire y984,
  output wire y985,
  output wire y986,
  output wire y987,
  output wire y988,
  output wire y989,
  output wire y990,
  output wire y991,
  output wire y992,
  output wire y993,
  output wire y994,
  output wire y995,
  output wire y996,
  output wire y997,
  output wire y998,
  output wire y999,
  output wire y1000,
  output wire y1001,
  output wire y1002,
  output wire y1003,
  output wire y1004,
  output wire y1005,
  output wire y1006,
  output wire y1007,
  output wire y1008,
  output wire y1009,
  output wire y1010,
  output wire y1011,
  output wire y1012,
  output wire y1013,
  output wire y1014,
  output wire y1015,
  output wire y1016,
  output wire y1017,
  output wire y1018,
  output wire y1019,
  output wire y1020,
  output wire y1021,
  output wire y1022,
  output wire y1023,
  output wire y1024,
  output wire y1025,
  output wire y1026,
  output wire y1027,
  output wire y1028,
  output wire y1029,
  output wire y1030,
  output wire y1031,
  output wire y1032,
  output wire y1033,
  output wire y1034,
  output wire y1035,
  output wire y1036,
  output wire y1037,
  output wire y1038,
  output wire y1039,
  output wire y1040,
  output wire y1041,
  output wire y1042,
  output wire y1043,
  output wire y1044,
  output wire y1045,
  output wire y1046,
  output wire y1047,
  output wire y1048,
  output wire y1049,
  output wire y1050,
  output wire y1051,
  output wire y1052,
  output wire y1053,
  output wire y1054,
  output wire y1055,
  output wire y1056,
  output wire y1057,
  output wire y1058,
  output wire y1059,
  output wire y1060,
  output wire y1061,
  output wire y1062,
  output wire y1063,
  output wire y1064,
  output wire y1065,
  output wire y1066,
  output wire y1067,
  output wire y1068,
  output wire y1069,
  output wire y1070,
  output wire y1071,
  output wire y1072,
  output wire y1073,
  output wire y1074,
  output wire y1075,
  output wire y1076,
  output wire y1077,
  output wire y1078,
  output wire y1079,
  output wire y1080,
  output wire y1081,
  output wire y1082,
  output wire y1083,
  output wire y1084,
  output wire y1085,
  output wire y1086,
  output wire y1087,
  output wire y1088,
  output wire y1089,
  output wire y1090,
  output wire y1091,
  output wire y1092,
  output wire y1093,
  output wire y1094,
  output wire y1095,
  output wire y1096,
  output wire y1097,
  output wire y1098,
  output wire y1099,
  output wire y1100,
  output wire y1101,
  output wire y1102,
  output wire y1103,
  output wire y1104,
  output wire y1105,
  output wire y1106,
  output wire y1107,
  output wire y1108,
  output wire y1109,
  output wire y1110,
  output wire y1111,
  output wire y1112,
  output wire y1113,
  output wire y1114,
  output wire y1115,
  output wire y1116,
  output wire y1117,
  output wire y1118,
  output wire y1119,
  output wire y1120,
  output wire y1121,
  output wire y1122,
  output wire y1123,
  output wire y1124,
  output wire y1125,
  output wire y1126,
  output wire y1127,
  output wire y1128,
  output wire y1129,
  output wire y1130,
  output wire y1131,
  output wire y1132,
  output wire y1133,
  output wire y1134,
  output wire y1135,
  output wire y1136,
  output wire y1137,
  output wire y1138,
  output wire y1139,
  output wire y1140,
  output wire y1141,
  output wire y1142,
  output wire y1143,
  output wire y1144,
  output wire y1145,
  output wire y1146,
  output wire y1147,
  output wire y1148,
  output wire y1149,
  output wire y1150,
  output wire y1151,
  output wire y1152,
  output wire y1153,
  output wire y1154,
  output wire y1155,
  output wire y1156,
  output wire y1157,
  output wire y1158,
  output wire y1159,
  output wire y1160,
  output wire y1161,
  output wire y1162,
  output wire y1163,
  output wire y1164,
  output wire y1165,
  output wire y1166,
  output wire y1167,
  output wire y1168,
  output wire y1169,
  output wire y1170,
  output wire y1171,
  output wire y1172,
  output wire y1173,
  output wire y1174,
  output wire y1175,
  output wire y1176,
  output wire y1177,
  output wire y1178,
  output wire y1179,
  output wire y1180,
  output wire y1181,
  output wire y1182,
  output wire y1183,
  output wire y1184,
  output wire y1185,
  output wire y1186,
  output wire y1187,
  output wire y1188,
  output wire y1189,
  output wire y1190,
  output wire y1191,
  output wire y1192,
  output wire y1193,
  output wire y1194,
  output wire y1195,
  output wire y1196,
  output wire y1197,
  output wire y1198,
  output wire y1199,
  output wire y1200,
  output wire y1201,
  output wire y1202,
  output wire y1203,
  output wire y1204,
  output wire y1205,
  output wire y1206,
  output wire y1207,
  output wire y1208,
  output wire y1209,
  output wire y1210,
  output wire y1211,
  output wire y1212,
  output wire y1213,
  output wire y1214,
  output wire y1215,
  output wire y1216,
  output wire y1217,
  output wire y1218,
  output wire y1219,
  output wire y1220,
  output wire y1221,
  output wire y1222,
  output wire y1223,
  output wire y1224,
  output wire y1225,
  output wire y1226,
  output wire y1227,
  output wire y1228,
  output wire y1229,
  output wire y1230,
  output wire y1231,
  output wire y1232,
  output wire y1233,
  output wire y1234,
  output wire y1235,
  output wire y1236,
  output wire y1237,
  output wire y1238,
  output wire y1239,
  output wire y1240,
  output wire y1241,
  output wire y1242,
  output wire y1243,
  output wire y1244,
  output wire y1245,
  output wire y1246,
  output wire y1247,
  output wire y1248,
  output wire y1249,
  output wire y1250,
  output wire y1251,
  output wire y1252,
  output wire y1253,
  output wire y1254,
  output wire y1255,
  output wire y1256,
  output wire y1257,
  output wire y1258,
  output wire y1259,
  output wire y1260,
  output wire y1261,
  output wire y1262,
  output wire y1263,
  output wire y1264,
  output wire y1265,
  output wire y1266,
  output wire y1267,
  output wire y1268,
  output wire y1269,
  output wire y1270,
  output wire y1271,
  output wire y1272,
  output wire y1273,
  output wire y1274,
  output wire y1275,
  output wire y1276,
  output wire y1277,
  output wire y1278,
  output wire y1279,
  output wire y1280,
  output wire y1281,
  output wire y1282,
  output wire y1283,
  output wire y1284,
  output wire y1285,
  output wire y1286,
  output wire y1287,
  output wire y1288,
  output wire y1289,
  output wire y1290,
  output wire y1291,
  output wire y1292,
  output wire y1293,
  output wire y1294,
  output wire y1295,
  output wire y1296,
  output wire y1297,
  output wire y1298,
  output wire y1299,
  output wire y1300,
  output wire y1301,
  output wire y1302,
  output wire y1303,
  output wire y1304,
  output wire y1305,
  output wire y1306,
  output wire y1307,
  output wire y1308,
  output wire y1309,
  output wire y1310,
  output wire y1311,
  output wire y1312,
  output wire y1313,
  output wire y1314,
  output wire y1315,
  output wire y1316,
  output wire y1317,
  output wire y1318,
  output wire y1319,
  output wire y1320,
  output wire y1321,
  output wire y1322,
  output wire y1323,
  output wire y1324,
  output wire y1325,
  output wire y1326,
  output wire y1327,
  output wire y1328,
  output wire y1329,
  output wire y1330,
  output wire y1331,
  output wire y1332,
  output wire y1333,
  output wire y1334,
  output wire y1335,
  output wire y1336,
  output wire y1337,
  output wire y1338,
  output wire y1339,
  output wire y1340,
  output wire y1341,
  output wire y1342,
  output wire y1343,
  output wire y1344,
  output wire y1345,
  output wire y1346,
  output wire y1347,
  output wire y1348,
  output wire y1349,
  output wire y1350,
  output wire y1351,
  output wire y1352,
  output wire y1353,
  output wire y1354,
  output wire y1355,
  output wire y1356,
  output wire y1357,
  output wire y1358,
  output wire y1359,
  output wire y1360,
  output wire y1361,
  output wire y1362,
  output wire y1363,
  output wire y1364,
  output wire y1365,
  output wire y1366,
  output wire y1367,
  output wire y1368,
  output wire y1369,
  output wire y1370,
  output wire y1371,
  output wire y1372,
  output wire y1373,
  output wire y1374,
  output wire y1375,
  output wire y1376,
  output wire y1377,
  output wire y1378,
  output wire y1379,
  output wire y1380,
  output wire y1381,
  output wire y1382,
  output wire y1383,
  output wire y1384,
  output wire y1385,
  output wire y1386,
  output wire y1387,
  output wire y1388,
  output wire y1389,
  output wire y1390,
  output wire y1391,
  output wire y1392,
  output wire y1393,
  output wire y1394,
  output wire y1395,
  output wire y1396,
  output wire y1397,
  output wire y1398,
  output wire y1399,
  output wire y1400,
  output wire y1401,
  output wire y1402,
  output wire y1403,
  output wire y1404,
  output wire y1405,
  output wire y1406,
  output wire y1407,
  output wire y1408,
  output wire y1409,
  output wire y1410,
  output wire y1411,
  output wire y1412,
  output wire y1413,
  output wire y1414,
  output wire y1415,
  output wire y1416,
  output wire y1417,
  output wire y1418,
  output wire y1419,
  output wire y1420,
  output wire y1421,
  output wire y1422,
  output wire y1423,
  output wire y1424,
  output wire y1425,
  output wire y1426,
  output wire y1427,
  output wire y1428,
  output wire y1429,
  output wire y1430,
  output wire y1431,
  output wire y1432,
  output wire y1433,
  output wire y1434,
  output wire y1435,
  output wire y1436,
  output wire y1437,
  output wire y1438,
  output wire y1439,
  output wire y1440,
  output wire y1441,
  output wire y1442,
  output wire y1443,
  output wire y1444,
  output wire y1445,
  output wire y1446,
  output wire y1447,
  output wire y1448,
  output wire y1449,
  output wire y1450,
  output wire y1451,
  output wire y1452,
  output wire y1453,
  output wire y1454,
  output wire y1455,
  output wire y1456,
  output wire y1457,
  output wire y1458,
  output wire y1459,
  output wire y1460,
  output wire y1461,
  output wire y1462,
  output wire y1463,
  output wire y1464,
  output wire y1465,
  output wire y1466,
  output wire y1467,
  output wire y1468,
  output wire y1469,
  output wire y1470,
  output wire y1471,
  output wire y1472,
  output wire y1473,
  output wire y1474,
  output wire y1475,
  output wire y1476,
  output wire y1477,
  output wire y1478,
  output wire y1479,
  output wire y1480,
  output wire y1481,
  output wire y1482,
  output wire y1483,
  output wire y1484,
  output wire y1485,
  output wire y1486,
  output wire y1487,
  output wire y1488,
  output wire y1489,
  output wire y1490,
  output wire y1491,
  output wire y1492,
  output wire y1493,
  output wire y1494,
  output wire y1495,
  output wire y1496,
  output wire y1497,
  output wire y1498,
  output wire y1499,
  output wire y1500,
  output wire y1501,
  output wire y1502,
  output wire y1503,
  output wire y1504,
  output wire y1505,
  output wire y1506,
  output wire y1507,
  output wire y1508,
  output wire y1509,
  output wire y1510,
  output wire y1511,
  output wire y1512,
  output wire y1513,
  output wire y1514,
  output wire y1515,
  output wire y1516,
  output wire y1517,
  output wire y1518,
  output wire y1519,
  output wire y1520,
  output wire y1521,
  output wire y1522,
  output wire y1523,
  output wire y1524,
  output wire y1525,
  output wire y1526,
  output wire y1527,
  output wire y1528,
  output wire y1529,
  output wire y1530,
  output wire y1531,
  output wire y1532,
  output wire y1533,
  output wire y1534,
  output wire y1535,
  output wire y1536,
  output wire y1537,
  output wire y1538,
  output wire y1539,
  output wire y1540,
  output wire y1541,
  output wire y1542,
  output wire y1543,
  output wire y1544,
  output wire y1545,
  output wire y1546,
  output wire y1547,
  output wire y1548,
  output wire y1549,
  output wire y1550,
  output wire y1551,
  output wire y1552,
  output wire y1553,
  output wire y1554,
  output wire y1555,
  output wire y1556,
  output wire y1557,
  output wire y1558,
  output wire y1559,
  output wire y1560,
  output wire y1561,
  output wire y1562,
  output wire y1563,
  output wire y1564,
  output wire y1565,
  output wire y1566,
  output wire y1567,
  output wire y1568,
  output wire y1569,
  output wire y1570,
  output wire y1571,
  output wire y1572,
  output wire y1573,
  output wire y1574,
  output wire y1575,
  output wire y1576,
  output wire y1577,
  output wire y1578,
  output wire y1579,
  output wire y1580,
  output wire y1581,
  output wire y1582,
  output wire y1583,
  output wire y1584,
  output wire y1585,
  output wire y1586,
  output wire y1587,
  output wire y1588,
  output wire y1589,
  output wire y1590,
  output wire y1591,
  output wire y1592,
  output wire y1593,
  output wire y1594,
  output wire y1595,
  output wire y1596,
  output wire y1597,
  output wire y1598,
  output wire y1599,
  output wire y1600,
  output wire y1601,
  output wire y1602,
  output wire y1603,
  output wire y1604,
  output wire y1605,
  output wire y1606,
  output wire y1607,
  output wire y1608,
  output wire y1609,
  output wire y1610,
  output wire y1611,
  output wire y1612,
  output wire y1613,
  output wire y1614,
  output wire y1615,
  output wire y1616,
  output wire y1617,
  output wire y1618,
  output wire y1619,
  output wire y1620,
  output wire y1621,
  output wire y1622,
  output wire y1623,
  output wire y1624,
  output wire y1625,
  output wire y1626,
  output wire y1627,
  output wire y1628,
  output wire y1629,
  output wire y1630,
  output wire y1631,
  output wire y1632,
  output wire y1633,
  output wire y1634,
  output wire y1635,
  output wire y1636,
  output wire y1637,
  output wire y1638,
  output wire y1639,
  output wire y1640,
  output wire y1641,
  output wire y1642,
  output wire y1643,
  output wire y1644,
  output wire y1645,
  output wire y1646,
  output wire y1647,
  output wire y1648,
  output wire y1649,
  output wire y1650,
  output wire y1651,
  output wire y1652,
  output wire y1653,
  output wire y1654,
  output wire y1655,
  output wire y1656,
  output wire y1657,
  output wire y1658,
  output wire y1659,
  output wire y1660,
  output wire y1661,
  output wire y1662,
  output wire y1663,
  output wire y1664,
  output wire y1665,
  output wire y1666,
  output wire y1667,
  output wire y1668,
  output wire y1669,
  output wire y1670,
  output wire y1671,
  output wire y1672,
  output wire y1673,
  output wire y1674,
  output wire y1675,
  output wire y1676,
  output wire y1677,
  output wire y1678,
  output wire y1679,
  output wire y1680,
  output wire y1681,
  output wire y1682,
  output wire y1683,
  output wire y1684,
  output wire y1685,
  output wire y1686,
  output wire y1687,
  output wire y1688,
  output wire y1689,
  output wire y1690,
  output wire y1691,
  output wire y1692,
  output wire y1693,
  output wire y1694,
  output wire y1695,
  output wire y1696,
  output wire y1697,
  output wire y1698,
  output wire y1699,
  output wire y1700,
  output wire y1701,
  output wire y1702,
  output wire y1703,
  output wire y1704,
  output wire y1705,
  output wire y1706,
  output wire y1707,
  output wire y1708,
  output wire y1709,
  output wire y1710,
  output wire y1711,
  output wire y1712,
  output wire y1713,
  output wire y1714,
  output wire y1715,
  output wire y1716,
  output wire y1717,
  output wire y1718,
  output wire y1719,
  output wire y1720,
  output wire y1721,
  output wire y1722,
  output wire y1723,
  output wire y1724,
  output wire y1725,
  output wire y1726,
  output wire y1727,
  output wire y1728,
  output wire y1729,
  output wire y1730,
  output wire y1731,
  output wire y1732,
  output wire y1733,
  output wire y1734,
  output wire y1735,
  output wire y1736,
  output wire y1737,
  output wire y1738,
  output wire y1739,
  output wire y1740,
  output wire y1741,
  output wire y1742,
  output wire y1743,
  output wire y1744,
  output wire y1745,
  output wire y1746,
  output wire y1747,
  output wire y1748,
  output wire y1749,
  output wire y1750,
  output wire y1751,
  output wire y1752,
  output wire y1753,
  output wire y1754,
  output wire y1755,
  output wire y1756,
  output wire y1757,
  output wire y1758,
  output wire y1759,
  output wire y1760,
  output wire y1761,
  output wire y1762,
  output wire y1763,
  output wire y1764,
  output wire y1765,
  output wire y1766,
  output wire y1767,
  output wire y1768,
  output wire y1769,
  output wire y1770,
  output wire y1771,
  output wire y1772,
  output wire y1773,
  output wire y1774,
  output wire y1775,
  output wire y1776,
  output wire y1777,
  output wire y1778,
  output wire y1779,
  output wire y1780,
  output wire y1781,
  output wire y1782,
  output wire y1783,
  output wire y1784,
  output wire y1785,
  output wire y1786,
  output wire y1787,
  output wire y1788,
  output wire y1789,
  output wire y1790,
  output wire y1791,
  output wire y1792,
  output wire y1793,
  output wire y1794,
  output wire y1795,
  output wire y1796,
  output wire y1797,
  output wire y1798,
  output wire y1799,
  output wire y1800,
  output wire y1801,
  output wire y1802,
  output wire y1803,
  output wire y1804,
  output wire y1805,
  output wire y1806,
  output wire y1807,
  output wire y1808,
  output wire y1809,
  output wire y1810,
  output wire y1811,
  output wire y1812,
  output wire y1813,
  output wire y1814,
  output wire y1815,
  output wire y1816,
  output wire y1817,
  output wire y1818,
  output wire y1819,
  output wire y1820,
  output wire y1821,
  output wire y1822,
  output wire y1823,
  output wire y1824,
  output wire y1825,
  output wire y1826,
  output wire y1827,
  output wire y1828,
  output wire y1829,
  output wire y1830,
  output wire y1831,
  output wire y1832,
  output wire y1833,
  output wire y1834,
  output wire y1835,
  output wire y1836,
  output wire y1837,
  output wire y1838,
  output wire y1839,
  output wire y1840,
  output wire y1841,
  output wire y1842,
  output wire y1843,
  output wire y1844,
  output wire y1845,
  output wire y1846,
  output wire y1847,
  output wire y1848,
  output wire y1849,
  output wire y1850,
  output wire y1851,
  output wire y1852,
  output wire y1853,
  output wire y1854,
  output wire y1855,
  output wire y1856,
  output wire y1857,
  output wire y1858,
  output wire y1859,
  output wire y1860,
  output wire y1861,
  output wire y1862,
  output wire y1863,
  output wire y1864,
  output wire y1865,
  output wire y1866,
  output wire y1867,
  output wire y1868,
  output wire y1869,
  output wire y1870,
  output wire y1871,
  output wire y1872,
  output wire y1873,
  output wire y1874,
  output wire y1875,
  output wire y1876,
  output wire y1877,
  output wire y1878,
  output wire y1879,
  output wire y1880,
  output wire y1881,
  output wire y1882,
  output wire y1883,
  output wire y1884,
  output wire y1885,
  output wire y1886,
  output wire y1887,
  output wire y1888,
  output wire y1889,
  output wire y1890,
  output wire y1891,
  output wire y1892,
  output wire y1893,
  output wire y1894,
  output wire y1895,
  output wire y1896,
  output wire y1897,
  output wire y1898,
  output wire y1899,
  output wire y1900,
  output wire y1901,
  output wire y1902,
  output wire y1903,
  output wire y1904,
  output wire y1905,
  output wire y1906,
  output wire y1907,
  output wire y1908,
  output wire y1909,
  output wire y1910,
  output wire y1911,
  output wire y1912,
  output wire y1913,
  output wire y1914,
  output wire y1915,
  output wire y1916,
  output wire y1917,
  output wire y1918,
  output wire y1919,
  output wire y1920,
  output wire y1921,
  output wire y1922,
  output wire y1923,
  output wire y1924,
  output wire y1925,
  output wire y1926,
  output wire y1927,
  output wire y1928,
  output wire y1929,
  output wire y1930,
  output wire y1931,
  output wire y1932,
  output wire y1933,
  output wire y1934,
  output wire y1935,
  output wire y1936,
  output wire y1937,
  output wire y1938,
  output wire y1939,
  output wire y1940,
  output wire y1941,
  output wire y1942,
  output wire y1943,
  output wire y1944,
  output wire y1945,
  output wire y1946,
  output wire y1947,
  output wire y1948,
  output wire y1949,
  output wire y1950,
  output wire y1951,
  output wire y1952,
  output wire y1953,
  output wire y1954,
  output wire y1955,
  output wire y1956,
  output wire y1957,
  output wire y1958,
  output wire y1959,
  output wire y1960,
  output wire y1961,
  output wire y1962,
  output wire y1963,
  output wire y1964,
  output wire y1965,
  output wire y1966,
  output wire y1967,
  output wire y1968,
  output wire y1969,
  output wire y1970,
  output wire y1971,
  output wire y1972,
  output wire y1973,
  output wire y1974,
  output wire y1975,
  output wire y1976,
  output wire y1977,
  output wire y1978,
  output wire y1979,
  output wire y1980,
  output wire y1981,
  output wire y1982,
  output wire y1983,
  output wire y1984,
  output wire y1985,
  output wire y1986,
  output wire y1987,
  output wire y1988,
  output wire y1989,
  output wire y1990,
  output wire y1991,
  output wire y1992,
  output wire y1993,
  output wire y1994,
  output wire y1995,
  output wire y1996,
  output wire y1997,
  output wire y1998,
  output wire y1999,
  output wire y2000,
  output wire y2001,
  output wire y2002,
  output wire y2003,
  output wire y2004,
  output wire y2005,
  output wire y2006,
  output wire y2007,
  output wire y2008,
  output wire y2009,
  output wire y2010,
  output wire y2011,
  output wire y2012,
  output wire y2013,
  output wire y2014,
  output wire y2015,
  output wire y2016,
  output wire y2017,
  output wire y2018,
  output wire y2019,
  output wire y2020,
  output wire y2021,
  output wire y2022,
  output wire y2023,
  output wire y2024,
  output wire y2025,
  output wire y2026,
  output wire y2027,
  output wire y2028,
  output wire y2029,
  output wire y2030,
  output wire y2031,
  output wire y2032,
  output wire y2033,
  output wire y2034,
  output wire y2035,
  output wire y2036,
  output wire y2037,
  output wire y2038,
  output wire y2039,
  output wire y2040,
  output wire y2041,
  output wire y2042,
  output wire y2043,
  output wire y2044,
  output wire y2045,
  output wire y2046,
  output wire y2047
);
  wire add_sel, sub_sel, and_sel, or_sel;
  assign add_sel = ~op1 & ~op0;
  assign sub_sel = ~op1 & op0;
  assign and_sel = op1 & ~op0;
  assign or_sel  = op1 & op0;
  wire c0;
  wire c1;
  wire c2;
  wire c3;
  wire c4;
  wire c5;
  wire c6;
  wire c7;
  wire c8;
  wire c9;
  wire c10;
  wire c11;
  wire c12;
  wire c13;
  wire c14;
  wire c15;
  wire c16;
  wire c17;
  wire c18;
  wire c19;
  wire c20;
  wire c21;
  wire c22;
  wire c23;
  wire c24;
  wire c25;
  wire c26;
  wire c27;
  wire c28;
  wire c29;
  wire c30;
  wire c31;
  wire c32;
  wire c33;
  wire c34;
  wire c35;
  wire c36;
  wire c37;
  wire c38;
  wire c39;
  wire c40;
  wire c41;
  wire c42;
  wire c43;
  wire c44;
  wire c45;
  wire c46;
  wire c47;
  wire c48;
  wire c49;
  wire c50;
  wire c51;
  wire c52;
  wire c53;
  wire c54;
  wire c55;
  wire c56;
  wire c57;
  wire c58;
  wire c59;
  wire c60;
  wire c61;
  wire c62;
  wire c63;
  wire c64;
  wire c65;
  wire c66;
  wire c67;
  wire c68;
  wire c69;
  wire c70;
  wire c71;
  wire c72;
  wire c73;
  wire c74;
  wire c75;
  wire c76;
  wire c77;
  wire c78;
  wire c79;
  wire c80;
  wire c81;
  wire c82;
  wire c83;
  wire c84;
  wire c85;
  wire c86;
  wire c87;
  wire c88;
  wire c89;
  wire c90;
  wire c91;
  wire c92;
  wire c93;
  wire c94;
  wire c95;
  wire c96;
  wire c97;
  wire c98;
  wire c99;
  wire c100;
  wire c101;
  wire c102;
  wire c103;
  wire c104;
  wire c105;
  wire c106;
  wire c107;
  wire c108;
  wire c109;
  wire c110;
  wire c111;
  wire c112;
  wire c113;
  wire c114;
  wire c115;
  wire c116;
  wire c117;
  wire c118;
  wire c119;
  wire c120;
  wire c121;
  wire c122;
  wire c123;
  wire c124;
  wire c125;
  wire c126;
  wire c127;
  wire c128;
  wire c129;
  wire c130;
  wire c131;
  wire c132;
  wire c133;
  wire c134;
  wire c135;
  wire c136;
  wire c137;
  wire c138;
  wire c139;
  wire c140;
  wire c141;
  wire c142;
  wire c143;
  wire c144;
  wire c145;
  wire c146;
  wire c147;
  wire c148;
  wire c149;
  wire c150;
  wire c151;
  wire c152;
  wire c153;
  wire c154;
  wire c155;
  wire c156;
  wire c157;
  wire c158;
  wire c159;
  wire c160;
  wire c161;
  wire c162;
  wire c163;
  wire c164;
  wire c165;
  wire c166;
  wire c167;
  wire c168;
  wire c169;
  wire c170;
  wire c171;
  wire c172;
  wire c173;
  wire c174;
  wire c175;
  wire c176;
  wire c177;
  wire c178;
  wire c179;
  wire c180;
  wire c181;
  wire c182;
  wire c183;
  wire c184;
  wire c185;
  wire c186;
  wire c187;
  wire c188;
  wire c189;
  wire c190;
  wire c191;
  wire c192;
  wire c193;
  wire c194;
  wire c195;
  wire c196;
  wire c197;
  wire c198;
  wire c199;
  wire c200;
  wire c201;
  wire c202;
  wire c203;
  wire c204;
  wire c205;
  wire c206;
  wire c207;
  wire c208;
  wire c209;
  wire c210;
  wire c211;
  wire c212;
  wire c213;
  wire c214;
  wire c215;
  wire c216;
  wire c217;
  wire c218;
  wire c219;
  wire c220;
  wire c221;
  wire c222;
  wire c223;
  wire c224;
  wire c225;
  wire c226;
  wire c227;
  wire c228;
  wire c229;
  wire c230;
  wire c231;
  wire c232;
  wire c233;
  wire c234;
  wire c235;
  wire c236;
  wire c237;
  wire c238;
  wire c239;
  wire c240;
  wire c241;
  wire c242;
  wire c243;
  wire c244;
  wire c245;
  wire c246;
  wire c247;
  wire c248;
  wire c249;
  wire c250;
  wire c251;
  wire c252;
  wire c253;
  wire c254;
  wire c255;
  wire c256;
  wire c257;
  wire c258;
  wire c259;
  wire c260;
  wire c261;
  wire c262;
  wire c263;
  wire c264;
  wire c265;
  wire c266;
  wire c267;
  wire c268;
  wire c269;
  wire c270;
  wire c271;
  wire c272;
  wire c273;
  wire c274;
  wire c275;
  wire c276;
  wire c277;
  wire c278;
  wire c279;
  wire c280;
  wire c281;
  wire c282;
  wire c283;
  wire c284;
  wire c285;
  wire c286;
  wire c287;
  wire c288;
  wire c289;
  wire c290;
  wire c291;
  wire c292;
  wire c293;
  wire c294;
  wire c295;
  wire c296;
  wire c297;
  wire c298;
  wire c299;
  wire c300;
  wire c301;
  wire c302;
  wire c303;
  wire c304;
  wire c305;
  wire c306;
  wire c307;
  wire c308;
  wire c309;
  wire c310;
  wire c311;
  wire c312;
  wire c313;
  wire c314;
  wire c315;
  wire c316;
  wire c317;
  wire c318;
  wire c319;
  wire c320;
  wire c321;
  wire c322;
  wire c323;
  wire c324;
  wire c325;
  wire c326;
  wire c327;
  wire c328;
  wire c329;
  wire c330;
  wire c331;
  wire c332;
  wire c333;
  wire c334;
  wire c335;
  wire c336;
  wire c337;
  wire c338;
  wire c339;
  wire c340;
  wire c341;
  wire c342;
  wire c343;
  wire c344;
  wire c345;
  wire c346;
  wire c347;
  wire c348;
  wire c349;
  wire c350;
  wire c351;
  wire c352;
  wire c353;
  wire c354;
  wire c355;
  wire c356;
  wire c357;
  wire c358;
  wire c359;
  wire c360;
  wire c361;
  wire c362;
  wire c363;
  wire c364;
  wire c365;
  wire c366;
  wire c367;
  wire c368;
  wire c369;
  wire c370;
  wire c371;
  wire c372;
  wire c373;
  wire c374;
  wire c375;
  wire c376;
  wire c377;
  wire c378;
  wire c379;
  wire c380;
  wire c381;
  wire c382;
  wire c383;
  wire c384;
  wire c385;
  wire c386;
  wire c387;
  wire c388;
  wire c389;
  wire c390;
  wire c391;
  wire c392;
  wire c393;
  wire c394;
  wire c395;
  wire c396;
  wire c397;
  wire c398;
  wire c399;
  wire c400;
  wire c401;
  wire c402;
  wire c403;
  wire c404;
  wire c405;
  wire c406;
  wire c407;
  wire c408;
  wire c409;
  wire c410;
  wire c411;
  wire c412;
  wire c413;
  wire c414;
  wire c415;
  wire c416;
  wire c417;
  wire c418;
  wire c419;
  wire c420;
  wire c421;
  wire c422;
  wire c423;
  wire c424;
  wire c425;
  wire c426;
  wire c427;
  wire c428;
  wire c429;
  wire c430;
  wire c431;
  wire c432;
  wire c433;
  wire c434;
  wire c435;
  wire c436;
  wire c437;
  wire c438;
  wire c439;
  wire c440;
  wire c441;
  wire c442;
  wire c443;
  wire c444;
  wire c445;
  wire c446;
  wire c447;
  wire c448;
  wire c449;
  wire c450;
  wire c451;
  wire c452;
  wire c453;
  wire c454;
  wire c455;
  wire c456;
  wire c457;
  wire c458;
  wire c459;
  wire c460;
  wire c461;
  wire c462;
  wire c463;
  wire c464;
  wire c465;
  wire c466;
  wire c467;
  wire c468;
  wire c469;
  wire c470;
  wire c471;
  wire c472;
  wire c473;
  wire c474;
  wire c475;
  wire c476;
  wire c477;
  wire c478;
  wire c479;
  wire c480;
  wire c481;
  wire c482;
  wire c483;
  wire c484;
  wire c485;
  wire c486;
  wire c487;
  wire c488;
  wire c489;
  wire c490;
  wire c491;
  wire c492;
  wire c493;
  wire c494;
  wire c495;
  wire c496;
  wire c497;
  wire c498;
  wire c499;
  wire c500;
  wire c501;
  wire c502;
  wire c503;
  wire c504;
  wire c505;
  wire c506;
  wire c507;
  wire c508;
  wire c509;
  wire c510;
  wire c511;
  wire c512;
  wire c513;
  wire c514;
  wire c515;
  wire c516;
  wire c517;
  wire c518;
  wire c519;
  wire c520;
  wire c521;
  wire c522;
  wire c523;
  wire c524;
  wire c525;
  wire c526;
  wire c527;
  wire c528;
  wire c529;
  wire c530;
  wire c531;
  wire c532;
  wire c533;
  wire c534;
  wire c535;
  wire c536;
  wire c537;
  wire c538;
  wire c539;
  wire c540;
  wire c541;
  wire c542;
  wire c543;
  wire c544;
  wire c545;
  wire c546;
  wire c547;
  wire c548;
  wire c549;
  wire c550;
  wire c551;
  wire c552;
  wire c553;
  wire c554;
  wire c555;
  wire c556;
  wire c557;
  wire c558;
  wire c559;
  wire c560;
  wire c561;
  wire c562;
  wire c563;
  wire c564;
  wire c565;
  wire c566;
  wire c567;
  wire c568;
  wire c569;
  wire c570;
  wire c571;
  wire c572;
  wire c573;
  wire c574;
  wire c575;
  wire c576;
  wire c577;
  wire c578;
  wire c579;
  wire c580;
  wire c581;
  wire c582;
  wire c583;
  wire c584;
  wire c585;
  wire c586;
  wire c587;
  wire c588;
  wire c589;
  wire c590;
  wire c591;
  wire c592;
  wire c593;
  wire c594;
  wire c595;
  wire c596;
  wire c597;
  wire c598;
  wire c599;
  wire c600;
  wire c601;
  wire c602;
  wire c603;
  wire c604;
  wire c605;
  wire c606;
  wire c607;
  wire c608;
  wire c609;
  wire c610;
  wire c611;
  wire c612;
  wire c613;
  wire c614;
  wire c615;
  wire c616;
  wire c617;
  wire c618;
  wire c619;
  wire c620;
  wire c621;
  wire c622;
  wire c623;
  wire c624;
  wire c625;
  wire c626;
  wire c627;
  wire c628;
  wire c629;
  wire c630;
  wire c631;
  wire c632;
  wire c633;
  wire c634;
  wire c635;
  wire c636;
  wire c637;
  wire c638;
  wire c639;
  wire c640;
  wire c641;
  wire c642;
  wire c643;
  wire c644;
  wire c645;
  wire c646;
  wire c647;
  wire c648;
  wire c649;
  wire c650;
  wire c651;
  wire c652;
  wire c653;
  wire c654;
  wire c655;
  wire c656;
  wire c657;
  wire c658;
  wire c659;
  wire c660;
  wire c661;
  wire c662;
  wire c663;
  wire c664;
  wire c665;
  wire c666;
  wire c667;
  wire c668;
  wire c669;
  wire c670;
  wire c671;
  wire c672;
  wire c673;
  wire c674;
  wire c675;
  wire c676;
  wire c677;
  wire c678;
  wire c679;
  wire c680;
  wire c681;
  wire c682;
  wire c683;
  wire c684;
  wire c685;
  wire c686;
  wire c687;
  wire c688;
  wire c689;
  wire c690;
  wire c691;
  wire c692;
  wire c693;
  wire c694;
  wire c695;
  wire c696;
  wire c697;
  wire c698;
  wire c699;
  wire c700;
  wire c701;
  wire c702;
  wire c703;
  wire c704;
  wire c705;
  wire c706;
  wire c707;
  wire c708;
  wire c709;
  wire c710;
  wire c711;
  wire c712;
  wire c713;
  wire c714;
  wire c715;
  wire c716;
  wire c717;
  wire c718;
  wire c719;
  wire c720;
  wire c721;
  wire c722;
  wire c723;
  wire c724;
  wire c725;
  wire c726;
  wire c727;
  wire c728;
  wire c729;
  wire c730;
  wire c731;
  wire c732;
  wire c733;
  wire c734;
  wire c735;
  wire c736;
  wire c737;
  wire c738;
  wire c739;
  wire c740;
  wire c741;
  wire c742;
  wire c743;
  wire c744;
  wire c745;
  wire c746;
  wire c747;
  wire c748;
  wire c749;
  wire c750;
  wire c751;
  wire c752;
  wire c753;
  wire c754;
  wire c755;
  wire c756;
  wire c757;
  wire c758;
  wire c759;
  wire c760;
  wire c761;
  wire c762;
  wire c763;
  wire c764;
  wire c765;
  wire c766;
  wire c767;
  wire c768;
  wire c769;
  wire c770;
  wire c771;
  wire c772;
  wire c773;
  wire c774;
  wire c775;
  wire c776;
  wire c777;
  wire c778;
  wire c779;
  wire c780;
  wire c781;
  wire c782;
  wire c783;
  wire c784;
  wire c785;
  wire c786;
  wire c787;
  wire c788;
  wire c789;
  wire c790;
  wire c791;
  wire c792;
  wire c793;
  wire c794;
  wire c795;
  wire c796;
  wire c797;
  wire c798;
  wire c799;
  wire c800;
  wire c801;
  wire c802;
  wire c803;
  wire c804;
  wire c805;
  wire c806;
  wire c807;
  wire c808;
  wire c809;
  wire c810;
  wire c811;
  wire c812;
  wire c813;
  wire c814;
  wire c815;
  wire c816;
  wire c817;
  wire c818;
  wire c819;
  wire c820;
  wire c821;
  wire c822;
  wire c823;
  wire c824;
  wire c825;
  wire c826;
  wire c827;
  wire c828;
  wire c829;
  wire c830;
  wire c831;
  wire c832;
  wire c833;
  wire c834;
  wire c835;
  wire c836;
  wire c837;
  wire c838;
  wire c839;
  wire c840;
  wire c841;
  wire c842;
  wire c843;
  wire c844;
  wire c845;
  wire c846;
  wire c847;
  wire c848;
  wire c849;
  wire c850;
  wire c851;
  wire c852;
  wire c853;
  wire c854;
  wire c855;
  wire c856;
  wire c857;
  wire c858;
  wire c859;
  wire c860;
  wire c861;
  wire c862;
  wire c863;
  wire c864;
  wire c865;
  wire c866;
  wire c867;
  wire c868;
  wire c869;
  wire c870;
  wire c871;
  wire c872;
  wire c873;
  wire c874;
  wire c875;
  wire c876;
  wire c877;
  wire c878;
  wire c879;
  wire c880;
  wire c881;
  wire c882;
  wire c883;
  wire c884;
  wire c885;
  wire c886;
  wire c887;
  wire c888;
  wire c889;
  wire c890;
  wire c891;
  wire c892;
  wire c893;
  wire c894;
  wire c895;
  wire c896;
  wire c897;
  wire c898;
  wire c899;
  wire c900;
  wire c901;
  wire c902;
  wire c903;
  wire c904;
  wire c905;
  wire c906;
  wire c907;
  wire c908;
  wire c909;
  wire c910;
  wire c911;
  wire c912;
  wire c913;
  wire c914;
  wire c915;
  wire c916;
  wire c917;
  wire c918;
  wire c919;
  wire c920;
  wire c921;
  wire c922;
  wire c923;
  wire c924;
  wire c925;
  wire c926;
  wire c927;
  wire c928;
  wire c929;
  wire c930;
  wire c931;
  wire c932;
  wire c933;
  wire c934;
  wire c935;
  wire c936;
  wire c937;
  wire c938;
  wire c939;
  wire c940;
  wire c941;
  wire c942;
  wire c943;
  wire c944;
  wire c945;
  wire c946;
  wire c947;
  wire c948;
  wire c949;
  wire c950;
  wire c951;
  wire c952;
  wire c953;
  wire c954;
  wire c955;
  wire c956;
  wire c957;
  wire c958;
  wire c959;
  wire c960;
  wire c961;
  wire c962;
  wire c963;
  wire c964;
  wire c965;
  wire c966;
  wire c967;
  wire c968;
  wire c969;
  wire c970;
  wire c971;
  wire c972;
  wire c973;
  wire c974;
  wire c975;
  wire c976;
  wire c977;
  wire c978;
  wire c979;
  wire c980;
  wire c981;
  wire c982;
  wire c983;
  wire c984;
  wire c985;
  wire c986;
  wire c987;
  wire c988;
  wire c989;
  wire c990;
  wire c991;
  wire c992;
  wire c993;
  wire c994;
  wire c995;
  wire c996;
  wire c997;
  wire c998;
  wire c999;
  wire c1000;
  wire c1001;
  wire c1002;
  wire c1003;
  wire c1004;
  wire c1005;
  wire c1006;
  wire c1007;
  wire c1008;
  wire c1009;
  wire c1010;
  wire c1011;
  wire c1012;
  wire c1013;
  wire c1014;
  wire c1015;
  wire c1016;
  wire c1017;
  wire c1018;
  wire c1019;
  wire c1020;
  wire c1021;
  wire c1022;
  wire c1023;
  wire c1024;
  wire c1025;
  wire c1026;
  wire c1027;
  wire c1028;
  wire c1029;
  wire c1030;
  wire c1031;
  wire c1032;
  wire c1033;
  wire c1034;
  wire c1035;
  wire c1036;
  wire c1037;
  wire c1038;
  wire c1039;
  wire c1040;
  wire c1041;
  wire c1042;
  wire c1043;
  wire c1044;
  wire c1045;
  wire c1046;
  wire c1047;
  wire c1048;
  wire c1049;
  wire c1050;
  wire c1051;
  wire c1052;
  wire c1053;
  wire c1054;
  wire c1055;
  wire c1056;
  wire c1057;
  wire c1058;
  wire c1059;
  wire c1060;
  wire c1061;
  wire c1062;
  wire c1063;
  wire c1064;
  wire c1065;
  wire c1066;
  wire c1067;
  wire c1068;
  wire c1069;
  wire c1070;
  wire c1071;
  wire c1072;
  wire c1073;
  wire c1074;
  wire c1075;
  wire c1076;
  wire c1077;
  wire c1078;
  wire c1079;
  wire c1080;
  wire c1081;
  wire c1082;
  wire c1083;
  wire c1084;
  wire c1085;
  wire c1086;
  wire c1087;
  wire c1088;
  wire c1089;
  wire c1090;
  wire c1091;
  wire c1092;
  wire c1093;
  wire c1094;
  wire c1095;
  wire c1096;
  wire c1097;
  wire c1098;
  wire c1099;
  wire c1100;
  wire c1101;
  wire c1102;
  wire c1103;
  wire c1104;
  wire c1105;
  wire c1106;
  wire c1107;
  wire c1108;
  wire c1109;
  wire c1110;
  wire c1111;
  wire c1112;
  wire c1113;
  wire c1114;
  wire c1115;
  wire c1116;
  wire c1117;
  wire c1118;
  wire c1119;
  wire c1120;
  wire c1121;
  wire c1122;
  wire c1123;
  wire c1124;
  wire c1125;
  wire c1126;
  wire c1127;
  wire c1128;
  wire c1129;
  wire c1130;
  wire c1131;
  wire c1132;
  wire c1133;
  wire c1134;
  wire c1135;
  wire c1136;
  wire c1137;
  wire c1138;
  wire c1139;
  wire c1140;
  wire c1141;
  wire c1142;
  wire c1143;
  wire c1144;
  wire c1145;
  wire c1146;
  wire c1147;
  wire c1148;
  wire c1149;
  wire c1150;
  wire c1151;
  wire c1152;
  wire c1153;
  wire c1154;
  wire c1155;
  wire c1156;
  wire c1157;
  wire c1158;
  wire c1159;
  wire c1160;
  wire c1161;
  wire c1162;
  wire c1163;
  wire c1164;
  wire c1165;
  wire c1166;
  wire c1167;
  wire c1168;
  wire c1169;
  wire c1170;
  wire c1171;
  wire c1172;
  wire c1173;
  wire c1174;
  wire c1175;
  wire c1176;
  wire c1177;
  wire c1178;
  wire c1179;
  wire c1180;
  wire c1181;
  wire c1182;
  wire c1183;
  wire c1184;
  wire c1185;
  wire c1186;
  wire c1187;
  wire c1188;
  wire c1189;
  wire c1190;
  wire c1191;
  wire c1192;
  wire c1193;
  wire c1194;
  wire c1195;
  wire c1196;
  wire c1197;
  wire c1198;
  wire c1199;
  wire c1200;
  wire c1201;
  wire c1202;
  wire c1203;
  wire c1204;
  wire c1205;
  wire c1206;
  wire c1207;
  wire c1208;
  wire c1209;
  wire c1210;
  wire c1211;
  wire c1212;
  wire c1213;
  wire c1214;
  wire c1215;
  wire c1216;
  wire c1217;
  wire c1218;
  wire c1219;
  wire c1220;
  wire c1221;
  wire c1222;
  wire c1223;
  wire c1224;
  wire c1225;
  wire c1226;
  wire c1227;
  wire c1228;
  wire c1229;
  wire c1230;
  wire c1231;
  wire c1232;
  wire c1233;
  wire c1234;
  wire c1235;
  wire c1236;
  wire c1237;
  wire c1238;
  wire c1239;
  wire c1240;
  wire c1241;
  wire c1242;
  wire c1243;
  wire c1244;
  wire c1245;
  wire c1246;
  wire c1247;
  wire c1248;
  wire c1249;
  wire c1250;
  wire c1251;
  wire c1252;
  wire c1253;
  wire c1254;
  wire c1255;
  wire c1256;
  wire c1257;
  wire c1258;
  wire c1259;
  wire c1260;
  wire c1261;
  wire c1262;
  wire c1263;
  wire c1264;
  wire c1265;
  wire c1266;
  wire c1267;
  wire c1268;
  wire c1269;
  wire c1270;
  wire c1271;
  wire c1272;
  wire c1273;
  wire c1274;
  wire c1275;
  wire c1276;
  wire c1277;
  wire c1278;
  wire c1279;
  wire c1280;
  wire c1281;
  wire c1282;
  wire c1283;
  wire c1284;
  wire c1285;
  wire c1286;
  wire c1287;
  wire c1288;
  wire c1289;
  wire c1290;
  wire c1291;
  wire c1292;
  wire c1293;
  wire c1294;
  wire c1295;
  wire c1296;
  wire c1297;
  wire c1298;
  wire c1299;
  wire c1300;
  wire c1301;
  wire c1302;
  wire c1303;
  wire c1304;
  wire c1305;
  wire c1306;
  wire c1307;
  wire c1308;
  wire c1309;
  wire c1310;
  wire c1311;
  wire c1312;
  wire c1313;
  wire c1314;
  wire c1315;
  wire c1316;
  wire c1317;
  wire c1318;
  wire c1319;
  wire c1320;
  wire c1321;
  wire c1322;
  wire c1323;
  wire c1324;
  wire c1325;
  wire c1326;
  wire c1327;
  wire c1328;
  wire c1329;
  wire c1330;
  wire c1331;
  wire c1332;
  wire c1333;
  wire c1334;
  wire c1335;
  wire c1336;
  wire c1337;
  wire c1338;
  wire c1339;
  wire c1340;
  wire c1341;
  wire c1342;
  wire c1343;
  wire c1344;
  wire c1345;
  wire c1346;
  wire c1347;
  wire c1348;
  wire c1349;
  wire c1350;
  wire c1351;
  wire c1352;
  wire c1353;
  wire c1354;
  wire c1355;
  wire c1356;
  wire c1357;
  wire c1358;
  wire c1359;
  wire c1360;
  wire c1361;
  wire c1362;
  wire c1363;
  wire c1364;
  wire c1365;
  wire c1366;
  wire c1367;
  wire c1368;
  wire c1369;
  wire c1370;
  wire c1371;
  wire c1372;
  wire c1373;
  wire c1374;
  wire c1375;
  wire c1376;
  wire c1377;
  wire c1378;
  wire c1379;
  wire c1380;
  wire c1381;
  wire c1382;
  wire c1383;
  wire c1384;
  wire c1385;
  wire c1386;
  wire c1387;
  wire c1388;
  wire c1389;
  wire c1390;
  wire c1391;
  wire c1392;
  wire c1393;
  wire c1394;
  wire c1395;
  wire c1396;
  wire c1397;
  wire c1398;
  wire c1399;
  wire c1400;
  wire c1401;
  wire c1402;
  wire c1403;
  wire c1404;
  wire c1405;
  wire c1406;
  wire c1407;
  wire c1408;
  wire c1409;
  wire c1410;
  wire c1411;
  wire c1412;
  wire c1413;
  wire c1414;
  wire c1415;
  wire c1416;
  wire c1417;
  wire c1418;
  wire c1419;
  wire c1420;
  wire c1421;
  wire c1422;
  wire c1423;
  wire c1424;
  wire c1425;
  wire c1426;
  wire c1427;
  wire c1428;
  wire c1429;
  wire c1430;
  wire c1431;
  wire c1432;
  wire c1433;
  wire c1434;
  wire c1435;
  wire c1436;
  wire c1437;
  wire c1438;
  wire c1439;
  wire c1440;
  wire c1441;
  wire c1442;
  wire c1443;
  wire c1444;
  wire c1445;
  wire c1446;
  wire c1447;
  wire c1448;
  wire c1449;
  wire c1450;
  wire c1451;
  wire c1452;
  wire c1453;
  wire c1454;
  wire c1455;
  wire c1456;
  wire c1457;
  wire c1458;
  wire c1459;
  wire c1460;
  wire c1461;
  wire c1462;
  wire c1463;
  wire c1464;
  wire c1465;
  wire c1466;
  wire c1467;
  wire c1468;
  wire c1469;
  wire c1470;
  wire c1471;
  wire c1472;
  wire c1473;
  wire c1474;
  wire c1475;
  wire c1476;
  wire c1477;
  wire c1478;
  wire c1479;
  wire c1480;
  wire c1481;
  wire c1482;
  wire c1483;
  wire c1484;
  wire c1485;
  wire c1486;
  wire c1487;
  wire c1488;
  wire c1489;
  wire c1490;
  wire c1491;
  wire c1492;
  wire c1493;
  wire c1494;
  wire c1495;
  wire c1496;
  wire c1497;
  wire c1498;
  wire c1499;
  wire c1500;
  wire c1501;
  wire c1502;
  wire c1503;
  wire c1504;
  wire c1505;
  wire c1506;
  wire c1507;
  wire c1508;
  wire c1509;
  wire c1510;
  wire c1511;
  wire c1512;
  wire c1513;
  wire c1514;
  wire c1515;
  wire c1516;
  wire c1517;
  wire c1518;
  wire c1519;
  wire c1520;
  wire c1521;
  wire c1522;
  wire c1523;
  wire c1524;
  wire c1525;
  wire c1526;
  wire c1527;
  wire c1528;
  wire c1529;
  wire c1530;
  wire c1531;
  wire c1532;
  wire c1533;
  wire c1534;
  wire c1535;
  wire c1536;
  wire c1537;
  wire c1538;
  wire c1539;
  wire c1540;
  wire c1541;
  wire c1542;
  wire c1543;
  wire c1544;
  wire c1545;
  wire c1546;
  wire c1547;
  wire c1548;
  wire c1549;
  wire c1550;
  wire c1551;
  wire c1552;
  wire c1553;
  wire c1554;
  wire c1555;
  wire c1556;
  wire c1557;
  wire c1558;
  wire c1559;
  wire c1560;
  wire c1561;
  wire c1562;
  wire c1563;
  wire c1564;
  wire c1565;
  wire c1566;
  wire c1567;
  wire c1568;
  wire c1569;
  wire c1570;
  wire c1571;
  wire c1572;
  wire c1573;
  wire c1574;
  wire c1575;
  wire c1576;
  wire c1577;
  wire c1578;
  wire c1579;
  wire c1580;
  wire c1581;
  wire c1582;
  wire c1583;
  wire c1584;
  wire c1585;
  wire c1586;
  wire c1587;
  wire c1588;
  wire c1589;
  wire c1590;
  wire c1591;
  wire c1592;
  wire c1593;
  wire c1594;
  wire c1595;
  wire c1596;
  wire c1597;
  wire c1598;
  wire c1599;
  wire c1600;
  wire c1601;
  wire c1602;
  wire c1603;
  wire c1604;
  wire c1605;
  wire c1606;
  wire c1607;
  wire c1608;
  wire c1609;
  wire c1610;
  wire c1611;
  wire c1612;
  wire c1613;
  wire c1614;
  wire c1615;
  wire c1616;
  wire c1617;
  wire c1618;
  wire c1619;
  wire c1620;
  wire c1621;
  wire c1622;
  wire c1623;
  wire c1624;
  wire c1625;
  wire c1626;
  wire c1627;
  wire c1628;
  wire c1629;
  wire c1630;
  wire c1631;
  wire c1632;
  wire c1633;
  wire c1634;
  wire c1635;
  wire c1636;
  wire c1637;
  wire c1638;
  wire c1639;
  wire c1640;
  wire c1641;
  wire c1642;
  wire c1643;
  wire c1644;
  wire c1645;
  wire c1646;
  wire c1647;
  wire c1648;
  wire c1649;
  wire c1650;
  wire c1651;
  wire c1652;
  wire c1653;
  wire c1654;
  wire c1655;
  wire c1656;
  wire c1657;
  wire c1658;
  wire c1659;
  wire c1660;
  wire c1661;
  wire c1662;
  wire c1663;
  wire c1664;
  wire c1665;
  wire c1666;
  wire c1667;
  wire c1668;
  wire c1669;
  wire c1670;
  wire c1671;
  wire c1672;
  wire c1673;
  wire c1674;
  wire c1675;
  wire c1676;
  wire c1677;
  wire c1678;
  wire c1679;
  wire c1680;
  wire c1681;
  wire c1682;
  wire c1683;
  wire c1684;
  wire c1685;
  wire c1686;
  wire c1687;
  wire c1688;
  wire c1689;
  wire c1690;
  wire c1691;
  wire c1692;
  wire c1693;
  wire c1694;
  wire c1695;
  wire c1696;
  wire c1697;
  wire c1698;
  wire c1699;
  wire c1700;
  wire c1701;
  wire c1702;
  wire c1703;
  wire c1704;
  wire c1705;
  wire c1706;
  wire c1707;
  wire c1708;
  wire c1709;
  wire c1710;
  wire c1711;
  wire c1712;
  wire c1713;
  wire c1714;
  wire c1715;
  wire c1716;
  wire c1717;
  wire c1718;
  wire c1719;
  wire c1720;
  wire c1721;
  wire c1722;
  wire c1723;
  wire c1724;
  wire c1725;
  wire c1726;
  wire c1727;
  wire c1728;
  wire c1729;
  wire c1730;
  wire c1731;
  wire c1732;
  wire c1733;
  wire c1734;
  wire c1735;
  wire c1736;
  wire c1737;
  wire c1738;
  wire c1739;
  wire c1740;
  wire c1741;
  wire c1742;
  wire c1743;
  wire c1744;
  wire c1745;
  wire c1746;
  wire c1747;
  wire c1748;
  wire c1749;
  wire c1750;
  wire c1751;
  wire c1752;
  wire c1753;
  wire c1754;
  wire c1755;
  wire c1756;
  wire c1757;
  wire c1758;
  wire c1759;
  wire c1760;
  wire c1761;
  wire c1762;
  wire c1763;
  wire c1764;
  wire c1765;
  wire c1766;
  wire c1767;
  wire c1768;
  wire c1769;
  wire c1770;
  wire c1771;
  wire c1772;
  wire c1773;
  wire c1774;
  wire c1775;
  wire c1776;
  wire c1777;
  wire c1778;
  wire c1779;
  wire c1780;
  wire c1781;
  wire c1782;
  wire c1783;
  wire c1784;
  wire c1785;
  wire c1786;
  wire c1787;
  wire c1788;
  wire c1789;
  wire c1790;
  wire c1791;
  wire c1792;
  wire c1793;
  wire c1794;
  wire c1795;
  wire c1796;
  wire c1797;
  wire c1798;
  wire c1799;
  wire c1800;
  wire c1801;
  wire c1802;
  wire c1803;
  wire c1804;
  wire c1805;
  wire c1806;
  wire c1807;
  wire c1808;
  wire c1809;
  wire c1810;
  wire c1811;
  wire c1812;
  wire c1813;
  wire c1814;
  wire c1815;
  wire c1816;
  wire c1817;
  wire c1818;
  wire c1819;
  wire c1820;
  wire c1821;
  wire c1822;
  wire c1823;
  wire c1824;
  wire c1825;
  wire c1826;
  wire c1827;
  wire c1828;
  wire c1829;
  wire c1830;
  wire c1831;
  wire c1832;
  wire c1833;
  wire c1834;
  wire c1835;
  wire c1836;
  wire c1837;
  wire c1838;
  wire c1839;
  wire c1840;
  wire c1841;
  wire c1842;
  wire c1843;
  wire c1844;
  wire c1845;
  wire c1846;
  wire c1847;
  wire c1848;
  wire c1849;
  wire c1850;
  wire c1851;
  wire c1852;
  wire c1853;
  wire c1854;
  wire c1855;
  wire c1856;
  wire c1857;
  wire c1858;
  wire c1859;
  wire c1860;
  wire c1861;
  wire c1862;
  wire c1863;
  wire c1864;
  wire c1865;
  wire c1866;
  wire c1867;
  wire c1868;
  wire c1869;
  wire c1870;
  wire c1871;
  wire c1872;
  wire c1873;
  wire c1874;
  wire c1875;
  wire c1876;
  wire c1877;
  wire c1878;
  wire c1879;
  wire c1880;
  wire c1881;
  wire c1882;
  wire c1883;
  wire c1884;
  wire c1885;
  wire c1886;
  wire c1887;
  wire c1888;
  wire c1889;
  wire c1890;
  wire c1891;
  wire c1892;
  wire c1893;
  wire c1894;
  wire c1895;
  wire c1896;
  wire c1897;
  wire c1898;
  wire c1899;
  wire c1900;
  wire c1901;
  wire c1902;
  wire c1903;
  wire c1904;
  wire c1905;
  wire c1906;
  wire c1907;
  wire c1908;
  wire c1909;
  wire c1910;
  wire c1911;
  wire c1912;
  wire c1913;
  wire c1914;
  wire c1915;
  wire c1916;
  wire c1917;
  wire c1918;
  wire c1919;
  wire c1920;
  wire c1921;
  wire c1922;
  wire c1923;
  wire c1924;
  wire c1925;
  wire c1926;
  wire c1927;
  wire c1928;
  wire c1929;
  wire c1930;
  wire c1931;
  wire c1932;
  wire c1933;
  wire c1934;
  wire c1935;
  wire c1936;
  wire c1937;
  wire c1938;
  wire c1939;
  wire c1940;
  wire c1941;
  wire c1942;
  wire c1943;
  wire c1944;
  wire c1945;
  wire c1946;
  wire c1947;
  wire c1948;
  wire c1949;
  wire c1950;
  wire c1951;
  wire c1952;
  wire c1953;
  wire c1954;
  wire c1955;
  wire c1956;
  wire c1957;
  wire c1958;
  wire c1959;
  wire c1960;
  wire c1961;
  wire c1962;
  wire c1963;
  wire c1964;
  wire c1965;
  wire c1966;
  wire c1967;
  wire c1968;
  wire c1969;
  wire c1970;
  wire c1971;
  wire c1972;
  wire c1973;
  wire c1974;
  wire c1975;
  wire c1976;
  wire c1977;
  wire c1978;
  wire c1979;
  wire c1980;
  wire c1981;
  wire c1982;
  wire c1983;
  wire c1984;
  wire c1985;
  wire c1986;
  wire c1987;
  wire c1988;
  wire c1989;
  wire c1990;
  wire c1991;
  wire c1992;
  wire c1993;
  wire c1994;
  wire c1995;
  wire c1996;
  wire c1997;
  wire c1998;
  wire c1999;
  wire c2000;
  wire c2001;
  wire c2002;
  wire c2003;
  wire c2004;
  wire c2005;
  wire c2006;
  wire c2007;
  wire c2008;
  wire c2009;
  wire c2010;
  wire c2011;
  wire c2012;
  wire c2013;
  wire c2014;
  wire c2015;
  wire c2016;
  wire c2017;
  wire c2018;
  wire c2019;
  wire c2020;
  wire c2021;
  wire c2022;
  wire c2023;
  wire c2024;
  wire c2025;
  wire c2026;
  wire c2027;
  wire c2028;
  wire c2029;
  wire c2030;
  wire c2031;
  wire c2032;
  wire c2033;
  wire c2034;
  wire c2035;
  wire c2036;
  wire c2037;
  wire c2038;
  wire c2039;
  wire c2040;
  wire c2041;
  wire c2042;
  wire c2043;
  wire c2044;
  wire c2045;
  wire c2046;
  wire c2047;
  wire c2048;
  assign c0 = 1'b0;
  wire s0, sub0, and0, or0;
  wire b_inv0;
  assign b_inv0 = ~b0;
  assign s0  = a0 ^ b0 ^ c0;
  assign sub0 = a0 ^ b_inv0 ^ c0;
  assign and0 = a0 & b0;
  assign or0  = a0 | b0;
  assign c1 = (a0 & b0) | (a0 & c0) | (b0 & c0);
  wire c_sub1;
  assign c_sub1 = (a0 & b_inv0) | (a0 & c0) | (b_inv0 & c0);
  wire s1, sub1, and1, or1;
  wire b_inv1;
  assign b_inv1 = ~b1;
  assign s1  = a1 ^ b1 ^ c1;
  assign sub1 = a1 ^ b_inv1 ^ c1;
  assign and1 = a1 & b1;
  assign or1  = a1 | b1;
  assign c2 = (a1 & b1) | (a1 & c1) | (b1 & c1);
  wire c_sub2;
  assign c_sub2 = (a1 & b_inv1) | (a1 & c1) | (b_inv1 & c1);
  wire s2, sub2, and2, or2;
  wire b_inv2;
  assign b_inv2 = ~b2;
  assign s2  = a2 ^ b2 ^ c2;
  assign sub2 = a2 ^ b_inv2 ^ c2;
  assign and2 = a2 & b2;
  assign or2  = a2 | b2;
  assign c3 = (a2 & b2) | (a2 & c2) | (b2 & c2);
  wire c_sub3;
  assign c_sub3 = (a2 & b_inv2) | (a2 & c2) | (b_inv2 & c2);
  wire s3, sub3, and3, or3;
  wire b_inv3;
  assign b_inv3 = ~b3;
  assign s3  = a3 ^ b3 ^ c3;
  assign sub3 = a3 ^ b_inv3 ^ c3;
  assign and3 = a3 & b3;
  assign or3  = a3 | b3;
  assign c4 = (a3 & b3) | (a3 & c3) | (b3 & c3);
  wire c_sub4;
  assign c_sub4 = (a3 & b_inv3) | (a3 & c3) | (b_inv3 & c3);
  wire s4, sub4, and4, or4;
  wire b_inv4;
  assign b_inv4 = ~b4;
  assign s4  = a4 ^ b4 ^ c4;
  assign sub4 = a4 ^ b_inv4 ^ c4;
  assign and4 = a4 & b4;
  assign or4  = a4 | b4;
  assign c5 = (a4 & b4) | (a4 & c4) | (b4 & c4);
  wire c_sub5;
  assign c_sub5 = (a4 & b_inv4) | (a4 & c4) | (b_inv4 & c4);
  wire s5, sub5, and5, or5;
  wire b_inv5;
  assign b_inv5 = ~b5;
  assign s5  = a5 ^ b5 ^ c5;
  assign sub5 = a5 ^ b_inv5 ^ c5;
  assign and5 = a5 & b5;
  assign or5  = a5 | b5;
  assign c6 = (a5 & b5) | (a5 & c5) | (b5 & c5);
  wire c_sub6;
  assign c_sub6 = (a5 & b_inv5) | (a5 & c5) | (b_inv5 & c5);
  wire s6, sub6, and6, or6;
  wire b_inv6;
  assign b_inv6 = ~b6;
  assign s6  = a6 ^ b6 ^ c6;
  assign sub6 = a6 ^ b_inv6 ^ c6;
  assign and6 = a6 & b6;
  assign or6  = a6 | b6;
  assign c7 = (a6 & b6) | (a6 & c6) | (b6 & c6);
  wire c_sub7;
  assign c_sub7 = (a6 & b_inv6) | (a6 & c6) | (b_inv6 & c6);
  wire s7, sub7, and7, or7;
  wire b_inv7;
  assign b_inv7 = ~b7;
  assign s7  = a7 ^ b7 ^ c7;
  assign sub7 = a7 ^ b_inv7 ^ c7;
  assign and7 = a7 & b7;
  assign or7  = a7 | b7;
  assign c8 = (a7 & b7) | (a7 & c7) | (b7 & c7);
  wire c_sub8;
  assign c_sub8 = (a7 & b_inv7) | (a7 & c7) | (b_inv7 & c7);
  wire s8, sub8, and8, or8;
  wire b_inv8;
  assign b_inv8 = ~b8;
  assign s8  = a8 ^ b8 ^ c8;
  assign sub8 = a8 ^ b_inv8 ^ c8;
  assign and8 = a8 & b8;
  assign or8  = a8 | b8;
  assign c9 = (a8 & b8) | (a8 & c8) | (b8 & c8);
  wire c_sub9;
  assign c_sub9 = (a8 & b_inv8) | (a8 & c8) | (b_inv8 & c8);
  wire s9, sub9, and9, or9;
  wire b_inv9;
  assign b_inv9 = ~b9;
  assign s9  = a9 ^ b9 ^ c9;
  assign sub9 = a9 ^ b_inv9 ^ c9;
  assign and9 = a9 & b9;
  assign or9  = a9 | b9;
  assign c10 = (a9 & b9) | (a9 & c9) | (b9 & c9);
  wire c_sub10;
  assign c_sub10 = (a9 & b_inv9) | (a9 & c9) | (b_inv9 & c9);
  wire s10, sub10, and10, or10;
  wire b_inv10;
  assign b_inv10 = ~b10;
  assign s10  = a10 ^ b10 ^ c10;
  assign sub10 = a10 ^ b_inv10 ^ c10;
  assign and10 = a10 & b10;
  assign or10  = a10 | b10;
  assign c11 = (a10 & b10) | (a10 & c10) | (b10 & c10);
  wire c_sub11;
  assign c_sub11 = (a10 & b_inv10) | (a10 & c10) | (b_inv10 & c10);
  wire s11, sub11, and11, or11;
  wire b_inv11;
  assign b_inv11 = ~b11;
  assign s11  = a11 ^ b11 ^ c11;
  assign sub11 = a11 ^ b_inv11 ^ c11;
  assign and11 = a11 & b11;
  assign or11  = a11 | b11;
  assign c12 = (a11 & b11) | (a11 & c11) | (b11 & c11);
  wire c_sub12;
  assign c_sub12 = (a11 & b_inv11) | (a11 & c11) | (b_inv11 & c11);
  wire s12, sub12, and12, or12;
  wire b_inv12;
  assign b_inv12 = ~b12;
  assign s12  = a12 ^ b12 ^ c12;
  assign sub12 = a12 ^ b_inv12 ^ c12;
  assign and12 = a12 & b12;
  assign or12  = a12 | b12;
  assign c13 = (a12 & b12) | (a12 & c12) | (b12 & c12);
  wire c_sub13;
  assign c_sub13 = (a12 & b_inv12) | (a12 & c12) | (b_inv12 & c12);
  wire s13, sub13, and13, or13;
  wire b_inv13;
  assign b_inv13 = ~b13;
  assign s13  = a13 ^ b13 ^ c13;
  assign sub13 = a13 ^ b_inv13 ^ c13;
  assign and13 = a13 & b13;
  assign or13  = a13 | b13;
  assign c14 = (a13 & b13) | (a13 & c13) | (b13 & c13);
  wire c_sub14;
  assign c_sub14 = (a13 & b_inv13) | (a13 & c13) | (b_inv13 & c13);
  wire s14, sub14, and14, or14;
  wire b_inv14;
  assign b_inv14 = ~b14;
  assign s14  = a14 ^ b14 ^ c14;
  assign sub14 = a14 ^ b_inv14 ^ c14;
  assign and14 = a14 & b14;
  assign or14  = a14 | b14;
  assign c15 = (a14 & b14) | (a14 & c14) | (b14 & c14);
  wire c_sub15;
  assign c_sub15 = (a14 & b_inv14) | (a14 & c14) | (b_inv14 & c14);
  wire s15, sub15, and15, or15;
  wire b_inv15;
  assign b_inv15 = ~b15;
  assign s15  = a15 ^ b15 ^ c15;
  assign sub15 = a15 ^ b_inv15 ^ c15;
  assign and15 = a15 & b15;
  assign or15  = a15 | b15;
  assign c16 = (a15 & b15) | (a15 & c15) | (b15 & c15);
  wire c_sub16;
  assign c_sub16 = (a15 & b_inv15) | (a15 & c15) | (b_inv15 & c15);
  wire s16, sub16, and16, or16;
  wire b_inv16;
  assign b_inv16 = ~b16;
  assign s16  = a16 ^ b16 ^ c16;
  assign sub16 = a16 ^ b_inv16 ^ c16;
  assign and16 = a16 & b16;
  assign or16  = a16 | b16;
  assign c17 = (a16 & b16) | (a16 & c16) | (b16 & c16);
  wire c_sub17;
  assign c_sub17 = (a16 & b_inv16) | (a16 & c16) | (b_inv16 & c16);
  wire s17, sub17, and17, or17;
  wire b_inv17;
  assign b_inv17 = ~b17;
  assign s17  = a17 ^ b17 ^ c17;
  assign sub17 = a17 ^ b_inv17 ^ c17;
  assign and17 = a17 & b17;
  assign or17  = a17 | b17;
  assign c18 = (a17 & b17) | (a17 & c17) | (b17 & c17);
  wire c_sub18;
  assign c_sub18 = (a17 & b_inv17) | (a17 & c17) | (b_inv17 & c17);
  wire s18, sub18, and18, or18;
  wire b_inv18;
  assign b_inv18 = ~b18;
  assign s18  = a18 ^ b18 ^ c18;
  assign sub18 = a18 ^ b_inv18 ^ c18;
  assign and18 = a18 & b18;
  assign or18  = a18 | b18;
  assign c19 = (a18 & b18) | (a18 & c18) | (b18 & c18);
  wire c_sub19;
  assign c_sub19 = (a18 & b_inv18) | (a18 & c18) | (b_inv18 & c18);
  wire s19, sub19, and19, or19;
  wire b_inv19;
  assign b_inv19 = ~b19;
  assign s19  = a19 ^ b19 ^ c19;
  assign sub19 = a19 ^ b_inv19 ^ c19;
  assign and19 = a19 & b19;
  assign or19  = a19 | b19;
  assign c20 = (a19 & b19) | (a19 & c19) | (b19 & c19);
  wire c_sub20;
  assign c_sub20 = (a19 & b_inv19) | (a19 & c19) | (b_inv19 & c19);
  wire s20, sub20, and20, or20;
  wire b_inv20;
  assign b_inv20 = ~b20;
  assign s20  = a20 ^ b20 ^ c20;
  assign sub20 = a20 ^ b_inv20 ^ c20;
  assign and20 = a20 & b20;
  assign or20  = a20 | b20;
  assign c21 = (a20 & b20) | (a20 & c20) | (b20 & c20);
  wire c_sub21;
  assign c_sub21 = (a20 & b_inv20) | (a20 & c20) | (b_inv20 & c20);
  wire s21, sub21, and21, or21;
  wire b_inv21;
  assign b_inv21 = ~b21;
  assign s21  = a21 ^ b21 ^ c21;
  assign sub21 = a21 ^ b_inv21 ^ c21;
  assign and21 = a21 & b21;
  assign or21  = a21 | b21;
  assign c22 = (a21 & b21) | (a21 & c21) | (b21 & c21);
  wire c_sub22;
  assign c_sub22 = (a21 & b_inv21) | (a21 & c21) | (b_inv21 & c21);
  wire s22, sub22, and22, or22;
  wire b_inv22;
  assign b_inv22 = ~b22;
  assign s22  = a22 ^ b22 ^ c22;
  assign sub22 = a22 ^ b_inv22 ^ c22;
  assign and22 = a22 & b22;
  assign or22  = a22 | b22;
  assign c23 = (a22 & b22) | (a22 & c22) | (b22 & c22);
  wire c_sub23;
  assign c_sub23 = (a22 & b_inv22) | (a22 & c22) | (b_inv22 & c22);
  wire s23, sub23, and23, or23;
  wire b_inv23;
  assign b_inv23 = ~b23;
  assign s23  = a23 ^ b23 ^ c23;
  assign sub23 = a23 ^ b_inv23 ^ c23;
  assign and23 = a23 & b23;
  assign or23  = a23 | b23;
  assign c24 = (a23 & b23) | (a23 & c23) | (b23 & c23);
  wire c_sub24;
  assign c_sub24 = (a23 & b_inv23) | (a23 & c23) | (b_inv23 & c23);
  wire s24, sub24, and24, or24;
  wire b_inv24;
  assign b_inv24 = ~b24;
  assign s24  = a24 ^ b24 ^ c24;
  assign sub24 = a24 ^ b_inv24 ^ c24;
  assign and24 = a24 & b24;
  assign or24  = a24 | b24;
  assign c25 = (a24 & b24) | (a24 & c24) | (b24 & c24);
  wire c_sub25;
  assign c_sub25 = (a24 & b_inv24) | (a24 & c24) | (b_inv24 & c24);
  wire s25, sub25, and25, or25;
  wire b_inv25;
  assign b_inv25 = ~b25;
  assign s25  = a25 ^ b25 ^ c25;
  assign sub25 = a25 ^ b_inv25 ^ c25;
  assign and25 = a25 & b25;
  assign or25  = a25 | b25;
  assign c26 = (a25 & b25) | (a25 & c25) | (b25 & c25);
  wire c_sub26;
  assign c_sub26 = (a25 & b_inv25) | (a25 & c25) | (b_inv25 & c25);
  wire s26, sub26, and26, or26;
  wire b_inv26;
  assign b_inv26 = ~b26;
  assign s26  = a26 ^ b26 ^ c26;
  assign sub26 = a26 ^ b_inv26 ^ c26;
  assign and26 = a26 & b26;
  assign or26  = a26 | b26;
  assign c27 = (a26 & b26) | (a26 & c26) | (b26 & c26);
  wire c_sub27;
  assign c_sub27 = (a26 & b_inv26) | (a26 & c26) | (b_inv26 & c26);
  wire s27, sub27, and27, or27;
  wire b_inv27;
  assign b_inv27 = ~b27;
  assign s27  = a27 ^ b27 ^ c27;
  assign sub27 = a27 ^ b_inv27 ^ c27;
  assign and27 = a27 & b27;
  assign or27  = a27 | b27;
  assign c28 = (a27 & b27) | (a27 & c27) | (b27 & c27);
  wire c_sub28;
  assign c_sub28 = (a27 & b_inv27) | (a27 & c27) | (b_inv27 & c27);
  wire s28, sub28, and28, or28;
  wire b_inv28;
  assign b_inv28 = ~b28;
  assign s28  = a28 ^ b28 ^ c28;
  assign sub28 = a28 ^ b_inv28 ^ c28;
  assign and28 = a28 & b28;
  assign or28  = a28 | b28;
  assign c29 = (a28 & b28) | (a28 & c28) | (b28 & c28);
  wire c_sub29;
  assign c_sub29 = (a28 & b_inv28) | (a28 & c28) | (b_inv28 & c28);
  wire s29, sub29, and29, or29;
  wire b_inv29;
  assign b_inv29 = ~b29;
  assign s29  = a29 ^ b29 ^ c29;
  assign sub29 = a29 ^ b_inv29 ^ c29;
  assign and29 = a29 & b29;
  assign or29  = a29 | b29;
  assign c30 = (a29 & b29) | (a29 & c29) | (b29 & c29);
  wire c_sub30;
  assign c_sub30 = (a29 & b_inv29) | (a29 & c29) | (b_inv29 & c29);
  wire s30, sub30, and30, or30;
  wire b_inv30;
  assign b_inv30 = ~b30;
  assign s30  = a30 ^ b30 ^ c30;
  assign sub30 = a30 ^ b_inv30 ^ c30;
  assign and30 = a30 & b30;
  assign or30  = a30 | b30;
  assign c31 = (a30 & b30) | (a30 & c30) | (b30 & c30);
  wire c_sub31;
  assign c_sub31 = (a30 & b_inv30) | (a30 & c30) | (b_inv30 & c30);
  wire s31, sub31, and31, or31;
  wire b_inv31;
  assign b_inv31 = ~b31;
  assign s31  = a31 ^ b31 ^ c31;
  assign sub31 = a31 ^ b_inv31 ^ c31;
  assign and31 = a31 & b31;
  assign or31  = a31 | b31;
  assign c32 = (a31 & b31) | (a31 & c31) | (b31 & c31);
  wire c_sub32;
  assign c_sub32 = (a31 & b_inv31) | (a31 & c31) | (b_inv31 & c31);
  wire s32, sub32, and32, or32;
  wire b_inv32;
  assign b_inv32 = ~b32;
  assign s32  = a32 ^ b32 ^ c32;
  assign sub32 = a32 ^ b_inv32 ^ c32;
  assign and32 = a32 & b32;
  assign or32  = a32 | b32;
  assign c33 = (a32 & b32) | (a32 & c32) | (b32 & c32);
  wire c_sub33;
  assign c_sub33 = (a32 & b_inv32) | (a32 & c32) | (b_inv32 & c32);
  wire s33, sub33, and33, or33;
  wire b_inv33;
  assign b_inv33 = ~b33;
  assign s33  = a33 ^ b33 ^ c33;
  assign sub33 = a33 ^ b_inv33 ^ c33;
  assign and33 = a33 & b33;
  assign or33  = a33 | b33;
  assign c34 = (a33 & b33) | (a33 & c33) | (b33 & c33);
  wire c_sub34;
  assign c_sub34 = (a33 & b_inv33) | (a33 & c33) | (b_inv33 & c33);
  wire s34, sub34, and34, or34;
  wire b_inv34;
  assign b_inv34 = ~b34;
  assign s34  = a34 ^ b34 ^ c34;
  assign sub34 = a34 ^ b_inv34 ^ c34;
  assign and34 = a34 & b34;
  assign or34  = a34 | b34;
  assign c35 = (a34 & b34) | (a34 & c34) | (b34 & c34);
  wire c_sub35;
  assign c_sub35 = (a34 & b_inv34) | (a34 & c34) | (b_inv34 & c34);
  wire s35, sub35, and35, or35;
  wire b_inv35;
  assign b_inv35 = ~b35;
  assign s35  = a35 ^ b35 ^ c35;
  assign sub35 = a35 ^ b_inv35 ^ c35;
  assign and35 = a35 & b35;
  assign or35  = a35 | b35;
  assign c36 = (a35 & b35) | (a35 & c35) | (b35 & c35);
  wire c_sub36;
  assign c_sub36 = (a35 & b_inv35) | (a35 & c35) | (b_inv35 & c35);
  wire s36, sub36, and36, or36;
  wire b_inv36;
  assign b_inv36 = ~b36;
  assign s36  = a36 ^ b36 ^ c36;
  assign sub36 = a36 ^ b_inv36 ^ c36;
  assign and36 = a36 & b36;
  assign or36  = a36 | b36;
  assign c37 = (a36 & b36) | (a36 & c36) | (b36 & c36);
  wire c_sub37;
  assign c_sub37 = (a36 & b_inv36) | (a36 & c36) | (b_inv36 & c36);
  wire s37, sub37, and37, or37;
  wire b_inv37;
  assign b_inv37 = ~b37;
  assign s37  = a37 ^ b37 ^ c37;
  assign sub37 = a37 ^ b_inv37 ^ c37;
  assign and37 = a37 & b37;
  assign or37  = a37 | b37;
  assign c38 = (a37 & b37) | (a37 & c37) | (b37 & c37);
  wire c_sub38;
  assign c_sub38 = (a37 & b_inv37) | (a37 & c37) | (b_inv37 & c37);
  wire s38, sub38, and38, or38;
  wire b_inv38;
  assign b_inv38 = ~b38;
  assign s38  = a38 ^ b38 ^ c38;
  assign sub38 = a38 ^ b_inv38 ^ c38;
  assign and38 = a38 & b38;
  assign or38  = a38 | b38;
  assign c39 = (a38 & b38) | (a38 & c38) | (b38 & c38);
  wire c_sub39;
  assign c_sub39 = (a38 & b_inv38) | (a38 & c38) | (b_inv38 & c38);
  wire s39, sub39, and39, or39;
  wire b_inv39;
  assign b_inv39 = ~b39;
  assign s39  = a39 ^ b39 ^ c39;
  assign sub39 = a39 ^ b_inv39 ^ c39;
  assign and39 = a39 & b39;
  assign or39  = a39 | b39;
  assign c40 = (a39 & b39) | (a39 & c39) | (b39 & c39);
  wire c_sub40;
  assign c_sub40 = (a39 & b_inv39) | (a39 & c39) | (b_inv39 & c39);
  wire s40, sub40, and40, or40;
  wire b_inv40;
  assign b_inv40 = ~b40;
  assign s40  = a40 ^ b40 ^ c40;
  assign sub40 = a40 ^ b_inv40 ^ c40;
  assign and40 = a40 & b40;
  assign or40  = a40 | b40;
  assign c41 = (a40 & b40) | (a40 & c40) | (b40 & c40);
  wire c_sub41;
  assign c_sub41 = (a40 & b_inv40) | (a40 & c40) | (b_inv40 & c40);
  wire s41, sub41, and41, or41;
  wire b_inv41;
  assign b_inv41 = ~b41;
  assign s41  = a41 ^ b41 ^ c41;
  assign sub41 = a41 ^ b_inv41 ^ c41;
  assign and41 = a41 & b41;
  assign or41  = a41 | b41;
  assign c42 = (a41 & b41) | (a41 & c41) | (b41 & c41);
  wire c_sub42;
  assign c_sub42 = (a41 & b_inv41) | (a41 & c41) | (b_inv41 & c41);
  wire s42, sub42, and42, or42;
  wire b_inv42;
  assign b_inv42 = ~b42;
  assign s42  = a42 ^ b42 ^ c42;
  assign sub42 = a42 ^ b_inv42 ^ c42;
  assign and42 = a42 & b42;
  assign or42  = a42 | b42;
  assign c43 = (a42 & b42) | (a42 & c42) | (b42 & c42);
  wire c_sub43;
  assign c_sub43 = (a42 & b_inv42) | (a42 & c42) | (b_inv42 & c42);
  wire s43, sub43, and43, or43;
  wire b_inv43;
  assign b_inv43 = ~b43;
  assign s43  = a43 ^ b43 ^ c43;
  assign sub43 = a43 ^ b_inv43 ^ c43;
  assign and43 = a43 & b43;
  assign or43  = a43 | b43;
  assign c44 = (a43 & b43) | (a43 & c43) | (b43 & c43);
  wire c_sub44;
  assign c_sub44 = (a43 & b_inv43) | (a43 & c43) | (b_inv43 & c43);
  wire s44, sub44, and44, or44;
  wire b_inv44;
  assign b_inv44 = ~b44;
  assign s44  = a44 ^ b44 ^ c44;
  assign sub44 = a44 ^ b_inv44 ^ c44;
  assign and44 = a44 & b44;
  assign or44  = a44 | b44;
  assign c45 = (a44 & b44) | (a44 & c44) | (b44 & c44);
  wire c_sub45;
  assign c_sub45 = (a44 & b_inv44) | (a44 & c44) | (b_inv44 & c44);
  wire s45, sub45, and45, or45;
  wire b_inv45;
  assign b_inv45 = ~b45;
  assign s45  = a45 ^ b45 ^ c45;
  assign sub45 = a45 ^ b_inv45 ^ c45;
  assign and45 = a45 & b45;
  assign or45  = a45 | b45;
  assign c46 = (a45 & b45) | (a45 & c45) | (b45 & c45);
  wire c_sub46;
  assign c_sub46 = (a45 & b_inv45) | (a45 & c45) | (b_inv45 & c45);
  wire s46, sub46, and46, or46;
  wire b_inv46;
  assign b_inv46 = ~b46;
  assign s46  = a46 ^ b46 ^ c46;
  assign sub46 = a46 ^ b_inv46 ^ c46;
  assign and46 = a46 & b46;
  assign or46  = a46 | b46;
  assign c47 = (a46 & b46) | (a46 & c46) | (b46 & c46);
  wire c_sub47;
  assign c_sub47 = (a46 & b_inv46) | (a46 & c46) | (b_inv46 & c46);
  wire s47, sub47, and47, or47;
  wire b_inv47;
  assign b_inv47 = ~b47;
  assign s47  = a47 ^ b47 ^ c47;
  assign sub47 = a47 ^ b_inv47 ^ c47;
  assign and47 = a47 & b47;
  assign or47  = a47 | b47;
  assign c48 = (a47 & b47) | (a47 & c47) | (b47 & c47);
  wire c_sub48;
  assign c_sub48 = (a47 & b_inv47) | (a47 & c47) | (b_inv47 & c47);
  wire s48, sub48, and48, or48;
  wire b_inv48;
  assign b_inv48 = ~b48;
  assign s48  = a48 ^ b48 ^ c48;
  assign sub48 = a48 ^ b_inv48 ^ c48;
  assign and48 = a48 & b48;
  assign or48  = a48 | b48;
  assign c49 = (a48 & b48) | (a48 & c48) | (b48 & c48);
  wire c_sub49;
  assign c_sub49 = (a48 & b_inv48) | (a48 & c48) | (b_inv48 & c48);
  wire s49, sub49, and49, or49;
  wire b_inv49;
  assign b_inv49 = ~b49;
  assign s49  = a49 ^ b49 ^ c49;
  assign sub49 = a49 ^ b_inv49 ^ c49;
  assign and49 = a49 & b49;
  assign or49  = a49 | b49;
  assign c50 = (a49 & b49) | (a49 & c49) | (b49 & c49);
  wire c_sub50;
  assign c_sub50 = (a49 & b_inv49) | (a49 & c49) | (b_inv49 & c49);
  wire s50, sub50, and50, or50;
  wire b_inv50;
  assign b_inv50 = ~b50;
  assign s50  = a50 ^ b50 ^ c50;
  assign sub50 = a50 ^ b_inv50 ^ c50;
  assign and50 = a50 & b50;
  assign or50  = a50 | b50;
  assign c51 = (a50 & b50) | (a50 & c50) | (b50 & c50);
  wire c_sub51;
  assign c_sub51 = (a50 & b_inv50) | (a50 & c50) | (b_inv50 & c50);
  wire s51, sub51, and51, or51;
  wire b_inv51;
  assign b_inv51 = ~b51;
  assign s51  = a51 ^ b51 ^ c51;
  assign sub51 = a51 ^ b_inv51 ^ c51;
  assign and51 = a51 & b51;
  assign or51  = a51 | b51;
  assign c52 = (a51 & b51) | (a51 & c51) | (b51 & c51);
  wire c_sub52;
  assign c_sub52 = (a51 & b_inv51) | (a51 & c51) | (b_inv51 & c51);
  wire s52, sub52, and52, or52;
  wire b_inv52;
  assign b_inv52 = ~b52;
  assign s52  = a52 ^ b52 ^ c52;
  assign sub52 = a52 ^ b_inv52 ^ c52;
  assign and52 = a52 & b52;
  assign or52  = a52 | b52;
  assign c53 = (a52 & b52) | (a52 & c52) | (b52 & c52);
  wire c_sub53;
  assign c_sub53 = (a52 & b_inv52) | (a52 & c52) | (b_inv52 & c52);
  wire s53, sub53, and53, or53;
  wire b_inv53;
  assign b_inv53 = ~b53;
  assign s53  = a53 ^ b53 ^ c53;
  assign sub53 = a53 ^ b_inv53 ^ c53;
  assign and53 = a53 & b53;
  assign or53  = a53 | b53;
  assign c54 = (a53 & b53) | (a53 & c53) | (b53 & c53);
  wire c_sub54;
  assign c_sub54 = (a53 & b_inv53) | (a53 & c53) | (b_inv53 & c53);
  wire s54, sub54, and54, or54;
  wire b_inv54;
  assign b_inv54 = ~b54;
  assign s54  = a54 ^ b54 ^ c54;
  assign sub54 = a54 ^ b_inv54 ^ c54;
  assign and54 = a54 & b54;
  assign or54  = a54 | b54;
  assign c55 = (a54 & b54) | (a54 & c54) | (b54 & c54);
  wire c_sub55;
  assign c_sub55 = (a54 & b_inv54) | (a54 & c54) | (b_inv54 & c54);
  wire s55, sub55, and55, or55;
  wire b_inv55;
  assign b_inv55 = ~b55;
  assign s55  = a55 ^ b55 ^ c55;
  assign sub55 = a55 ^ b_inv55 ^ c55;
  assign and55 = a55 & b55;
  assign or55  = a55 | b55;
  assign c56 = (a55 & b55) | (a55 & c55) | (b55 & c55);
  wire c_sub56;
  assign c_sub56 = (a55 & b_inv55) | (a55 & c55) | (b_inv55 & c55);
  wire s56, sub56, and56, or56;
  wire b_inv56;
  assign b_inv56 = ~b56;
  assign s56  = a56 ^ b56 ^ c56;
  assign sub56 = a56 ^ b_inv56 ^ c56;
  assign and56 = a56 & b56;
  assign or56  = a56 | b56;
  assign c57 = (a56 & b56) | (a56 & c56) | (b56 & c56);
  wire c_sub57;
  assign c_sub57 = (a56 & b_inv56) | (a56 & c56) | (b_inv56 & c56);
  wire s57, sub57, and57, or57;
  wire b_inv57;
  assign b_inv57 = ~b57;
  assign s57  = a57 ^ b57 ^ c57;
  assign sub57 = a57 ^ b_inv57 ^ c57;
  assign and57 = a57 & b57;
  assign or57  = a57 | b57;
  assign c58 = (a57 & b57) | (a57 & c57) | (b57 & c57);
  wire c_sub58;
  assign c_sub58 = (a57 & b_inv57) | (a57 & c57) | (b_inv57 & c57);
  wire s58, sub58, and58, or58;
  wire b_inv58;
  assign b_inv58 = ~b58;
  assign s58  = a58 ^ b58 ^ c58;
  assign sub58 = a58 ^ b_inv58 ^ c58;
  assign and58 = a58 & b58;
  assign or58  = a58 | b58;
  assign c59 = (a58 & b58) | (a58 & c58) | (b58 & c58);
  wire c_sub59;
  assign c_sub59 = (a58 & b_inv58) | (a58 & c58) | (b_inv58 & c58);
  wire s59, sub59, and59, or59;
  wire b_inv59;
  assign b_inv59 = ~b59;
  assign s59  = a59 ^ b59 ^ c59;
  assign sub59 = a59 ^ b_inv59 ^ c59;
  assign and59 = a59 & b59;
  assign or59  = a59 | b59;
  assign c60 = (a59 & b59) | (a59 & c59) | (b59 & c59);
  wire c_sub60;
  assign c_sub60 = (a59 & b_inv59) | (a59 & c59) | (b_inv59 & c59);
  wire s60, sub60, and60, or60;
  wire b_inv60;
  assign b_inv60 = ~b60;
  assign s60  = a60 ^ b60 ^ c60;
  assign sub60 = a60 ^ b_inv60 ^ c60;
  assign and60 = a60 & b60;
  assign or60  = a60 | b60;
  assign c61 = (a60 & b60) | (a60 & c60) | (b60 & c60);
  wire c_sub61;
  assign c_sub61 = (a60 & b_inv60) | (a60 & c60) | (b_inv60 & c60);
  wire s61, sub61, and61, or61;
  wire b_inv61;
  assign b_inv61 = ~b61;
  assign s61  = a61 ^ b61 ^ c61;
  assign sub61 = a61 ^ b_inv61 ^ c61;
  assign and61 = a61 & b61;
  assign or61  = a61 | b61;
  assign c62 = (a61 & b61) | (a61 & c61) | (b61 & c61);
  wire c_sub62;
  assign c_sub62 = (a61 & b_inv61) | (a61 & c61) | (b_inv61 & c61);
  wire s62, sub62, and62, or62;
  wire b_inv62;
  assign b_inv62 = ~b62;
  assign s62  = a62 ^ b62 ^ c62;
  assign sub62 = a62 ^ b_inv62 ^ c62;
  assign and62 = a62 & b62;
  assign or62  = a62 | b62;
  assign c63 = (a62 & b62) | (a62 & c62) | (b62 & c62);
  wire c_sub63;
  assign c_sub63 = (a62 & b_inv62) | (a62 & c62) | (b_inv62 & c62);
  wire s63, sub63, and63, or63;
  wire b_inv63;
  assign b_inv63 = ~b63;
  assign s63  = a63 ^ b63 ^ c63;
  assign sub63 = a63 ^ b_inv63 ^ c63;
  assign and63 = a63 & b63;
  assign or63  = a63 | b63;
  assign c64 = (a63 & b63) | (a63 & c63) | (b63 & c63);
  wire c_sub64;
  assign c_sub64 = (a63 & b_inv63) | (a63 & c63) | (b_inv63 & c63);
  wire s64, sub64, and64, or64;
  wire b_inv64;
  assign b_inv64 = ~b64;
  assign s64  = a64 ^ b64 ^ c64;
  assign sub64 = a64 ^ b_inv64 ^ c64;
  assign and64 = a64 & b64;
  assign or64  = a64 | b64;
  assign c65 = (a64 & b64) | (a64 & c64) | (b64 & c64);
  wire c_sub65;
  assign c_sub65 = (a64 & b_inv64) | (a64 & c64) | (b_inv64 & c64);
  wire s65, sub65, and65, or65;
  wire b_inv65;
  assign b_inv65 = ~b65;
  assign s65  = a65 ^ b65 ^ c65;
  assign sub65 = a65 ^ b_inv65 ^ c65;
  assign and65 = a65 & b65;
  assign or65  = a65 | b65;
  assign c66 = (a65 & b65) | (a65 & c65) | (b65 & c65);
  wire c_sub66;
  assign c_sub66 = (a65 & b_inv65) | (a65 & c65) | (b_inv65 & c65);
  wire s66, sub66, and66, or66;
  wire b_inv66;
  assign b_inv66 = ~b66;
  assign s66  = a66 ^ b66 ^ c66;
  assign sub66 = a66 ^ b_inv66 ^ c66;
  assign and66 = a66 & b66;
  assign or66  = a66 | b66;
  assign c67 = (a66 & b66) | (a66 & c66) | (b66 & c66);
  wire c_sub67;
  assign c_sub67 = (a66 & b_inv66) | (a66 & c66) | (b_inv66 & c66);
  wire s67, sub67, and67, or67;
  wire b_inv67;
  assign b_inv67 = ~b67;
  assign s67  = a67 ^ b67 ^ c67;
  assign sub67 = a67 ^ b_inv67 ^ c67;
  assign and67 = a67 & b67;
  assign or67  = a67 | b67;
  assign c68 = (a67 & b67) | (a67 & c67) | (b67 & c67);
  wire c_sub68;
  assign c_sub68 = (a67 & b_inv67) | (a67 & c67) | (b_inv67 & c67);
  wire s68, sub68, and68, or68;
  wire b_inv68;
  assign b_inv68 = ~b68;
  assign s68  = a68 ^ b68 ^ c68;
  assign sub68 = a68 ^ b_inv68 ^ c68;
  assign and68 = a68 & b68;
  assign or68  = a68 | b68;
  assign c69 = (a68 & b68) | (a68 & c68) | (b68 & c68);
  wire c_sub69;
  assign c_sub69 = (a68 & b_inv68) | (a68 & c68) | (b_inv68 & c68);
  wire s69, sub69, and69, or69;
  wire b_inv69;
  assign b_inv69 = ~b69;
  assign s69  = a69 ^ b69 ^ c69;
  assign sub69 = a69 ^ b_inv69 ^ c69;
  assign and69 = a69 & b69;
  assign or69  = a69 | b69;
  assign c70 = (a69 & b69) | (a69 & c69) | (b69 & c69);
  wire c_sub70;
  assign c_sub70 = (a69 & b_inv69) | (a69 & c69) | (b_inv69 & c69);
  wire s70, sub70, and70, or70;
  wire b_inv70;
  assign b_inv70 = ~b70;
  assign s70  = a70 ^ b70 ^ c70;
  assign sub70 = a70 ^ b_inv70 ^ c70;
  assign and70 = a70 & b70;
  assign or70  = a70 | b70;
  assign c71 = (a70 & b70) | (a70 & c70) | (b70 & c70);
  wire c_sub71;
  assign c_sub71 = (a70 & b_inv70) | (a70 & c70) | (b_inv70 & c70);
  wire s71, sub71, and71, or71;
  wire b_inv71;
  assign b_inv71 = ~b71;
  assign s71  = a71 ^ b71 ^ c71;
  assign sub71 = a71 ^ b_inv71 ^ c71;
  assign and71 = a71 & b71;
  assign or71  = a71 | b71;
  assign c72 = (a71 & b71) | (a71 & c71) | (b71 & c71);
  wire c_sub72;
  assign c_sub72 = (a71 & b_inv71) | (a71 & c71) | (b_inv71 & c71);
  wire s72, sub72, and72, or72;
  wire b_inv72;
  assign b_inv72 = ~b72;
  assign s72  = a72 ^ b72 ^ c72;
  assign sub72 = a72 ^ b_inv72 ^ c72;
  assign and72 = a72 & b72;
  assign or72  = a72 | b72;
  assign c73 = (a72 & b72) | (a72 & c72) | (b72 & c72);
  wire c_sub73;
  assign c_sub73 = (a72 & b_inv72) | (a72 & c72) | (b_inv72 & c72);
  wire s73, sub73, and73, or73;
  wire b_inv73;
  assign b_inv73 = ~b73;
  assign s73  = a73 ^ b73 ^ c73;
  assign sub73 = a73 ^ b_inv73 ^ c73;
  assign and73 = a73 & b73;
  assign or73  = a73 | b73;
  assign c74 = (a73 & b73) | (a73 & c73) | (b73 & c73);
  wire c_sub74;
  assign c_sub74 = (a73 & b_inv73) | (a73 & c73) | (b_inv73 & c73);
  wire s74, sub74, and74, or74;
  wire b_inv74;
  assign b_inv74 = ~b74;
  assign s74  = a74 ^ b74 ^ c74;
  assign sub74 = a74 ^ b_inv74 ^ c74;
  assign and74 = a74 & b74;
  assign or74  = a74 | b74;
  assign c75 = (a74 & b74) | (a74 & c74) | (b74 & c74);
  wire c_sub75;
  assign c_sub75 = (a74 & b_inv74) | (a74 & c74) | (b_inv74 & c74);
  wire s75, sub75, and75, or75;
  wire b_inv75;
  assign b_inv75 = ~b75;
  assign s75  = a75 ^ b75 ^ c75;
  assign sub75 = a75 ^ b_inv75 ^ c75;
  assign and75 = a75 & b75;
  assign or75  = a75 | b75;
  assign c76 = (a75 & b75) | (a75 & c75) | (b75 & c75);
  wire c_sub76;
  assign c_sub76 = (a75 & b_inv75) | (a75 & c75) | (b_inv75 & c75);
  wire s76, sub76, and76, or76;
  wire b_inv76;
  assign b_inv76 = ~b76;
  assign s76  = a76 ^ b76 ^ c76;
  assign sub76 = a76 ^ b_inv76 ^ c76;
  assign and76 = a76 & b76;
  assign or76  = a76 | b76;
  assign c77 = (a76 & b76) | (a76 & c76) | (b76 & c76);
  wire c_sub77;
  assign c_sub77 = (a76 & b_inv76) | (a76 & c76) | (b_inv76 & c76);
  wire s77, sub77, and77, or77;
  wire b_inv77;
  assign b_inv77 = ~b77;
  assign s77  = a77 ^ b77 ^ c77;
  assign sub77 = a77 ^ b_inv77 ^ c77;
  assign and77 = a77 & b77;
  assign or77  = a77 | b77;
  assign c78 = (a77 & b77) | (a77 & c77) | (b77 & c77);
  wire c_sub78;
  assign c_sub78 = (a77 & b_inv77) | (a77 & c77) | (b_inv77 & c77);
  wire s78, sub78, and78, or78;
  wire b_inv78;
  assign b_inv78 = ~b78;
  assign s78  = a78 ^ b78 ^ c78;
  assign sub78 = a78 ^ b_inv78 ^ c78;
  assign and78 = a78 & b78;
  assign or78  = a78 | b78;
  assign c79 = (a78 & b78) | (a78 & c78) | (b78 & c78);
  wire c_sub79;
  assign c_sub79 = (a78 & b_inv78) | (a78 & c78) | (b_inv78 & c78);
  wire s79, sub79, and79, or79;
  wire b_inv79;
  assign b_inv79 = ~b79;
  assign s79  = a79 ^ b79 ^ c79;
  assign sub79 = a79 ^ b_inv79 ^ c79;
  assign and79 = a79 & b79;
  assign or79  = a79 | b79;
  assign c80 = (a79 & b79) | (a79 & c79) | (b79 & c79);
  wire c_sub80;
  assign c_sub80 = (a79 & b_inv79) | (a79 & c79) | (b_inv79 & c79);
  wire s80, sub80, and80, or80;
  wire b_inv80;
  assign b_inv80 = ~b80;
  assign s80  = a80 ^ b80 ^ c80;
  assign sub80 = a80 ^ b_inv80 ^ c80;
  assign and80 = a80 & b80;
  assign or80  = a80 | b80;
  assign c81 = (a80 & b80) | (a80 & c80) | (b80 & c80);
  wire c_sub81;
  assign c_sub81 = (a80 & b_inv80) | (a80 & c80) | (b_inv80 & c80);
  wire s81, sub81, and81, or81;
  wire b_inv81;
  assign b_inv81 = ~b81;
  assign s81  = a81 ^ b81 ^ c81;
  assign sub81 = a81 ^ b_inv81 ^ c81;
  assign and81 = a81 & b81;
  assign or81  = a81 | b81;
  assign c82 = (a81 & b81) | (a81 & c81) | (b81 & c81);
  wire c_sub82;
  assign c_sub82 = (a81 & b_inv81) | (a81 & c81) | (b_inv81 & c81);
  wire s82, sub82, and82, or82;
  wire b_inv82;
  assign b_inv82 = ~b82;
  assign s82  = a82 ^ b82 ^ c82;
  assign sub82 = a82 ^ b_inv82 ^ c82;
  assign and82 = a82 & b82;
  assign or82  = a82 | b82;
  assign c83 = (a82 & b82) | (a82 & c82) | (b82 & c82);
  wire c_sub83;
  assign c_sub83 = (a82 & b_inv82) | (a82 & c82) | (b_inv82 & c82);
  wire s83, sub83, and83, or83;
  wire b_inv83;
  assign b_inv83 = ~b83;
  assign s83  = a83 ^ b83 ^ c83;
  assign sub83 = a83 ^ b_inv83 ^ c83;
  assign and83 = a83 & b83;
  assign or83  = a83 | b83;
  assign c84 = (a83 & b83) | (a83 & c83) | (b83 & c83);
  wire c_sub84;
  assign c_sub84 = (a83 & b_inv83) | (a83 & c83) | (b_inv83 & c83);
  wire s84, sub84, and84, or84;
  wire b_inv84;
  assign b_inv84 = ~b84;
  assign s84  = a84 ^ b84 ^ c84;
  assign sub84 = a84 ^ b_inv84 ^ c84;
  assign and84 = a84 & b84;
  assign or84  = a84 | b84;
  assign c85 = (a84 & b84) | (a84 & c84) | (b84 & c84);
  wire c_sub85;
  assign c_sub85 = (a84 & b_inv84) | (a84 & c84) | (b_inv84 & c84);
  wire s85, sub85, and85, or85;
  wire b_inv85;
  assign b_inv85 = ~b85;
  assign s85  = a85 ^ b85 ^ c85;
  assign sub85 = a85 ^ b_inv85 ^ c85;
  assign and85 = a85 & b85;
  assign or85  = a85 | b85;
  assign c86 = (a85 & b85) | (a85 & c85) | (b85 & c85);
  wire c_sub86;
  assign c_sub86 = (a85 & b_inv85) | (a85 & c85) | (b_inv85 & c85);
  wire s86, sub86, and86, or86;
  wire b_inv86;
  assign b_inv86 = ~b86;
  assign s86  = a86 ^ b86 ^ c86;
  assign sub86 = a86 ^ b_inv86 ^ c86;
  assign and86 = a86 & b86;
  assign or86  = a86 | b86;
  assign c87 = (a86 & b86) | (a86 & c86) | (b86 & c86);
  wire c_sub87;
  assign c_sub87 = (a86 & b_inv86) | (a86 & c86) | (b_inv86 & c86);
  wire s87, sub87, and87, or87;
  wire b_inv87;
  assign b_inv87 = ~b87;
  assign s87  = a87 ^ b87 ^ c87;
  assign sub87 = a87 ^ b_inv87 ^ c87;
  assign and87 = a87 & b87;
  assign or87  = a87 | b87;
  assign c88 = (a87 & b87) | (a87 & c87) | (b87 & c87);
  wire c_sub88;
  assign c_sub88 = (a87 & b_inv87) | (a87 & c87) | (b_inv87 & c87);
  wire s88, sub88, and88, or88;
  wire b_inv88;
  assign b_inv88 = ~b88;
  assign s88  = a88 ^ b88 ^ c88;
  assign sub88 = a88 ^ b_inv88 ^ c88;
  assign and88 = a88 & b88;
  assign or88  = a88 | b88;
  assign c89 = (a88 & b88) | (a88 & c88) | (b88 & c88);
  wire c_sub89;
  assign c_sub89 = (a88 & b_inv88) | (a88 & c88) | (b_inv88 & c88);
  wire s89, sub89, and89, or89;
  wire b_inv89;
  assign b_inv89 = ~b89;
  assign s89  = a89 ^ b89 ^ c89;
  assign sub89 = a89 ^ b_inv89 ^ c89;
  assign and89 = a89 & b89;
  assign or89  = a89 | b89;
  assign c90 = (a89 & b89) | (a89 & c89) | (b89 & c89);
  wire c_sub90;
  assign c_sub90 = (a89 & b_inv89) | (a89 & c89) | (b_inv89 & c89);
  wire s90, sub90, and90, or90;
  wire b_inv90;
  assign b_inv90 = ~b90;
  assign s90  = a90 ^ b90 ^ c90;
  assign sub90 = a90 ^ b_inv90 ^ c90;
  assign and90 = a90 & b90;
  assign or90  = a90 | b90;
  assign c91 = (a90 & b90) | (a90 & c90) | (b90 & c90);
  wire c_sub91;
  assign c_sub91 = (a90 & b_inv90) | (a90 & c90) | (b_inv90 & c90);
  wire s91, sub91, and91, or91;
  wire b_inv91;
  assign b_inv91 = ~b91;
  assign s91  = a91 ^ b91 ^ c91;
  assign sub91 = a91 ^ b_inv91 ^ c91;
  assign and91 = a91 & b91;
  assign or91  = a91 | b91;
  assign c92 = (a91 & b91) | (a91 & c91) | (b91 & c91);
  wire c_sub92;
  assign c_sub92 = (a91 & b_inv91) | (a91 & c91) | (b_inv91 & c91);
  wire s92, sub92, and92, or92;
  wire b_inv92;
  assign b_inv92 = ~b92;
  assign s92  = a92 ^ b92 ^ c92;
  assign sub92 = a92 ^ b_inv92 ^ c92;
  assign and92 = a92 & b92;
  assign or92  = a92 | b92;
  assign c93 = (a92 & b92) | (a92 & c92) | (b92 & c92);
  wire c_sub93;
  assign c_sub93 = (a92 & b_inv92) | (a92 & c92) | (b_inv92 & c92);
  wire s93, sub93, and93, or93;
  wire b_inv93;
  assign b_inv93 = ~b93;
  assign s93  = a93 ^ b93 ^ c93;
  assign sub93 = a93 ^ b_inv93 ^ c93;
  assign and93 = a93 & b93;
  assign or93  = a93 | b93;
  assign c94 = (a93 & b93) | (a93 & c93) | (b93 & c93);
  wire c_sub94;
  assign c_sub94 = (a93 & b_inv93) | (a93 & c93) | (b_inv93 & c93);
  wire s94, sub94, and94, or94;
  wire b_inv94;
  assign b_inv94 = ~b94;
  assign s94  = a94 ^ b94 ^ c94;
  assign sub94 = a94 ^ b_inv94 ^ c94;
  assign and94 = a94 & b94;
  assign or94  = a94 | b94;
  assign c95 = (a94 & b94) | (a94 & c94) | (b94 & c94);
  wire c_sub95;
  assign c_sub95 = (a94 & b_inv94) | (a94 & c94) | (b_inv94 & c94);
  wire s95, sub95, and95, or95;
  wire b_inv95;
  assign b_inv95 = ~b95;
  assign s95  = a95 ^ b95 ^ c95;
  assign sub95 = a95 ^ b_inv95 ^ c95;
  assign and95 = a95 & b95;
  assign or95  = a95 | b95;
  assign c96 = (a95 & b95) | (a95 & c95) | (b95 & c95);
  wire c_sub96;
  assign c_sub96 = (a95 & b_inv95) | (a95 & c95) | (b_inv95 & c95);
  wire s96, sub96, and96, or96;
  wire b_inv96;
  assign b_inv96 = ~b96;
  assign s96  = a96 ^ b96 ^ c96;
  assign sub96 = a96 ^ b_inv96 ^ c96;
  assign and96 = a96 & b96;
  assign or96  = a96 | b96;
  assign c97 = (a96 & b96) | (a96 & c96) | (b96 & c96);
  wire c_sub97;
  assign c_sub97 = (a96 & b_inv96) | (a96 & c96) | (b_inv96 & c96);
  wire s97, sub97, and97, or97;
  wire b_inv97;
  assign b_inv97 = ~b97;
  assign s97  = a97 ^ b97 ^ c97;
  assign sub97 = a97 ^ b_inv97 ^ c97;
  assign and97 = a97 & b97;
  assign or97  = a97 | b97;
  assign c98 = (a97 & b97) | (a97 & c97) | (b97 & c97);
  wire c_sub98;
  assign c_sub98 = (a97 & b_inv97) | (a97 & c97) | (b_inv97 & c97);
  wire s98, sub98, and98, or98;
  wire b_inv98;
  assign b_inv98 = ~b98;
  assign s98  = a98 ^ b98 ^ c98;
  assign sub98 = a98 ^ b_inv98 ^ c98;
  assign and98 = a98 & b98;
  assign or98  = a98 | b98;
  assign c99 = (a98 & b98) | (a98 & c98) | (b98 & c98);
  wire c_sub99;
  assign c_sub99 = (a98 & b_inv98) | (a98 & c98) | (b_inv98 & c98);
  wire s99, sub99, and99, or99;
  wire b_inv99;
  assign b_inv99 = ~b99;
  assign s99  = a99 ^ b99 ^ c99;
  assign sub99 = a99 ^ b_inv99 ^ c99;
  assign and99 = a99 & b99;
  assign or99  = a99 | b99;
  assign c100 = (a99 & b99) | (a99 & c99) | (b99 & c99);
  wire c_sub100;
  assign c_sub100 = (a99 & b_inv99) | (a99 & c99) | (b_inv99 & c99);
  wire s100, sub100, and100, or100;
  wire b_inv100;
  assign b_inv100 = ~b100;
  assign s100  = a100 ^ b100 ^ c100;
  assign sub100 = a100 ^ b_inv100 ^ c100;
  assign and100 = a100 & b100;
  assign or100  = a100 | b100;
  assign c101 = (a100 & b100) | (a100 & c100) | (b100 & c100);
  wire c_sub101;
  assign c_sub101 = (a100 & b_inv100) | (a100 & c100) | (b_inv100 & c100);
  wire s101, sub101, and101, or101;
  wire b_inv101;
  assign b_inv101 = ~b101;
  assign s101  = a101 ^ b101 ^ c101;
  assign sub101 = a101 ^ b_inv101 ^ c101;
  assign and101 = a101 & b101;
  assign or101  = a101 | b101;
  assign c102 = (a101 & b101) | (a101 & c101) | (b101 & c101);
  wire c_sub102;
  assign c_sub102 = (a101 & b_inv101) | (a101 & c101) | (b_inv101 & c101);
  wire s102, sub102, and102, or102;
  wire b_inv102;
  assign b_inv102 = ~b102;
  assign s102  = a102 ^ b102 ^ c102;
  assign sub102 = a102 ^ b_inv102 ^ c102;
  assign and102 = a102 & b102;
  assign or102  = a102 | b102;
  assign c103 = (a102 & b102) | (a102 & c102) | (b102 & c102);
  wire c_sub103;
  assign c_sub103 = (a102 & b_inv102) | (a102 & c102) | (b_inv102 & c102);
  wire s103, sub103, and103, or103;
  wire b_inv103;
  assign b_inv103 = ~b103;
  assign s103  = a103 ^ b103 ^ c103;
  assign sub103 = a103 ^ b_inv103 ^ c103;
  assign and103 = a103 & b103;
  assign or103  = a103 | b103;
  assign c104 = (a103 & b103) | (a103 & c103) | (b103 & c103);
  wire c_sub104;
  assign c_sub104 = (a103 & b_inv103) | (a103 & c103) | (b_inv103 & c103);
  wire s104, sub104, and104, or104;
  wire b_inv104;
  assign b_inv104 = ~b104;
  assign s104  = a104 ^ b104 ^ c104;
  assign sub104 = a104 ^ b_inv104 ^ c104;
  assign and104 = a104 & b104;
  assign or104  = a104 | b104;
  assign c105 = (a104 & b104) | (a104 & c104) | (b104 & c104);
  wire c_sub105;
  assign c_sub105 = (a104 & b_inv104) | (a104 & c104) | (b_inv104 & c104);
  wire s105, sub105, and105, or105;
  wire b_inv105;
  assign b_inv105 = ~b105;
  assign s105  = a105 ^ b105 ^ c105;
  assign sub105 = a105 ^ b_inv105 ^ c105;
  assign and105 = a105 & b105;
  assign or105  = a105 | b105;
  assign c106 = (a105 & b105) | (a105 & c105) | (b105 & c105);
  wire c_sub106;
  assign c_sub106 = (a105 & b_inv105) | (a105 & c105) | (b_inv105 & c105);
  wire s106, sub106, and106, or106;
  wire b_inv106;
  assign b_inv106 = ~b106;
  assign s106  = a106 ^ b106 ^ c106;
  assign sub106 = a106 ^ b_inv106 ^ c106;
  assign and106 = a106 & b106;
  assign or106  = a106 | b106;
  assign c107 = (a106 & b106) | (a106 & c106) | (b106 & c106);
  wire c_sub107;
  assign c_sub107 = (a106 & b_inv106) | (a106 & c106) | (b_inv106 & c106);
  wire s107, sub107, and107, or107;
  wire b_inv107;
  assign b_inv107 = ~b107;
  assign s107  = a107 ^ b107 ^ c107;
  assign sub107 = a107 ^ b_inv107 ^ c107;
  assign and107 = a107 & b107;
  assign or107  = a107 | b107;
  assign c108 = (a107 & b107) | (a107 & c107) | (b107 & c107);
  wire c_sub108;
  assign c_sub108 = (a107 & b_inv107) | (a107 & c107) | (b_inv107 & c107);
  wire s108, sub108, and108, or108;
  wire b_inv108;
  assign b_inv108 = ~b108;
  assign s108  = a108 ^ b108 ^ c108;
  assign sub108 = a108 ^ b_inv108 ^ c108;
  assign and108 = a108 & b108;
  assign or108  = a108 | b108;
  assign c109 = (a108 & b108) | (a108 & c108) | (b108 & c108);
  wire c_sub109;
  assign c_sub109 = (a108 & b_inv108) | (a108 & c108) | (b_inv108 & c108);
  wire s109, sub109, and109, or109;
  wire b_inv109;
  assign b_inv109 = ~b109;
  assign s109  = a109 ^ b109 ^ c109;
  assign sub109 = a109 ^ b_inv109 ^ c109;
  assign and109 = a109 & b109;
  assign or109  = a109 | b109;
  assign c110 = (a109 & b109) | (a109 & c109) | (b109 & c109);
  wire c_sub110;
  assign c_sub110 = (a109 & b_inv109) | (a109 & c109) | (b_inv109 & c109);
  wire s110, sub110, and110, or110;
  wire b_inv110;
  assign b_inv110 = ~b110;
  assign s110  = a110 ^ b110 ^ c110;
  assign sub110 = a110 ^ b_inv110 ^ c110;
  assign and110 = a110 & b110;
  assign or110  = a110 | b110;
  assign c111 = (a110 & b110) | (a110 & c110) | (b110 & c110);
  wire c_sub111;
  assign c_sub111 = (a110 & b_inv110) | (a110 & c110) | (b_inv110 & c110);
  wire s111, sub111, and111, or111;
  wire b_inv111;
  assign b_inv111 = ~b111;
  assign s111  = a111 ^ b111 ^ c111;
  assign sub111 = a111 ^ b_inv111 ^ c111;
  assign and111 = a111 & b111;
  assign or111  = a111 | b111;
  assign c112 = (a111 & b111) | (a111 & c111) | (b111 & c111);
  wire c_sub112;
  assign c_sub112 = (a111 & b_inv111) | (a111 & c111) | (b_inv111 & c111);
  wire s112, sub112, and112, or112;
  wire b_inv112;
  assign b_inv112 = ~b112;
  assign s112  = a112 ^ b112 ^ c112;
  assign sub112 = a112 ^ b_inv112 ^ c112;
  assign and112 = a112 & b112;
  assign or112  = a112 | b112;
  assign c113 = (a112 & b112) | (a112 & c112) | (b112 & c112);
  wire c_sub113;
  assign c_sub113 = (a112 & b_inv112) | (a112 & c112) | (b_inv112 & c112);
  wire s113, sub113, and113, or113;
  wire b_inv113;
  assign b_inv113 = ~b113;
  assign s113  = a113 ^ b113 ^ c113;
  assign sub113 = a113 ^ b_inv113 ^ c113;
  assign and113 = a113 & b113;
  assign or113  = a113 | b113;
  assign c114 = (a113 & b113) | (a113 & c113) | (b113 & c113);
  wire c_sub114;
  assign c_sub114 = (a113 & b_inv113) | (a113 & c113) | (b_inv113 & c113);
  wire s114, sub114, and114, or114;
  wire b_inv114;
  assign b_inv114 = ~b114;
  assign s114  = a114 ^ b114 ^ c114;
  assign sub114 = a114 ^ b_inv114 ^ c114;
  assign and114 = a114 & b114;
  assign or114  = a114 | b114;
  assign c115 = (a114 & b114) | (a114 & c114) | (b114 & c114);
  wire c_sub115;
  assign c_sub115 = (a114 & b_inv114) | (a114 & c114) | (b_inv114 & c114);
  wire s115, sub115, and115, or115;
  wire b_inv115;
  assign b_inv115 = ~b115;
  assign s115  = a115 ^ b115 ^ c115;
  assign sub115 = a115 ^ b_inv115 ^ c115;
  assign and115 = a115 & b115;
  assign or115  = a115 | b115;
  assign c116 = (a115 & b115) | (a115 & c115) | (b115 & c115);
  wire c_sub116;
  assign c_sub116 = (a115 & b_inv115) | (a115 & c115) | (b_inv115 & c115);
  wire s116, sub116, and116, or116;
  wire b_inv116;
  assign b_inv116 = ~b116;
  assign s116  = a116 ^ b116 ^ c116;
  assign sub116 = a116 ^ b_inv116 ^ c116;
  assign and116 = a116 & b116;
  assign or116  = a116 | b116;
  assign c117 = (a116 & b116) | (a116 & c116) | (b116 & c116);
  wire c_sub117;
  assign c_sub117 = (a116 & b_inv116) | (a116 & c116) | (b_inv116 & c116);
  wire s117, sub117, and117, or117;
  wire b_inv117;
  assign b_inv117 = ~b117;
  assign s117  = a117 ^ b117 ^ c117;
  assign sub117 = a117 ^ b_inv117 ^ c117;
  assign and117 = a117 & b117;
  assign or117  = a117 | b117;
  assign c118 = (a117 & b117) | (a117 & c117) | (b117 & c117);
  wire c_sub118;
  assign c_sub118 = (a117 & b_inv117) | (a117 & c117) | (b_inv117 & c117);
  wire s118, sub118, and118, or118;
  wire b_inv118;
  assign b_inv118 = ~b118;
  assign s118  = a118 ^ b118 ^ c118;
  assign sub118 = a118 ^ b_inv118 ^ c118;
  assign and118 = a118 & b118;
  assign or118  = a118 | b118;
  assign c119 = (a118 & b118) | (a118 & c118) | (b118 & c118);
  wire c_sub119;
  assign c_sub119 = (a118 & b_inv118) | (a118 & c118) | (b_inv118 & c118);
  wire s119, sub119, and119, or119;
  wire b_inv119;
  assign b_inv119 = ~b119;
  assign s119  = a119 ^ b119 ^ c119;
  assign sub119 = a119 ^ b_inv119 ^ c119;
  assign and119 = a119 & b119;
  assign or119  = a119 | b119;
  assign c120 = (a119 & b119) | (a119 & c119) | (b119 & c119);
  wire c_sub120;
  assign c_sub120 = (a119 & b_inv119) | (a119 & c119) | (b_inv119 & c119);
  wire s120, sub120, and120, or120;
  wire b_inv120;
  assign b_inv120 = ~b120;
  assign s120  = a120 ^ b120 ^ c120;
  assign sub120 = a120 ^ b_inv120 ^ c120;
  assign and120 = a120 & b120;
  assign or120  = a120 | b120;
  assign c121 = (a120 & b120) | (a120 & c120) | (b120 & c120);
  wire c_sub121;
  assign c_sub121 = (a120 & b_inv120) | (a120 & c120) | (b_inv120 & c120);
  wire s121, sub121, and121, or121;
  wire b_inv121;
  assign b_inv121 = ~b121;
  assign s121  = a121 ^ b121 ^ c121;
  assign sub121 = a121 ^ b_inv121 ^ c121;
  assign and121 = a121 & b121;
  assign or121  = a121 | b121;
  assign c122 = (a121 & b121) | (a121 & c121) | (b121 & c121);
  wire c_sub122;
  assign c_sub122 = (a121 & b_inv121) | (a121 & c121) | (b_inv121 & c121);
  wire s122, sub122, and122, or122;
  wire b_inv122;
  assign b_inv122 = ~b122;
  assign s122  = a122 ^ b122 ^ c122;
  assign sub122 = a122 ^ b_inv122 ^ c122;
  assign and122 = a122 & b122;
  assign or122  = a122 | b122;
  assign c123 = (a122 & b122) | (a122 & c122) | (b122 & c122);
  wire c_sub123;
  assign c_sub123 = (a122 & b_inv122) | (a122 & c122) | (b_inv122 & c122);
  wire s123, sub123, and123, or123;
  wire b_inv123;
  assign b_inv123 = ~b123;
  assign s123  = a123 ^ b123 ^ c123;
  assign sub123 = a123 ^ b_inv123 ^ c123;
  assign and123 = a123 & b123;
  assign or123  = a123 | b123;
  assign c124 = (a123 & b123) | (a123 & c123) | (b123 & c123);
  wire c_sub124;
  assign c_sub124 = (a123 & b_inv123) | (a123 & c123) | (b_inv123 & c123);
  wire s124, sub124, and124, or124;
  wire b_inv124;
  assign b_inv124 = ~b124;
  assign s124  = a124 ^ b124 ^ c124;
  assign sub124 = a124 ^ b_inv124 ^ c124;
  assign and124 = a124 & b124;
  assign or124  = a124 | b124;
  assign c125 = (a124 & b124) | (a124 & c124) | (b124 & c124);
  wire c_sub125;
  assign c_sub125 = (a124 & b_inv124) | (a124 & c124) | (b_inv124 & c124);
  wire s125, sub125, and125, or125;
  wire b_inv125;
  assign b_inv125 = ~b125;
  assign s125  = a125 ^ b125 ^ c125;
  assign sub125 = a125 ^ b_inv125 ^ c125;
  assign and125 = a125 & b125;
  assign or125  = a125 | b125;
  assign c126 = (a125 & b125) | (a125 & c125) | (b125 & c125);
  wire c_sub126;
  assign c_sub126 = (a125 & b_inv125) | (a125 & c125) | (b_inv125 & c125);
  wire s126, sub126, and126, or126;
  wire b_inv126;
  assign b_inv126 = ~b126;
  assign s126  = a126 ^ b126 ^ c126;
  assign sub126 = a126 ^ b_inv126 ^ c126;
  assign and126 = a126 & b126;
  assign or126  = a126 | b126;
  assign c127 = (a126 & b126) | (a126 & c126) | (b126 & c126);
  wire c_sub127;
  assign c_sub127 = (a126 & b_inv126) | (a126 & c126) | (b_inv126 & c126);
  wire s127, sub127, and127, or127;
  wire b_inv127;
  assign b_inv127 = ~b127;
  assign s127  = a127 ^ b127 ^ c127;
  assign sub127 = a127 ^ b_inv127 ^ c127;
  assign and127 = a127 & b127;
  assign or127  = a127 | b127;
  assign c128 = (a127 & b127) | (a127 & c127) | (b127 & c127);
  wire c_sub128;
  assign c_sub128 = (a127 & b_inv127) | (a127 & c127) | (b_inv127 & c127);
  wire s128, sub128, and128, or128;
  wire b_inv128;
  assign b_inv128 = ~b128;
  assign s128  = a128 ^ b128 ^ c128;
  assign sub128 = a128 ^ b_inv128 ^ c128;
  assign and128 = a128 & b128;
  assign or128  = a128 | b128;
  assign c129 = (a128 & b128) | (a128 & c128) | (b128 & c128);
  wire c_sub129;
  assign c_sub129 = (a128 & b_inv128) | (a128 & c128) | (b_inv128 & c128);
  wire s129, sub129, and129, or129;
  wire b_inv129;
  assign b_inv129 = ~b129;
  assign s129  = a129 ^ b129 ^ c129;
  assign sub129 = a129 ^ b_inv129 ^ c129;
  assign and129 = a129 & b129;
  assign or129  = a129 | b129;
  assign c130 = (a129 & b129) | (a129 & c129) | (b129 & c129);
  wire c_sub130;
  assign c_sub130 = (a129 & b_inv129) | (a129 & c129) | (b_inv129 & c129);
  wire s130, sub130, and130, or130;
  wire b_inv130;
  assign b_inv130 = ~b130;
  assign s130  = a130 ^ b130 ^ c130;
  assign sub130 = a130 ^ b_inv130 ^ c130;
  assign and130 = a130 & b130;
  assign or130  = a130 | b130;
  assign c131 = (a130 & b130) | (a130 & c130) | (b130 & c130);
  wire c_sub131;
  assign c_sub131 = (a130 & b_inv130) | (a130 & c130) | (b_inv130 & c130);
  wire s131, sub131, and131, or131;
  wire b_inv131;
  assign b_inv131 = ~b131;
  assign s131  = a131 ^ b131 ^ c131;
  assign sub131 = a131 ^ b_inv131 ^ c131;
  assign and131 = a131 & b131;
  assign or131  = a131 | b131;
  assign c132 = (a131 & b131) | (a131 & c131) | (b131 & c131);
  wire c_sub132;
  assign c_sub132 = (a131 & b_inv131) | (a131 & c131) | (b_inv131 & c131);
  wire s132, sub132, and132, or132;
  wire b_inv132;
  assign b_inv132 = ~b132;
  assign s132  = a132 ^ b132 ^ c132;
  assign sub132 = a132 ^ b_inv132 ^ c132;
  assign and132 = a132 & b132;
  assign or132  = a132 | b132;
  assign c133 = (a132 & b132) | (a132 & c132) | (b132 & c132);
  wire c_sub133;
  assign c_sub133 = (a132 & b_inv132) | (a132 & c132) | (b_inv132 & c132);
  wire s133, sub133, and133, or133;
  wire b_inv133;
  assign b_inv133 = ~b133;
  assign s133  = a133 ^ b133 ^ c133;
  assign sub133 = a133 ^ b_inv133 ^ c133;
  assign and133 = a133 & b133;
  assign or133  = a133 | b133;
  assign c134 = (a133 & b133) | (a133 & c133) | (b133 & c133);
  wire c_sub134;
  assign c_sub134 = (a133 & b_inv133) | (a133 & c133) | (b_inv133 & c133);
  wire s134, sub134, and134, or134;
  wire b_inv134;
  assign b_inv134 = ~b134;
  assign s134  = a134 ^ b134 ^ c134;
  assign sub134 = a134 ^ b_inv134 ^ c134;
  assign and134 = a134 & b134;
  assign or134  = a134 | b134;
  assign c135 = (a134 & b134) | (a134 & c134) | (b134 & c134);
  wire c_sub135;
  assign c_sub135 = (a134 & b_inv134) | (a134 & c134) | (b_inv134 & c134);
  wire s135, sub135, and135, or135;
  wire b_inv135;
  assign b_inv135 = ~b135;
  assign s135  = a135 ^ b135 ^ c135;
  assign sub135 = a135 ^ b_inv135 ^ c135;
  assign and135 = a135 & b135;
  assign or135  = a135 | b135;
  assign c136 = (a135 & b135) | (a135 & c135) | (b135 & c135);
  wire c_sub136;
  assign c_sub136 = (a135 & b_inv135) | (a135 & c135) | (b_inv135 & c135);
  wire s136, sub136, and136, or136;
  wire b_inv136;
  assign b_inv136 = ~b136;
  assign s136  = a136 ^ b136 ^ c136;
  assign sub136 = a136 ^ b_inv136 ^ c136;
  assign and136 = a136 & b136;
  assign or136  = a136 | b136;
  assign c137 = (a136 & b136) | (a136 & c136) | (b136 & c136);
  wire c_sub137;
  assign c_sub137 = (a136 & b_inv136) | (a136 & c136) | (b_inv136 & c136);
  wire s137, sub137, and137, or137;
  wire b_inv137;
  assign b_inv137 = ~b137;
  assign s137  = a137 ^ b137 ^ c137;
  assign sub137 = a137 ^ b_inv137 ^ c137;
  assign and137 = a137 & b137;
  assign or137  = a137 | b137;
  assign c138 = (a137 & b137) | (a137 & c137) | (b137 & c137);
  wire c_sub138;
  assign c_sub138 = (a137 & b_inv137) | (a137 & c137) | (b_inv137 & c137);
  wire s138, sub138, and138, or138;
  wire b_inv138;
  assign b_inv138 = ~b138;
  assign s138  = a138 ^ b138 ^ c138;
  assign sub138 = a138 ^ b_inv138 ^ c138;
  assign and138 = a138 & b138;
  assign or138  = a138 | b138;
  assign c139 = (a138 & b138) | (a138 & c138) | (b138 & c138);
  wire c_sub139;
  assign c_sub139 = (a138 & b_inv138) | (a138 & c138) | (b_inv138 & c138);
  wire s139, sub139, and139, or139;
  wire b_inv139;
  assign b_inv139 = ~b139;
  assign s139  = a139 ^ b139 ^ c139;
  assign sub139 = a139 ^ b_inv139 ^ c139;
  assign and139 = a139 & b139;
  assign or139  = a139 | b139;
  assign c140 = (a139 & b139) | (a139 & c139) | (b139 & c139);
  wire c_sub140;
  assign c_sub140 = (a139 & b_inv139) | (a139 & c139) | (b_inv139 & c139);
  wire s140, sub140, and140, or140;
  wire b_inv140;
  assign b_inv140 = ~b140;
  assign s140  = a140 ^ b140 ^ c140;
  assign sub140 = a140 ^ b_inv140 ^ c140;
  assign and140 = a140 & b140;
  assign or140  = a140 | b140;
  assign c141 = (a140 & b140) | (a140 & c140) | (b140 & c140);
  wire c_sub141;
  assign c_sub141 = (a140 & b_inv140) | (a140 & c140) | (b_inv140 & c140);
  wire s141, sub141, and141, or141;
  wire b_inv141;
  assign b_inv141 = ~b141;
  assign s141  = a141 ^ b141 ^ c141;
  assign sub141 = a141 ^ b_inv141 ^ c141;
  assign and141 = a141 & b141;
  assign or141  = a141 | b141;
  assign c142 = (a141 & b141) | (a141 & c141) | (b141 & c141);
  wire c_sub142;
  assign c_sub142 = (a141 & b_inv141) | (a141 & c141) | (b_inv141 & c141);
  wire s142, sub142, and142, or142;
  wire b_inv142;
  assign b_inv142 = ~b142;
  assign s142  = a142 ^ b142 ^ c142;
  assign sub142 = a142 ^ b_inv142 ^ c142;
  assign and142 = a142 & b142;
  assign or142  = a142 | b142;
  assign c143 = (a142 & b142) | (a142 & c142) | (b142 & c142);
  wire c_sub143;
  assign c_sub143 = (a142 & b_inv142) | (a142 & c142) | (b_inv142 & c142);
  wire s143, sub143, and143, or143;
  wire b_inv143;
  assign b_inv143 = ~b143;
  assign s143  = a143 ^ b143 ^ c143;
  assign sub143 = a143 ^ b_inv143 ^ c143;
  assign and143 = a143 & b143;
  assign or143  = a143 | b143;
  assign c144 = (a143 & b143) | (a143 & c143) | (b143 & c143);
  wire c_sub144;
  assign c_sub144 = (a143 & b_inv143) | (a143 & c143) | (b_inv143 & c143);
  wire s144, sub144, and144, or144;
  wire b_inv144;
  assign b_inv144 = ~b144;
  assign s144  = a144 ^ b144 ^ c144;
  assign sub144 = a144 ^ b_inv144 ^ c144;
  assign and144 = a144 & b144;
  assign or144  = a144 | b144;
  assign c145 = (a144 & b144) | (a144 & c144) | (b144 & c144);
  wire c_sub145;
  assign c_sub145 = (a144 & b_inv144) | (a144 & c144) | (b_inv144 & c144);
  wire s145, sub145, and145, or145;
  wire b_inv145;
  assign b_inv145 = ~b145;
  assign s145  = a145 ^ b145 ^ c145;
  assign sub145 = a145 ^ b_inv145 ^ c145;
  assign and145 = a145 & b145;
  assign or145  = a145 | b145;
  assign c146 = (a145 & b145) | (a145 & c145) | (b145 & c145);
  wire c_sub146;
  assign c_sub146 = (a145 & b_inv145) | (a145 & c145) | (b_inv145 & c145);
  wire s146, sub146, and146, or146;
  wire b_inv146;
  assign b_inv146 = ~b146;
  assign s146  = a146 ^ b146 ^ c146;
  assign sub146 = a146 ^ b_inv146 ^ c146;
  assign and146 = a146 & b146;
  assign or146  = a146 | b146;
  assign c147 = (a146 & b146) | (a146 & c146) | (b146 & c146);
  wire c_sub147;
  assign c_sub147 = (a146 & b_inv146) | (a146 & c146) | (b_inv146 & c146);
  wire s147, sub147, and147, or147;
  wire b_inv147;
  assign b_inv147 = ~b147;
  assign s147  = a147 ^ b147 ^ c147;
  assign sub147 = a147 ^ b_inv147 ^ c147;
  assign and147 = a147 & b147;
  assign or147  = a147 | b147;
  assign c148 = (a147 & b147) | (a147 & c147) | (b147 & c147);
  wire c_sub148;
  assign c_sub148 = (a147 & b_inv147) | (a147 & c147) | (b_inv147 & c147);
  wire s148, sub148, and148, or148;
  wire b_inv148;
  assign b_inv148 = ~b148;
  assign s148  = a148 ^ b148 ^ c148;
  assign sub148 = a148 ^ b_inv148 ^ c148;
  assign and148 = a148 & b148;
  assign or148  = a148 | b148;
  assign c149 = (a148 & b148) | (a148 & c148) | (b148 & c148);
  wire c_sub149;
  assign c_sub149 = (a148 & b_inv148) | (a148 & c148) | (b_inv148 & c148);
  wire s149, sub149, and149, or149;
  wire b_inv149;
  assign b_inv149 = ~b149;
  assign s149  = a149 ^ b149 ^ c149;
  assign sub149 = a149 ^ b_inv149 ^ c149;
  assign and149 = a149 & b149;
  assign or149  = a149 | b149;
  assign c150 = (a149 & b149) | (a149 & c149) | (b149 & c149);
  wire c_sub150;
  assign c_sub150 = (a149 & b_inv149) | (a149 & c149) | (b_inv149 & c149);
  wire s150, sub150, and150, or150;
  wire b_inv150;
  assign b_inv150 = ~b150;
  assign s150  = a150 ^ b150 ^ c150;
  assign sub150 = a150 ^ b_inv150 ^ c150;
  assign and150 = a150 & b150;
  assign or150  = a150 | b150;
  assign c151 = (a150 & b150) | (a150 & c150) | (b150 & c150);
  wire c_sub151;
  assign c_sub151 = (a150 & b_inv150) | (a150 & c150) | (b_inv150 & c150);
  wire s151, sub151, and151, or151;
  wire b_inv151;
  assign b_inv151 = ~b151;
  assign s151  = a151 ^ b151 ^ c151;
  assign sub151 = a151 ^ b_inv151 ^ c151;
  assign and151 = a151 & b151;
  assign or151  = a151 | b151;
  assign c152 = (a151 & b151) | (a151 & c151) | (b151 & c151);
  wire c_sub152;
  assign c_sub152 = (a151 & b_inv151) | (a151 & c151) | (b_inv151 & c151);
  wire s152, sub152, and152, or152;
  wire b_inv152;
  assign b_inv152 = ~b152;
  assign s152  = a152 ^ b152 ^ c152;
  assign sub152 = a152 ^ b_inv152 ^ c152;
  assign and152 = a152 & b152;
  assign or152  = a152 | b152;
  assign c153 = (a152 & b152) | (a152 & c152) | (b152 & c152);
  wire c_sub153;
  assign c_sub153 = (a152 & b_inv152) | (a152 & c152) | (b_inv152 & c152);
  wire s153, sub153, and153, or153;
  wire b_inv153;
  assign b_inv153 = ~b153;
  assign s153  = a153 ^ b153 ^ c153;
  assign sub153 = a153 ^ b_inv153 ^ c153;
  assign and153 = a153 & b153;
  assign or153  = a153 | b153;
  assign c154 = (a153 & b153) | (a153 & c153) | (b153 & c153);
  wire c_sub154;
  assign c_sub154 = (a153 & b_inv153) | (a153 & c153) | (b_inv153 & c153);
  wire s154, sub154, and154, or154;
  wire b_inv154;
  assign b_inv154 = ~b154;
  assign s154  = a154 ^ b154 ^ c154;
  assign sub154 = a154 ^ b_inv154 ^ c154;
  assign and154 = a154 & b154;
  assign or154  = a154 | b154;
  assign c155 = (a154 & b154) | (a154 & c154) | (b154 & c154);
  wire c_sub155;
  assign c_sub155 = (a154 & b_inv154) | (a154 & c154) | (b_inv154 & c154);
  wire s155, sub155, and155, or155;
  wire b_inv155;
  assign b_inv155 = ~b155;
  assign s155  = a155 ^ b155 ^ c155;
  assign sub155 = a155 ^ b_inv155 ^ c155;
  assign and155 = a155 & b155;
  assign or155  = a155 | b155;
  assign c156 = (a155 & b155) | (a155 & c155) | (b155 & c155);
  wire c_sub156;
  assign c_sub156 = (a155 & b_inv155) | (a155 & c155) | (b_inv155 & c155);
  wire s156, sub156, and156, or156;
  wire b_inv156;
  assign b_inv156 = ~b156;
  assign s156  = a156 ^ b156 ^ c156;
  assign sub156 = a156 ^ b_inv156 ^ c156;
  assign and156 = a156 & b156;
  assign or156  = a156 | b156;
  assign c157 = (a156 & b156) | (a156 & c156) | (b156 & c156);
  wire c_sub157;
  assign c_sub157 = (a156 & b_inv156) | (a156 & c156) | (b_inv156 & c156);
  wire s157, sub157, and157, or157;
  wire b_inv157;
  assign b_inv157 = ~b157;
  assign s157  = a157 ^ b157 ^ c157;
  assign sub157 = a157 ^ b_inv157 ^ c157;
  assign and157 = a157 & b157;
  assign or157  = a157 | b157;
  assign c158 = (a157 & b157) | (a157 & c157) | (b157 & c157);
  wire c_sub158;
  assign c_sub158 = (a157 & b_inv157) | (a157 & c157) | (b_inv157 & c157);
  wire s158, sub158, and158, or158;
  wire b_inv158;
  assign b_inv158 = ~b158;
  assign s158  = a158 ^ b158 ^ c158;
  assign sub158 = a158 ^ b_inv158 ^ c158;
  assign and158 = a158 & b158;
  assign or158  = a158 | b158;
  assign c159 = (a158 & b158) | (a158 & c158) | (b158 & c158);
  wire c_sub159;
  assign c_sub159 = (a158 & b_inv158) | (a158 & c158) | (b_inv158 & c158);
  wire s159, sub159, and159, or159;
  wire b_inv159;
  assign b_inv159 = ~b159;
  assign s159  = a159 ^ b159 ^ c159;
  assign sub159 = a159 ^ b_inv159 ^ c159;
  assign and159 = a159 & b159;
  assign or159  = a159 | b159;
  assign c160 = (a159 & b159) | (a159 & c159) | (b159 & c159);
  wire c_sub160;
  assign c_sub160 = (a159 & b_inv159) | (a159 & c159) | (b_inv159 & c159);
  wire s160, sub160, and160, or160;
  wire b_inv160;
  assign b_inv160 = ~b160;
  assign s160  = a160 ^ b160 ^ c160;
  assign sub160 = a160 ^ b_inv160 ^ c160;
  assign and160 = a160 & b160;
  assign or160  = a160 | b160;
  assign c161 = (a160 & b160) | (a160 & c160) | (b160 & c160);
  wire c_sub161;
  assign c_sub161 = (a160 & b_inv160) | (a160 & c160) | (b_inv160 & c160);
  wire s161, sub161, and161, or161;
  wire b_inv161;
  assign b_inv161 = ~b161;
  assign s161  = a161 ^ b161 ^ c161;
  assign sub161 = a161 ^ b_inv161 ^ c161;
  assign and161 = a161 & b161;
  assign or161  = a161 | b161;
  assign c162 = (a161 & b161) | (a161 & c161) | (b161 & c161);
  wire c_sub162;
  assign c_sub162 = (a161 & b_inv161) | (a161 & c161) | (b_inv161 & c161);
  wire s162, sub162, and162, or162;
  wire b_inv162;
  assign b_inv162 = ~b162;
  assign s162  = a162 ^ b162 ^ c162;
  assign sub162 = a162 ^ b_inv162 ^ c162;
  assign and162 = a162 & b162;
  assign or162  = a162 | b162;
  assign c163 = (a162 & b162) | (a162 & c162) | (b162 & c162);
  wire c_sub163;
  assign c_sub163 = (a162 & b_inv162) | (a162 & c162) | (b_inv162 & c162);
  wire s163, sub163, and163, or163;
  wire b_inv163;
  assign b_inv163 = ~b163;
  assign s163  = a163 ^ b163 ^ c163;
  assign sub163 = a163 ^ b_inv163 ^ c163;
  assign and163 = a163 & b163;
  assign or163  = a163 | b163;
  assign c164 = (a163 & b163) | (a163 & c163) | (b163 & c163);
  wire c_sub164;
  assign c_sub164 = (a163 & b_inv163) | (a163 & c163) | (b_inv163 & c163);
  wire s164, sub164, and164, or164;
  wire b_inv164;
  assign b_inv164 = ~b164;
  assign s164  = a164 ^ b164 ^ c164;
  assign sub164 = a164 ^ b_inv164 ^ c164;
  assign and164 = a164 & b164;
  assign or164  = a164 | b164;
  assign c165 = (a164 & b164) | (a164 & c164) | (b164 & c164);
  wire c_sub165;
  assign c_sub165 = (a164 & b_inv164) | (a164 & c164) | (b_inv164 & c164);
  wire s165, sub165, and165, or165;
  wire b_inv165;
  assign b_inv165 = ~b165;
  assign s165  = a165 ^ b165 ^ c165;
  assign sub165 = a165 ^ b_inv165 ^ c165;
  assign and165 = a165 & b165;
  assign or165  = a165 | b165;
  assign c166 = (a165 & b165) | (a165 & c165) | (b165 & c165);
  wire c_sub166;
  assign c_sub166 = (a165 & b_inv165) | (a165 & c165) | (b_inv165 & c165);
  wire s166, sub166, and166, or166;
  wire b_inv166;
  assign b_inv166 = ~b166;
  assign s166  = a166 ^ b166 ^ c166;
  assign sub166 = a166 ^ b_inv166 ^ c166;
  assign and166 = a166 & b166;
  assign or166  = a166 | b166;
  assign c167 = (a166 & b166) | (a166 & c166) | (b166 & c166);
  wire c_sub167;
  assign c_sub167 = (a166 & b_inv166) | (a166 & c166) | (b_inv166 & c166);
  wire s167, sub167, and167, or167;
  wire b_inv167;
  assign b_inv167 = ~b167;
  assign s167  = a167 ^ b167 ^ c167;
  assign sub167 = a167 ^ b_inv167 ^ c167;
  assign and167 = a167 & b167;
  assign or167  = a167 | b167;
  assign c168 = (a167 & b167) | (a167 & c167) | (b167 & c167);
  wire c_sub168;
  assign c_sub168 = (a167 & b_inv167) | (a167 & c167) | (b_inv167 & c167);
  wire s168, sub168, and168, or168;
  wire b_inv168;
  assign b_inv168 = ~b168;
  assign s168  = a168 ^ b168 ^ c168;
  assign sub168 = a168 ^ b_inv168 ^ c168;
  assign and168 = a168 & b168;
  assign or168  = a168 | b168;
  assign c169 = (a168 & b168) | (a168 & c168) | (b168 & c168);
  wire c_sub169;
  assign c_sub169 = (a168 & b_inv168) | (a168 & c168) | (b_inv168 & c168);
  wire s169, sub169, and169, or169;
  wire b_inv169;
  assign b_inv169 = ~b169;
  assign s169  = a169 ^ b169 ^ c169;
  assign sub169 = a169 ^ b_inv169 ^ c169;
  assign and169 = a169 & b169;
  assign or169  = a169 | b169;
  assign c170 = (a169 & b169) | (a169 & c169) | (b169 & c169);
  wire c_sub170;
  assign c_sub170 = (a169 & b_inv169) | (a169 & c169) | (b_inv169 & c169);
  wire s170, sub170, and170, or170;
  wire b_inv170;
  assign b_inv170 = ~b170;
  assign s170  = a170 ^ b170 ^ c170;
  assign sub170 = a170 ^ b_inv170 ^ c170;
  assign and170 = a170 & b170;
  assign or170  = a170 | b170;
  assign c171 = (a170 & b170) | (a170 & c170) | (b170 & c170);
  wire c_sub171;
  assign c_sub171 = (a170 & b_inv170) | (a170 & c170) | (b_inv170 & c170);
  wire s171, sub171, and171, or171;
  wire b_inv171;
  assign b_inv171 = ~b171;
  assign s171  = a171 ^ b171 ^ c171;
  assign sub171 = a171 ^ b_inv171 ^ c171;
  assign and171 = a171 & b171;
  assign or171  = a171 | b171;
  assign c172 = (a171 & b171) | (a171 & c171) | (b171 & c171);
  wire c_sub172;
  assign c_sub172 = (a171 & b_inv171) | (a171 & c171) | (b_inv171 & c171);
  wire s172, sub172, and172, or172;
  wire b_inv172;
  assign b_inv172 = ~b172;
  assign s172  = a172 ^ b172 ^ c172;
  assign sub172 = a172 ^ b_inv172 ^ c172;
  assign and172 = a172 & b172;
  assign or172  = a172 | b172;
  assign c173 = (a172 & b172) | (a172 & c172) | (b172 & c172);
  wire c_sub173;
  assign c_sub173 = (a172 & b_inv172) | (a172 & c172) | (b_inv172 & c172);
  wire s173, sub173, and173, or173;
  wire b_inv173;
  assign b_inv173 = ~b173;
  assign s173  = a173 ^ b173 ^ c173;
  assign sub173 = a173 ^ b_inv173 ^ c173;
  assign and173 = a173 & b173;
  assign or173  = a173 | b173;
  assign c174 = (a173 & b173) | (a173 & c173) | (b173 & c173);
  wire c_sub174;
  assign c_sub174 = (a173 & b_inv173) | (a173 & c173) | (b_inv173 & c173);
  wire s174, sub174, and174, or174;
  wire b_inv174;
  assign b_inv174 = ~b174;
  assign s174  = a174 ^ b174 ^ c174;
  assign sub174 = a174 ^ b_inv174 ^ c174;
  assign and174 = a174 & b174;
  assign or174  = a174 | b174;
  assign c175 = (a174 & b174) | (a174 & c174) | (b174 & c174);
  wire c_sub175;
  assign c_sub175 = (a174 & b_inv174) | (a174 & c174) | (b_inv174 & c174);
  wire s175, sub175, and175, or175;
  wire b_inv175;
  assign b_inv175 = ~b175;
  assign s175  = a175 ^ b175 ^ c175;
  assign sub175 = a175 ^ b_inv175 ^ c175;
  assign and175 = a175 & b175;
  assign or175  = a175 | b175;
  assign c176 = (a175 & b175) | (a175 & c175) | (b175 & c175);
  wire c_sub176;
  assign c_sub176 = (a175 & b_inv175) | (a175 & c175) | (b_inv175 & c175);
  wire s176, sub176, and176, or176;
  wire b_inv176;
  assign b_inv176 = ~b176;
  assign s176  = a176 ^ b176 ^ c176;
  assign sub176 = a176 ^ b_inv176 ^ c176;
  assign and176 = a176 & b176;
  assign or176  = a176 | b176;
  assign c177 = (a176 & b176) | (a176 & c176) | (b176 & c176);
  wire c_sub177;
  assign c_sub177 = (a176 & b_inv176) | (a176 & c176) | (b_inv176 & c176);
  wire s177, sub177, and177, or177;
  wire b_inv177;
  assign b_inv177 = ~b177;
  assign s177  = a177 ^ b177 ^ c177;
  assign sub177 = a177 ^ b_inv177 ^ c177;
  assign and177 = a177 & b177;
  assign or177  = a177 | b177;
  assign c178 = (a177 & b177) | (a177 & c177) | (b177 & c177);
  wire c_sub178;
  assign c_sub178 = (a177 & b_inv177) | (a177 & c177) | (b_inv177 & c177);
  wire s178, sub178, and178, or178;
  wire b_inv178;
  assign b_inv178 = ~b178;
  assign s178  = a178 ^ b178 ^ c178;
  assign sub178 = a178 ^ b_inv178 ^ c178;
  assign and178 = a178 & b178;
  assign or178  = a178 | b178;
  assign c179 = (a178 & b178) | (a178 & c178) | (b178 & c178);
  wire c_sub179;
  assign c_sub179 = (a178 & b_inv178) | (a178 & c178) | (b_inv178 & c178);
  wire s179, sub179, and179, or179;
  wire b_inv179;
  assign b_inv179 = ~b179;
  assign s179  = a179 ^ b179 ^ c179;
  assign sub179 = a179 ^ b_inv179 ^ c179;
  assign and179 = a179 & b179;
  assign or179  = a179 | b179;
  assign c180 = (a179 & b179) | (a179 & c179) | (b179 & c179);
  wire c_sub180;
  assign c_sub180 = (a179 & b_inv179) | (a179 & c179) | (b_inv179 & c179);
  wire s180, sub180, and180, or180;
  wire b_inv180;
  assign b_inv180 = ~b180;
  assign s180  = a180 ^ b180 ^ c180;
  assign sub180 = a180 ^ b_inv180 ^ c180;
  assign and180 = a180 & b180;
  assign or180  = a180 | b180;
  assign c181 = (a180 & b180) | (a180 & c180) | (b180 & c180);
  wire c_sub181;
  assign c_sub181 = (a180 & b_inv180) | (a180 & c180) | (b_inv180 & c180);
  wire s181, sub181, and181, or181;
  wire b_inv181;
  assign b_inv181 = ~b181;
  assign s181  = a181 ^ b181 ^ c181;
  assign sub181 = a181 ^ b_inv181 ^ c181;
  assign and181 = a181 & b181;
  assign or181  = a181 | b181;
  assign c182 = (a181 & b181) | (a181 & c181) | (b181 & c181);
  wire c_sub182;
  assign c_sub182 = (a181 & b_inv181) | (a181 & c181) | (b_inv181 & c181);
  wire s182, sub182, and182, or182;
  wire b_inv182;
  assign b_inv182 = ~b182;
  assign s182  = a182 ^ b182 ^ c182;
  assign sub182 = a182 ^ b_inv182 ^ c182;
  assign and182 = a182 & b182;
  assign or182  = a182 | b182;
  assign c183 = (a182 & b182) | (a182 & c182) | (b182 & c182);
  wire c_sub183;
  assign c_sub183 = (a182 & b_inv182) | (a182 & c182) | (b_inv182 & c182);
  wire s183, sub183, and183, or183;
  wire b_inv183;
  assign b_inv183 = ~b183;
  assign s183  = a183 ^ b183 ^ c183;
  assign sub183 = a183 ^ b_inv183 ^ c183;
  assign and183 = a183 & b183;
  assign or183  = a183 | b183;
  assign c184 = (a183 & b183) | (a183 & c183) | (b183 & c183);
  wire c_sub184;
  assign c_sub184 = (a183 & b_inv183) | (a183 & c183) | (b_inv183 & c183);
  wire s184, sub184, and184, or184;
  wire b_inv184;
  assign b_inv184 = ~b184;
  assign s184  = a184 ^ b184 ^ c184;
  assign sub184 = a184 ^ b_inv184 ^ c184;
  assign and184 = a184 & b184;
  assign or184  = a184 | b184;
  assign c185 = (a184 & b184) | (a184 & c184) | (b184 & c184);
  wire c_sub185;
  assign c_sub185 = (a184 & b_inv184) | (a184 & c184) | (b_inv184 & c184);
  wire s185, sub185, and185, or185;
  wire b_inv185;
  assign b_inv185 = ~b185;
  assign s185  = a185 ^ b185 ^ c185;
  assign sub185 = a185 ^ b_inv185 ^ c185;
  assign and185 = a185 & b185;
  assign or185  = a185 | b185;
  assign c186 = (a185 & b185) | (a185 & c185) | (b185 & c185);
  wire c_sub186;
  assign c_sub186 = (a185 & b_inv185) | (a185 & c185) | (b_inv185 & c185);
  wire s186, sub186, and186, or186;
  wire b_inv186;
  assign b_inv186 = ~b186;
  assign s186  = a186 ^ b186 ^ c186;
  assign sub186 = a186 ^ b_inv186 ^ c186;
  assign and186 = a186 & b186;
  assign or186  = a186 | b186;
  assign c187 = (a186 & b186) | (a186 & c186) | (b186 & c186);
  wire c_sub187;
  assign c_sub187 = (a186 & b_inv186) | (a186 & c186) | (b_inv186 & c186);
  wire s187, sub187, and187, or187;
  wire b_inv187;
  assign b_inv187 = ~b187;
  assign s187  = a187 ^ b187 ^ c187;
  assign sub187 = a187 ^ b_inv187 ^ c187;
  assign and187 = a187 & b187;
  assign or187  = a187 | b187;
  assign c188 = (a187 & b187) | (a187 & c187) | (b187 & c187);
  wire c_sub188;
  assign c_sub188 = (a187 & b_inv187) | (a187 & c187) | (b_inv187 & c187);
  wire s188, sub188, and188, or188;
  wire b_inv188;
  assign b_inv188 = ~b188;
  assign s188  = a188 ^ b188 ^ c188;
  assign sub188 = a188 ^ b_inv188 ^ c188;
  assign and188 = a188 & b188;
  assign or188  = a188 | b188;
  assign c189 = (a188 & b188) | (a188 & c188) | (b188 & c188);
  wire c_sub189;
  assign c_sub189 = (a188 & b_inv188) | (a188 & c188) | (b_inv188 & c188);
  wire s189, sub189, and189, or189;
  wire b_inv189;
  assign b_inv189 = ~b189;
  assign s189  = a189 ^ b189 ^ c189;
  assign sub189 = a189 ^ b_inv189 ^ c189;
  assign and189 = a189 & b189;
  assign or189  = a189 | b189;
  assign c190 = (a189 & b189) | (a189 & c189) | (b189 & c189);
  wire c_sub190;
  assign c_sub190 = (a189 & b_inv189) | (a189 & c189) | (b_inv189 & c189);
  wire s190, sub190, and190, or190;
  wire b_inv190;
  assign b_inv190 = ~b190;
  assign s190  = a190 ^ b190 ^ c190;
  assign sub190 = a190 ^ b_inv190 ^ c190;
  assign and190 = a190 & b190;
  assign or190  = a190 | b190;
  assign c191 = (a190 & b190) | (a190 & c190) | (b190 & c190);
  wire c_sub191;
  assign c_sub191 = (a190 & b_inv190) | (a190 & c190) | (b_inv190 & c190);
  wire s191, sub191, and191, or191;
  wire b_inv191;
  assign b_inv191 = ~b191;
  assign s191  = a191 ^ b191 ^ c191;
  assign sub191 = a191 ^ b_inv191 ^ c191;
  assign and191 = a191 & b191;
  assign or191  = a191 | b191;
  assign c192 = (a191 & b191) | (a191 & c191) | (b191 & c191);
  wire c_sub192;
  assign c_sub192 = (a191 & b_inv191) | (a191 & c191) | (b_inv191 & c191);
  wire s192, sub192, and192, or192;
  wire b_inv192;
  assign b_inv192 = ~b192;
  assign s192  = a192 ^ b192 ^ c192;
  assign sub192 = a192 ^ b_inv192 ^ c192;
  assign and192 = a192 & b192;
  assign or192  = a192 | b192;
  assign c193 = (a192 & b192) | (a192 & c192) | (b192 & c192);
  wire c_sub193;
  assign c_sub193 = (a192 & b_inv192) | (a192 & c192) | (b_inv192 & c192);
  wire s193, sub193, and193, or193;
  wire b_inv193;
  assign b_inv193 = ~b193;
  assign s193  = a193 ^ b193 ^ c193;
  assign sub193 = a193 ^ b_inv193 ^ c193;
  assign and193 = a193 & b193;
  assign or193  = a193 | b193;
  assign c194 = (a193 & b193) | (a193 & c193) | (b193 & c193);
  wire c_sub194;
  assign c_sub194 = (a193 & b_inv193) | (a193 & c193) | (b_inv193 & c193);
  wire s194, sub194, and194, or194;
  wire b_inv194;
  assign b_inv194 = ~b194;
  assign s194  = a194 ^ b194 ^ c194;
  assign sub194 = a194 ^ b_inv194 ^ c194;
  assign and194 = a194 & b194;
  assign or194  = a194 | b194;
  assign c195 = (a194 & b194) | (a194 & c194) | (b194 & c194);
  wire c_sub195;
  assign c_sub195 = (a194 & b_inv194) | (a194 & c194) | (b_inv194 & c194);
  wire s195, sub195, and195, or195;
  wire b_inv195;
  assign b_inv195 = ~b195;
  assign s195  = a195 ^ b195 ^ c195;
  assign sub195 = a195 ^ b_inv195 ^ c195;
  assign and195 = a195 & b195;
  assign or195  = a195 | b195;
  assign c196 = (a195 & b195) | (a195 & c195) | (b195 & c195);
  wire c_sub196;
  assign c_sub196 = (a195 & b_inv195) | (a195 & c195) | (b_inv195 & c195);
  wire s196, sub196, and196, or196;
  wire b_inv196;
  assign b_inv196 = ~b196;
  assign s196  = a196 ^ b196 ^ c196;
  assign sub196 = a196 ^ b_inv196 ^ c196;
  assign and196 = a196 & b196;
  assign or196  = a196 | b196;
  assign c197 = (a196 & b196) | (a196 & c196) | (b196 & c196);
  wire c_sub197;
  assign c_sub197 = (a196 & b_inv196) | (a196 & c196) | (b_inv196 & c196);
  wire s197, sub197, and197, or197;
  wire b_inv197;
  assign b_inv197 = ~b197;
  assign s197  = a197 ^ b197 ^ c197;
  assign sub197 = a197 ^ b_inv197 ^ c197;
  assign and197 = a197 & b197;
  assign or197  = a197 | b197;
  assign c198 = (a197 & b197) | (a197 & c197) | (b197 & c197);
  wire c_sub198;
  assign c_sub198 = (a197 & b_inv197) | (a197 & c197) | (b_inv197 & c197);
  wire s198, sub198, and198, or198;
  wire b_inv198;
  assign b_inv198 = ~b198;
  assign s198  = a198 ^ b198 ^ c198;
  assign sub198 = a198 ^ b_inv198 ^ c198;
  assign and198 = a198 & b198;
  assign or198  = a198 | b198;
  assign c199 = (a198 & b198) | (a198 & c198) | (b198 & c198);
  wire c_sub199;
  assign c_sub199 = (a198 & b_inv198) | (a198 & c198) | (b_inv198 & c198);
  wire s199, sub199, and199, or199;
  wire b_inv199;
  assign b_inv199 = ~b199;
  assign s199  = a199 ^ b199 ^ c199;
  assign sub199 = a199 ^ b_inv199 ^ c199;
  assign and199 = a199 & b199;
  assign or199  = a199 | b199;
  assign c200 = (a199 & b199) | (a199 & c199) | (b199 & c199);
  wire c_sub200;
  assign c_sub200 = (a199 & b_inv199) | (a199 & c199) | (b_inv199 & c199);
  wire s200, sub200, and200, or200;
  wire b_inv200;
  assign b_inv200 = ~b200;
  assign s200  = a200 ^ b200 ^ c200;
  assign sub200 = a200 ^ b_inv200 ^ c200;
  assign and200 = a200 & b200;
  assign or200  = a200 | b200;
  assign c201 = (a200 & b200) | (a200 & c200) | (b200 & c200);
  wire c_sub201;
  assign c_sub201 = (a200 & b_inv200) | (a200 & c200) | (b_inv200 & c200);
  wire s201, sub201, and201, or201;
  wire b_inv201;
  assign b_inv201 = ~b201;
  assign s201  = a201 ^ b201 ^ c201;
  assign sub201 = a201 ^ b_inv201 ^ c201;
  assign and201 = a201 & b201;
  assign or201  = a201 | b201;
  assign c202 = (a201 & b201) | (a201 & c201) | (b201 & c201);
  wire c_sub202;
  assign c_sub202 = (a201 & b_inv201) | (a201 & c201) | (b_inv201 & c201);
  wire s202, sub202, and202, or202;
  wire b_inv202;
  assign b_inv202 = ~b202;
  assign s202  = a202 ^ b202 ^ c202;
  assign sub202 = a202 ^ b_inv202 ^ c202;
  assign and202 = a202 & b202;
  assign or202  = a202 | b202;
  assign c203 = (a202 & b202) | (a202 & c202) | (b202 & c202);
  wire c_sub203;
  assign c_sub203 = (a202 & b_inv202) | (a202 & c202) | (b_inv202 & c202);
  wire s203, sub203, and203, or203;
  wire b_inv203;
  assign b_inv203 = ~b203;
  assign s203  = a203 ^ b203 ^ c203;
  assign sub203 = a203 ^ b_inv203 ^ c203;
  assign and203 = a203 & b203;
  assign or203  = a203 | b203;
  assign c204 = (a203 & b203) | (a203 & c203) | (b203 & c203);
  wire c_sub204;
  assign c_sub204 = (a203 & b_inv203) | (a203 & c203) | (b_inv203 & c203);
  wire s204, sub204, and204, or204;
  wire b_inv204;
  assign b_inv204 = ~b204;
  assign s204  = a204 ^ b204 ^ c204;
  assign sub204 = a204 ^ b_inv204 ^ c204;
  assign and204 = a204 & b204;
  assign or204  = a204 | b204;
  assign c205 = (a204 & b204) | (a204 & c204) | (b204 & c204);
  wire c_sub205;
  assign c_sub205 = (a204 & b_inv204) | (a204 & c204) | (b_inv204 & c204);
  wire s205, sub205, and205, or205;
  wire b_inv205;
  assign b_inv205 = ~b205;
  assign s205  = a205 ^ b205 ^ c205;
  assign sub205 = a205 ^ b_inv205 ^ c205;
  assign and205 = a205 & b205;
  assign or205  = a205 | b205;
  assign c206 = (a205 & b205) | (a205 & c205) | (b205 & c205);
  wire c_sub206;
  assign c_sub206 = (a205 & b_inv205) | (a205 & c205) | (b_inv205 & c205);
  wire s206, sub206, and206, or206;
  wire b_inv206;
  assign b_inv206 = ~b206;
  assign s206  = a206 ^ b206 ^ c206;
  assign sub206 = a206 ^ b_inv206 ^ c206;
  assign and206 = a206 & b206;
  assign or206  = a206 | b206;
  assign c207 = (a206 & b206) | (a206 & c206) | (b206 & c206);
  wire c_sub207;
  assign c_sub207 = (a206 & b_inv206) | (a206 & c206) | (b_inv206 & c206);
  wire s207, sub207, and207, or207;
  wire b_inv207;
  assign b_inv207 = ~b207;
  assign s207  = a207 ^ b207 ^ c207;
  assign sub207 = a207 ^ b_inv207 ^ c207;
  assign and207 = a207 & b207;
  assign or207  = a207 | b207;
  assign c208 = (a207 & b207) | (a207 & c207) | (b207 & c207);
  wire c_sub208;
  assign c_sub208 = (a207 & b_inv207) | (a207 & c207) | (b_inv207 & c207);
  wire s208, sub208, and208, or208;
  wire b_inv208;
  assign b_inv208 = ~b208;
  assign s208  = a208 ^ b208 ^ c208;
  assign sub208 = a208 ^ b_inv208 ^ c208;
  assign and208 = a208 & b208;
  assign or208  = a208 | b208;
  assign c209 = (a208 & b208) | (a208 & c208) | (b208 & c208);
  wire c_sub209;
  assign c_sub209 = (a208 & b_inv208) | (a208 & c208) | (b_inv208 & c208);
  wire s209, sub209, and209, or209;
  wire b_inv209;
  assign b_inv209 = ~b209;
  assign s209  = a209 ^ b209 ^ c209;
  assign sub209 = a209 ^ b_inv209 ^ c209;
  assign and209 = a209 & b209;
  assign or209  = a209 | b209;
  assign c210 = (a209 & b209) | (a209 & c209) | (b209 & c209);
  wire c_sub210;
  assign c_sub210 = (a209 & b_inv209) | (a209 & c209) | (b_inv209 & c209);
  wire s210, sub210, and210, or210;
  wire b_inv210;
  assign b_inv210 = ~b210;
  assign s210  = a210 ^ b210 ^ c210;
  assign sub210 = a210 ^ b_inv210 ^ c210;
  assign and210 = a210 & b210;
  assign or210  = a210 | b210;
  assign c211 = (a210 & b210) | (a210 & c210) | (b210 & c210);
  wire c_sub211;
  assign c_sub211 = (a210 & b_inv210) | (a210 & c210) | (b_inv210 & c210);
  wire s211, sub211, and211, or211;
  wire b_inv211;
  assign b_inv211 = ~b211;
  assign s211  = a211 ^ b211 ^ c211;
  assign sub211 = a211 ^ b_inv211 ^ c211;
  assign and211 = a211 & b211;
  assign or211  = a211 | b211;
  assign c212 = (a211 & b211) | (a211 & c211) | (b211 & c211);
  wire c_sub212;
  assign c_sub212 = (a211 & b_inv211) | (a211 & c211) | (b_inv211 & c211);
  wire s212, sub212, and212, or212;
  wire b_inv212;
  assign b_inv212 = ~b212;
  assign s212  = a212 ^ b212 ^ c212;
  assign sub212 = a212 ^ b_inv212 ^ c212;
  assign and212 = a212 & b212;
  assign or212  = a212 | b212;
  assign c213 = (a212 & b212) | (a212 & c212) | (b212 & c212);
  wire c_sub213;
  assign c_sub213 = (a212 & b_inv212) | (a212 & c212) | (b_inv212 & c212);
  wire s213, sub213, and213, or213;
  wire b_inv213;
  assign b_inv213 = ~b213;
  assign s213  = a213 ^ b213 ^ c213;
  assign sub213 = a213 ^ b_inv213 ^ c213;
  assign and213 = a213 & b213;
  assign or213  = a213 | b213;
  assign c214 = (a213 & b213) | (a213 & c213) | (b213 & c213);
  wire c_sub214;
  assign c_sub214 = (a213 & b_inv213) | (a213 & c213) | (b_inv213 & c213);
  wire s214, sub214, and214, or214;
  wire b_inv214;
  assign b_inv214 = ~b214;
  assign s214  = a214 ^ b214 ^ c214;
  assign sub214 = a214 ^ b_inv214 ^ c214;
  assign and214 = a214 & b214;
  assign or214  = a214 | b214;
  assign c215 = (a214 & b214) | (a214 & c214) | (b214 & c214);
  wire c_sub215;
  assign c_sub215 = (a214 & b_inv214) | (a214 & c214) | (b_inv214 & c214);
  wire s215, sub215, and215, or215;
  wire b_inv215;
  assign b_inv215 = ~b215;
  assign s215  = a215 ^ b215 ^ c215;
  assign sub215 = a215 ^ b_inv215 ^ c215;
  assign and215 = a215 & b215;
  assign or215  = a215 | b215;
  assign c216 = (a215 & b215) | (a215 & c215) | (b215 & c215);
  wire c_sub216;
  assign c_sub216 = (a215 & b_inv215) | (a215 & c215) | (b_inv215 & c215);
  wire s216, sub216, and216, or216;
  wire b_inv216;
  assign b_inv216 = ~b216;
  assign s216  = a216 ^ b216 ^ c216;
  assign sub216 = a216 ^ b_inv216 ^ c216;
  assign and216 = a216 & b216;
  assign or216  = a216 | b216;
  assign c217 = (a216 & b216) | (a216 & c216) | (b216 & c216);
  wire c_sub217;
  assign c_sub217 = (a216 & b_inv216) | (a216 & c216) | (b_inv216 & c216);
  wire s217, sub217, and217, or217;
  wire b_inv217;
  assign b_inv217 = ~b217;
  assign s217  = a217 ^ b217 ^ c217;
  assign sub217 = a217 ^ b_inv217 ^ c217;
  assign and217 = a217 & b217;
  assign or217  = a217 | b217;
  assign c218 = (a217 & b217) | (a217 & c217) | (b217 & c217);
  wire c_sub218;
  assign c_sub218 = (a217 & b_inv217) | (a217 & c217) | (b_inv217 & c217);
  wire s218, sub218, and218, or218;
  wire b_inv218;
  assign b_inv218 = ~b218;
  assign s218  = a218 ^ b218 ^ c218;
  assign sub218 = a218 ^ b_inv218 ^ c218;
  assign and218 = a218 & b218;
  assign or218  = a218 | b218;
  assign c219 = (a218 & b218) | (a218 & c218) | (b218 & c218);
  wire c_sub219;
  assign c_sub219 = (a218 & b_inv218) | (a218 & c218) | (b_inv218 & c218);
  wire s219, sub219, and219, or219;
  wire b_inv219;
  assign b_inv219 = ~b219;
  assign s219  = a219 ^ b219 ^ c219;
  assign sub219 = a219 ^ b_inv219 ^ c219;
  assign and219 = a219 & b219;
  assign or219  = a219 | b219;
  assign c220 = (a219 & b219) | (a219 & c219) | (b219 & c219);
  wire c_sub220;
  assign c_sub220 = (a219 & b_inv219) | (a219 & c219) | (b_inv219 & c219);
  wire s220, sub220, and220, or220;
  wire b_inv220;
  assign b_inv220 = ~b220;
  assign s220  = a220 ^ b220 ^ c220;
  assign sub220 = a220 ^ b_inv220 ^ c220;
  assign and220 = a220 & b220;
  assign or220  = a220 | b220;
  assign c221 = (a220 & b220) | (a220 & c220) | (b220 & c220);
  wire c_sub221;
  assign c_sub221 = (a220 & b_inv220) | (a220 & c220) | (b_inv220 & c220);
  wire s221, sub221, and221, or221;
  wire b_inv221;
  assign b_inv221 = ~b221;
  assign s221  = a221 ^ b221 ^ c221;
  assign sub221 = a221 ^ b_inv221 ^ c221;
  assign and221 = a221 & b221;
  assign or221  = a221 | b221;
  assign c222 = (a221 & b221) | (a221 & c221) | (b221 & c221);
  wire c_sub222;
  assign c_sub222 = (a221 & b_inv221) | (a221 & c221) | (b_inv221 & c221);
  wire s222, sub222, and222, or222;
  wire b_inv222;
  assign b_inv222 = ~b222;
  assign s222  = a222 ^ b222 ^ c222;
  assign sub222 = a222 ^ b_inv222 ^ c222;
  assign and222 = a222 & b222;
  assign or222  = a222 | b222;
  assign c223 = (a222 & b222) | (a222 & c222) | (b222 & c222);
  wire c_sub223;
  assign c_sub223 = (a222 & b_inv222) | (a222 & c222) | (b_inv222 & c222);
  wire s223, sub223, and223, or223;
  wire b_inv223;
  assign b_inv223 = ~b223;
  assign s223  = a223 ^ b223 ^ c223;
  assign sub223 = a223 ^ b_inv223 ^ c223;
  assign and223 = a223 & b223;
  assign or223  = a223 | b223;
  assign c224 = (a223 & b223) | (a223 & c223) | (b223 & c223);
  wire c_sub224;
  assign c_sub224 = (a223 & b_inv223) | (a223 & c223) | (b_inv223 & c223);
  wire s224, sub224, and224, or224;
  wire b_inv224;
  assign b_inv224 = ~b224;
  assign s224  = a224 ^ b224 ^ c224;
  assign sub224 = a224 ^ b_inv224 ^ c224;
  assign and224 = a224 & b224;
  assign or224  = a224 | b224;
  assign c225 = (a224 & b224) | (a224 & c224) | (b224 & c224);
  wire c_sub225;
  assign c_sub225 = (a224 & b_inv224) | (a224 & c224) | (b_inv224 & c224);
  wire s225, sub225, and225, or225;
  wire b_inv225;
  assign b_inv225 = ~b225;
  assign s225  = a225 ^ b225 ^ c225;
  assign sub225 = a225 ^ b_inv225 ^ c225;
  assign and225 = a225 & b225;
  assign or225  = a225 | b225;
  assign c226 = (a225 & b225) | (a225 & c225) | (b225 & c225);
  wire c_sub226;
  assign c_sub226 = (a225 & b_inv225) | (a225 & c225) | (b_inv225 & c225);
  wire s226, sub226, and226, or226;
  wire b_inv226;
  assign b_inv226 = ~b226;
  assign s226  = a226 ^ b226 ^ c226;
  assign sub226 = a226 ^ b_inv226 ^ c226;
  assign and226 = a226 & b226;
  assign or226  = a226 | b226;
  assign c227 = (a226 & b226) | (a226 & c226) | (b226 & c226);
  wire c_sub227;
  assign c_sub227 = (a226 & b_inv226) | (a226 & c226) | (b_inv226 & c226);
  wire s227, sub227, and227, or227;
  wire b_inv227;
  assign b_inv227 = ~b227;
  assign s227  = a227 ^ b227 ^ c227;
  assign sub227 = a227 ^ b_inv227 ^ c227;
  assign and227 = a227 & b227;
  assign or227  = a227 | b227;
  assign c228 = (a227 & b227) | (a227 & c227) | (b227 & c227);
  wire c_sub228;
  assign c_sub228 = (a227 & b_inv227) | (a227 & c227) | (b_inv227 & c227);
  wire s228, sub228, and228, or228;
  wire b_inv228;
  assign b_inv228 = ~b228;
  assign s228  = a228 ^ b228 ^ c228;
  assign sub228 = a228 ^ b_inv228 ^ c228;
  assign and228 = a228 & b228;
  assign or228  = a228 | b228;
  assign c229 = (a228 & b228) | (a228 & c228) | (b228 & c228);
  wire c_sub229;
  assign c_sub229 = (a228 & b_inv228) | (a228 & c228) | (b_inv228 & c228);
  wire s229, sub229, and229, or229;
  wire b_inv229;
  assign b_inv229 = ~b229;
  assign s229  = a229 ^ b229 ^ c229;
  assign sub229 = a229 ^ b_inv229 ^ c229;
  assign and229 = a229 & b229;
  assign or229  = a229 | b229;
  assign c230 = (a229 & b229) | (a229 & c229) | (b229 & c229);
  wire c_sub230;
  assign c_sub230 = (a229 & b_inv229) | (a229 & c229) | (b_inv229 & c229);
  wire s230, sub230, and230, or230;
  wire b_inv230;
  assign b_inv230 = ~b230;
  assign s230  = a230 ^ b230 ^ c230;
  assign sub230 = a230 ^ b_inv230 ^ c230;
  assign and230 = a230 & b230;
  assign or230  = a230 | b230;
  assign c231 = (a230 & b230) | (a230 & c230) | (b230 & c230);
  wire c_sub231;
  assign c_sub231 = (a230 & b_inv230) | (a230 & c230) | (b_inv230 & c230);
  wire s231, sub231, and231, or231;
  wire b_inv231;
  assign b_inv231 = ~b231;
  assign s231  = a231 ^ b231 ^ c231;
  assign sub231 = a231 ^ b_inv231 ^ c231;
  assign and231 = a231 & b231;
  assign or231  = a231 | b231;
  assign c232 = (a231 & b231) | (a231 & c231) | (b231 & c231);
  wire c_sub232;
  assign c_sub232 = (a231 & b_inv231) | (a231 & c231) | (b_inv231 & c231);
  wire s232, sub232, and232, or232;
  wire b_inv232;
  assign b_inv232 = ~b232;
  assign s232  = a232 ^ b232 ^ c232;
  assign sub232 = a232 ^ b_inv232 ^ c232;
  assign and232 = a232 & b232;
  assign or232  = a232 | b232;
  assign c233 = (a232 & b232) | (a232 & c232) | (b232 & c232);
  wire c_sub233;
  assign c_sub233 = (a232 & b_inv232) | (a232 & c232) | (b_inv232 & c232);
  wire s233, sub233, and233, or233;
  wire b_inv233;
  assign b_inv233 = ~b233;
  assign s233  = a233 ^ b233 ^ c233;
  assign sub233 = a233 ^ b_inv233 ^ c233;
  assign and233 = a233 & b233;
  assign or233  = a233 | b233;
  assign c234 = (a233 & b233) | (a233 & c233) | (b233 & c233);
  wire c_sub234;
  assign c_sub234 = (a233 & b_inv233) | (a233 & c233) | (b_inv233 & c233);
  wire s234, sub234, and234, or234;
  wire b_inv234;
  assign b_inv234 = ~b234;
  assign s234  = a234 ^ b234 ^ c234;
  assign sub234 = a234 ^ b_inv234 ^ c234;
  assign and234 = a234 & b234;
  assign or234  = a234 | b234;
  assign c235 = (a234 & b234) | (a234 & c234) | (b234 & c234);
  wire c_sub235;
  assign c_sub235 = (a234 & b_inv234) | (a234 & c234) | (b_inv234 & c234);
  wire s235, sub235, and235, or235;
  wire b_inv235;
  assign b_inv235 = ~b235;
  assign s235  = a235 ^ b235 ^ c235;
  assign sub235 = a235 ^ b_inv235 ^ c235;
  assign and235 = a235 & b235;
  assign or235  = a235 | b235;
  assign c236 = (a235 & b235) | (a235 & c235) | (b235 & c235);
  wire c_sub236;
  assign c_sub236 = (a235 & b_inv235) | (a235 & c235) | (b_inv235 & c235);
  wire s236, sub236, and236, or236;
  wire b_inv236;
  assign b_inv236 = ~b236;
  assign s236  = a236 ^ b236 ^ c236;
  assign sub236 = a236 ^ b_inv236 ^ c236;
  assign and236 = a236 & b236;
  assign or236  = a236 | b236;
  assign c237 = (a236 & b236) | (a236 & c236) | (b236 & c236);
  wire c_sub237;
  assign c_sub237 = (a236 & b_inv236) | (a236 & c236) | (b_inv236 & c236);
  wire s237, sub237, and237, or237;
  wire b_inv237;
  assign b_inv237 = ~b237;
  assign s237  = a237 ^ b237 ^ c237;
  assign sub237 = a237 ^ b_inv237 ^ c237;
  assign and237 = a237 & b237;
  assign or237  = a237 | b237;
  assign c238 = (a237 & b237) | (a237 & c237) | (b237 & c237);
  wire c_sub238;
  assign c_sub238 = (a237 & b_inv237) | (a237 & c237) | (b_inv237 & c237);
  wire s238, sub238, and238, or238;
  wire b_inv238;
  assign b_inv238 = ~b238;
  assign s238  = a238 ^ b238 ^ c238;
  assign sub238 = a238 ^ b_inv238 ^ c238;
  assign and238 = a238 & b238;
  assign or238  = a238 | b238;
  assign c239 = (a238 & b238) | (a238 & c238) | (b238 & c238);
  wire c_sub239;
  assign c_sub239 = (a238 & b_inv238) | (a238 & c238) | (b_inv238 & c238);
  wire s239, sub239, and239, or239;
  wire b_inv239;
  assign b_inv239 = ~b239;
  assign s239  = a239 ^ b239 ^ c239;
  assign sub239 = a239 ^ b_inv239 ^ c239;
  assign and239 = a239 & b239;
  assign or239  = a239 | b239;
  assign c240 = (a239 & b239) | (a239 & c239) | (b239 & c239);
  wire c_sub240;
  assign c_sub240 = (a239 & b_inv239) | (a239 & c239) | (b_inv239 & c239);
  wire s240, sub240, and240, or240;
  wire b_inv240;
  assign b_inv240 = ~b240;
  assign s240  = a240 ^ b240 ^ c240;
  assign sub240 = a240 ^ b_inv240 ^ c240;
  assign and240 = a240 & b240;
  assign or240  = a240 | b240;
  assign c241 = (a240 & b240) | (a240 & c240) | (b240 & c240);
  wire c_sub241;
  assign c_sub241 = (a240 & b_inv240) | (a240 & c240) | (b_inv240 & c240);
  wire s241, sub241, and241, or241;
  wire b_inv241;
  assign b_inv241 = ~b241;
  assign s241  = a241 ^ b241 ^ c241;
  assign sub241 = a241 ^ b_inv241 ^ c241;
  assign and241 = a241 & b241;
  assign or241  = a241 | b241;
  assign c242 = (a241 & b241) | (a241 & c241) | (b241 & c241);
  wire c_sub242;
  assign c_sub242 = (a241 & b_inv241) | (a241 & c241) | (b_inv241 & c241);
  wire s242, sub242, and242, or242;
  wire b_inv242;
  assign b_inv242 = ~b242;
  assign s242  = a242 ^ b242 ^ c242;
  assign sub242 = a242 ^ b_inv242 ^ c242;
  assign and242 = a242 & b242;
  assign or242  = a242 | b242;
  assign c243 = (a242 & b242) | (a242 & c242) | (b242 & c242);
  wire c_sub243;
  assign c_sub243 = (a242 & b_inv242) | (a242 & c242) | (b_inv242 & c242);
  wire s243, sub243, and243, or243;
  wire b_inv243;
  assign b_inv243 = ~b243;
  assign s243  = a243 ^ b243 ^ c243;
  assign sub243 = a243 ^ b_inv243 ^ c243;
  assign and243 = a243 & b243;
  assign or243  = a243 | b243;
  assign c244 = (a243 & b243) | (a243 & c243) | (b243 & c243);
  wire c_sub244;
  assign c_sub244 = (a243 & b_inv243) | (a243 & c243) | (b_inv243 & c243);
  wire s244, sub244, and244, or244;
  wire b_inv244;
  assign b_inv244 = ~b244;
  assign s244  = a244 ^ b244 ^ c244;
  assign sub244 = a244 ^ b_inv244 ^ c244;
  assign and244 = a244 & b244;
  assign or244  = a244 | b244;
  assign c245 = (a244 & b244) | (a244 & c244) | (b244 & c244);
  wire c_sub245;
  assign c_sub245 = (a244 & b_inv244) | (a244 & c244) | (b_inv244 & c244);
  wire s245, sub245, and245, or245;
  wire b_inv245;
  assign b_inv245 = ~b245;
  assign s245  = a245 ^ b245 ^ c245;
  assign sub245 = a245 ^ b_inv245 ^ c245;
  assign and245 = a245 & b245;
  assign or245  = a245 | b245;
  assign c246 = (a245 & b245) | (a245 & c245) | (b245 & c245);
  wire c_sub246;
  assign c_sub246 = (a245 & b_inv245) | (a245 & c245) | (b_inv245 & c245);
  wire s246, sub246, and246, or246;
  wire b_inv246;
  assign b_inv246 = ~b246;
  assign s246  = a246 ^ b246 ^ c246;
  assign sub246 = a246 ^ b_inv246 ^ c246;
  assign and246 = a246 & b246;
  assign or246  = a246 | b246;
  assign c247 = (a246 & b246) | (a246 & c246) | (b246 & c246);
  wire c_sub247;
  assign c_sub247 = (a246 & b_inv246) | (a246 & c246) | (b_inv246 & c246);
  wire s247, sub247, and247, or247;
  wire b_inv247;
  assign b_inv247 = ~b247;
  assign s247  = a247 ^ b247 ^ c247;
  assign sub247 = a247 ^ b_inv247 ^ c247;
  assign and247 = a247 & b247;
  assign or247  = a247 | b247;
  assign c248 = (a247 & b247) | (a247 & c247) | (b247 & c247);
  wire c_sub248;
  assign c_sub248 = (a247 & b_inv247) | (a247 & c247) | (b_inv247 & c247);
  wire s248, sub248, and248, or248;
  wire b_inv248;
  assign b_inv248 = ~b248;
  assign s248  = a248 ^ b248 ^ c248;
  assign sub248 = a248 ^ b_inv248 ^ c248;
  assign and248 = a248 & b248;
  assign or248  = a248 | b248;
  assign c249 = (a248 & b248) | (a248 & c248) | (b248 & c248);
  wire c_sub249;
  assign c_sub249 = (a248 & b_inv248) | (a248 & c248) | (b_inv248 & c248);
  wire s249, sub249, and249, or249;
  wire b_inv249;
  assign b_inv249 = ~b249;
  assign s249  = a249 ^ b249 ^ c249;
  assign sub249 = a249 ^ b_inv249 ^ c249;
  assign and249 = a249 & b249;
  assign or249  = a249 | b249;
  assign c250 = (a249 & b249) | (a249 & c249) | (b249 & c249);
  wire c_sub250;
  assign c_sub250 = (a249 & b_inv249) | (a249 & c249) | (b_inv249 & c249);
  wire s250, sub250, and250, or250;
  wire b_inv250;
  assign b_inv250 = ~b250;
  assign s250  = a250 ^ b250 ^ c250;
  assign sub250 = a250 ^ b_inv250 ^ c250;
  assign and250 = a250 & b250;
  assign or250  = a250 | b250;
  assign c251 = (a250 & b250) | (a250 & c250) | (b250 & c250);
  wire c_sub251;
  assign c_sub251 = (a250 & b_inv250) | (a250 & c250) | (b_inv250 & c250);
  wire s251, sub251, and251, or251;
  wire b_inv251;
  assign b_inv251 = ~b251;
  assign s251  = a251 ^ b251 ^ c251;
  assign sub251 = a251 ^ b_inv251 ^ c251;
  assign and251 = a251 & b251;
  assign or251  = a251 | b251;
  assign c252 = (a251 & b251) | (a251 & c251) | (b251 & c251);
  wire c_sub252;
  assign c_sub252 = (a251 & b_inv251) | (a251 & c251) | (b_inv251 & c251);
  wire s252, sub252, and252, or252;
  wire b_inv252;
  assign b_inv252 = ~b252;
  assign s252  = a252 ^ b252 ^ c252;
  assign sub252 = a252 ^ b_inv252 ^ c252;
  assign and252 = a252 & b252;
  assign or252  = a252 | b252;
  assign c253 = (a252 & b252) | (a252 & c252) | (b252 & c252);
  wire c_sub253;
  assign c_sub253 = (a252 & b_inv252) | (a252 & c252) | (b_inv252 & c252);
  wire s253, sub253, and253, or253;
  wire b_inv253;
  assign b_inv253 = ~b253;
  assign s253  = a253 ^ b253 ^ c253;
  assign sub253 = a253 ^ b_inv253 ^ c253;
  assign and253 = a253 & b253;
  assign or253  = a253 | b253;
  assign c254 = (a253 & b253) | (a253 & c253) | (b253 & c253);
  wire c_sub254;
  assign c_sub254 = (a253 & b_inv253) | (a253 & c253) | (b_inv253 & c253);
  wire s254, sub254, and254, or254;
  wire b_inv254;
  assign b_inv254 = ~b254;
  assign s254  = a254 ^ b254 ^ c254;
  assign sub254 = a254 ^ b_inv254 ^ c254;
  assign and254 = a254 & b254;
  assign or254  = a254 | b254;
  assign c255 = (a254 & b254) | (a254 & c254) | (b254 & c254);
  wire c_sub255;
  assign c_sub255 = (a254 & b_inv254) | (a254 & c254) | (b_inv254 & c254);
  wire s255, sub255, and255, or255;
  wire b_inv255;
  assign b_inv255 = ~b255;
  assign s255  = a255 ^ b255 ^ c255;
  assign sub255 = a255 ^ b_inv255 ^ c255;
  assign and255 = a255 & b255;
  assign or255  = a255 | b255;
  assign c256 = (a255 & b255) | (a255 & c255) | (b255 & c255);
  wire c_sub256;
  assign c_sub256 = (a255 & b_inv255) | (a255 & c255) | (b_inv255 & c255);
  wire s256, sub256, and256, or256;
  wire b_inv256;
  assign b_inv256 = ~b256;
  assign s256  = a256 ^ b256 ^ c256;
  assign sub256 = a256 ^ b_inv256 ^ c256;
  assign and256 = a256 & b256;
  assign or256  = a256 | b256;
  assign c257 = (a256 & b256) | (a256 & c256) | (b256 & c256);
  wire c_sub257;
  assign c_sub257 = (a256 & b_inv256) | (a256 & c256) | (b_inv256 & c256);
  wire s257, sub257, and257, or257;
  wire b_inv257;
  assign b_inv257 = ~b257;
  assign s257  = a257 ^ b257 ^ c257;
  assign sub257 = a257 ^ b_inv257 ^ c257;
  assign and257 = a257 & b257;
  assign or257  = a257 | b257;
  assign c258 = (a257 & b257) | (a257 & c257) | (b257 & c257);
  wire c_sub258;
  assign c_sub258 = (a257 & b_inv257) | (a257 & c257) | (b_inv257 & c257);
  wire s258, sub258, and258, or258;
  wire b_inv258;
  assign b_inv258 = ~b258;
  assign s258  = a258 ^ b258 ^ c258;
  assign sub258 = a258 ^ b_inv258 ^ c258;
  assign and258 = a258 & b258;
  assign or258  = a258 | b258;
  assign c259 = (a258 & b258) | (a258 & c258) | (b258 & c258);
  wire c_sub259;
  assign c_sub259 = (a258 & b_inv258) | (a258 & c258) | (b_inv258 & c258);
  wire s259, sub259, and259, or259;
  wire b_inv259;
  assign b_inv259 = ~b259;
  assign s259  = a259 ^ b259 ^ c259;
  assign sub259 = a259 ^ b_inv259 ^ c259;
  assign and259 = a259 & b259;
  assign or259  = a259 | b259;
  assign c260 = (a259 & b259) | (a259 & c259) | (b259 & c259);
  wire c_sub260;
  assign c_sub260 = (a259 & b_inv259) | (a259 & c259) | (b_inv259 & c259);
  wire s260, sub260, and260, or260;
  wire b_inv260;
  assign b_inv260 = ~b260;
  assign s260  = a260 ^ b260 ^ c260;
  assign sub260 = a260 ^ b_inv260 ^ c260;
  assign and260 = a260 & b260;
  assign or260  = a260 | b260;
  assign c261 = (a260 & b260) | (a260 & c260) | (b260 & c260);
  wire c_sub261;
  assign c_sub261 = (a260 & b_inv260) | (a260 & c260) | (b_inv260 & c260);
  wire s261, sub261, and261, or261;
  wire b_inv261;
  assign b_inv261 = ~b261;
  assign s261  = a261 ^ b261 ^ c261;
  assign sub261 = a261 ^ b_inv261 ^ c261;
  assign and261 = a261 & b261;
  assign or261  = a261 | b261;
  assign c262 = (a261 & b261) | (a261 & c261) | (b261 & c261);
  wire c_sub262;
  assign c_sub262 = (a261 & b_inv261) | (a261 & c261) | (b_inv261 & c261);
  wire s262, sub262, and262, or262;
  wire b_inv262;
  assign b_inv262 = ~b262;
  assign s262  = a262 ^ b262 ^ c262;
  assign sub262 = a262 ^ b_inv262 ^ c262;
  assign and262 = a262 & b262;
  assign or262  = a262 | b262;
  assign c263 = (a262 & b262) | (a262 & c262) | (b262 & c262);
  wire c_sub263;
  assign c_sub263 = (a262 & b_inv262) | (a262 & c262) | (b_inv262 & c262);
  wire s263, sub263, and263, or263;
  wire b_inv263;
  assign b_inv263 = ~b263;
  assign s263  = a263 ^ b263 ^ c263;
  assign sub263 = a263 ^ b_inv263 ^ c263;
  assign and263 = a263 & b263;
  assign or263  = a263 | b263;
  assign c264 = (a263 & b263) | (a263 & c263) | (b263 & c263);
  wire c_sub264;
  assign c_sub264 = (a263 & b_inv263) | (a263 & c263) | (b_inv263 & c263);
  wire s264, sub264, and264, or264;
  wire b_inv264;
  assign b_inv264 = ~b264;
  assign s264  = a264 ^ b264 ^ c264;
  assign sub264 = a264 ^ b_inv264 ^ c264;
  assign and264 = a264 & b264;
  assign or264  = a264 | b264;
  assign c265 = (a264 & b264) | (a264 & c264) | (b264 & c264);
  wire c_sub265;
  assign c_sub265 = (a264 & b_inv264) | (a264 & c264) | (b_inv264 & c264);
  wire s265, sub265, and265, or265;
  wire b_inv265;
  assign b_inv265 = ~b265;
  assign s265  = a265 ^ b265 ^ c265;
  assign sub265 = a265 ^ b_inv265 ^ c265;
  assign and265 = a265 & b265;
  assign or265  = a265 | b265;
  assign c266 = (a265 & b265) | (a265 & c265) | (b265 & c265);
  wire c_sub266;
  assign c_sub266 = (a265 & b_inv265) | (a265 & c265) | (b_inv265 & c265);
  wire s266, sub266, and266, or266;
  wire b_inv266;
  assign b_inv266 = ~b266;
  assign s266  = a266 ^ b266 ^ c266;
  assign sub266 = a266 ^ b_inv266 ^ c266;
  assign and266 = a266 & b266;
  assign or266  = a266 | b266;
  assign c267 = (a266 & b266) | (a266 & c266) | (b266 & c266);
  wire c_sub267;
  assign c_sub267 = (a266 & b_inv266) | (a266 & c266) | (b_inv266 & c266);
  wire s267, sub267, and267, or267;
  wire b_inv267;
  assign b_inv267 = ~b267;
  assign s267  = a267 ^ b267 ^ c267;
  assign sub267 = a267 ^ b_inv267 ^ c267;
  assign and267 = a267 & b267;
  assign or267  = a267 | b267;
  assign c268 = (a267 & b267) | (a267 & c267) | (b267 & c267);
  wire c_sub268;
  assign c_sub268 = (a267 & b_inv267) | (a267 & c267) | (b_inv267 & c267);
  wire s268, sub268, and268, or268;
  wire b_inv268;
  assign b_inv268 = ~b268;
  assign s268  = a268 ^ b268 ^ c268;
  assign sub268 = a268 ^ b_inv268 ^ c268;
  assign and268 = a268 & b268;
  assign or268  = a268 | b268;
  assign c269 = (a268 & b268) | (a268 & c268) | (b268 & c268);
  wire c_sub269;
  assign c_sub269 = (a268 & b_inv268) | (a268 & c268) | (b_inv268 & c268);
  wire s269, sub269, and269, or269;
  wire b_inv269;
  assign b_inv269 = ~b269;
  assign s269  = a269 ^ b269 ^ c269;
  assign sub269 = a269 ^ b_inv269 ^ c269;
  assign and269 = a269 & b269;
  assign or269  = a269 | b269;
  assign c270 = (a269 & b269) | (a269 & c269) | (b269 & c269);
  wire c_sub270;
  assign c_sub270 = (a269 & b_inv269) | (a269 & c269) | (b_inv269 & c269);
  wire s270, sub270, and270, or270;
  wire b_inv270;
  assign b_inv270 = ~b270;
  assign s270  = a270 ^ b270 ^ c270;
  assign sub270 = a270 ^ b_inv270 ^ c270;
  assign and270 = a270 & b270;
  assign or270  = a270 | b270;
  assign c271 = (a270 & b270) | (a270 & c270) | (b270 & c270);
  wire c_sub271;
  assign c_sub271 = (a270 & b_inv270) | (a270 & c270) | (b_inv270 & c270);
  wire s271, sub271, and271, or271;
  wire b_inv271;
  assign b_inv271 = ~b271;
  assign s271  = a271 ^ b271 ^ c271;
  assign sub271 = a271 ^ b_inv271 ^ c271;
  assign and271 = a271 & b271;
  assign or271  = a271 | b271;
  assign c272 = (a271 & b271) | (a271 & c271) | (b271 & c271);
  wire c_sub272;
  assign c_sub272 = (a271 & b_inv271) | (a271 & c271) | (b_inv271 & c271);
  wire s272, sub272, and272, or272;
  wire b_inv272;
  assign b_inv272 = ~b272;
  assign s272  = a272 ^ b272 ^ c272;
  assign sub272 = a272 ^ b_inv272 ^ c272;
  assign and272 = a272 & b272;
  assign or272  = a272 | b272;
  assign c273 = (a272 & b272) | (a272 & c272) | (b272 & c272);
  wire c_sub273;
  assign c_sub273 = (a272 & b_inv272) | (a272 & c272) | (b_inv272 & c272);
  wire s273, sub273, and273, or273;
  wire b_inv273;
  assign b_inv273 = ~b273;
  assign s273  = a273 ^ b273 ^ c273;
  assign sub273 = a273 ^ b_inv273 ^ c273;
  assign and273 = a273 & b273;
  assign or273  = a273 | b273;
  assign c274 = (a273 & b273) | (a273 & c273) | (b273 & c273);
  wire c_sub274;
  assign c_sub274 = (a273 & b_inv273) | (a273 & c273) | (b_inv273 & c273);
  wire s274, sub274, and274, or274;
  wire b_inv274;
  assign b_inv274 = ~b274;
  assign s274  = a274 ^ b274 ^ c274;
  assign sub274 = a274 ^ b_inv274 ^ c274;
  assign and274 = a274 & b274;
  assign or274  = a274 | b274;
  assign c275 = (a274 & b274) | (a274 & c274) | (b274 & c274);
  wire c_sub275;
  assign c_sub275 = (a274 & b_inv274) | (a274 & c274) | (b_inv274 & c274);
  wire s275, sub275, and275, or275;
  wire b_inv275;
  assign b_inv275 = ~b275;
  assign s275  = a275 ^ b275 ^ c275;
  assign sub275 = a275 ^ b_inv275 ^ c275;
  assign and275 = a275 & b275;
  assign or275  = a275 | b275;
  assign c276 = (a275 & b275) | (a275 & c275) | (b275 & c275);
  wire c_sub276;
  assign c_sub276 = (a275 & b_inv275) | (a275 & c275) | (b_inv275 & c275);
  wire s276, sub276, and276, or276;
  wire b_inv276;
  assign b_inv276 = ~b276;
  assign s276  = a276 ^ b276 ^ c276;
  assign sub276 = a276 ^ b_inv276 ^ c276;
  assign and276 = a276 & b276;
  assign or276  = a276 | b276;
  assign c277 = (a276 & b276) | (a276 & c276) | (b276 & c276);
  wire c_sub277;
  assign c_sub277 = (a276 & b_inv276) | (a276 & c276) | (b_inv276 & c276);
  wire s277, sub277, and277, or277;
  wire b_inv277;
  assign b_inv277 = ~b277;
  assign s277  = a277 ^ b277 ^ c277;
  assign sub277 = a277 ^ b_inv277 ^ c277;
  assign and277 = a277 & b277;
  assign or277  = a277 | b277;
  assign c278 = (a277 & b277) | (a277 & c277) | (b277 & c277);
  wire c_sub278;
  assign c_sub278 = (a277 & b_inv277) | (a277 & c277) | (b_inv277 & c277);
  wire s278, sub278, and278, or278;
  wire b_inv278;
  assign b_inv278 = ~b278;
  assign s278  = a278 ^ b278 ^ c278;
  assign sub278 = a278 ^ b_inv278 ^ c278;
  assign and278 = a278 & b278;
  assign or278  = a278 | b278;
  assign c279 = (a278 & b278) | (a278 & c278) | (b278 & c278);
  wire c_sub279;
  assign c_sub279 = (a278 & b_inv278) | (a278 & c278) | (b_inv278 & c278);
  wire s279, sub279, and279, or279;
  wire b_inv279;
  assign b_inv279 = ~b279;
  assign s279  = a279 ^ b279 ^ c279;
  assign sub279 = a279 ^ b_inv279 ^ c279;
  assign and279 = a279 & b279;
  assign or279  = a279 | b279;
  assign c280 = (a279 & b279) | (a279 & c279) | (b279 & c279);
  wire c_sub280;
  assign c_sub280 = (a279 & b_inv279) | (a279 & c279) | (b_inv279 & c279);
  wire s280, sub280, and280, or280;
  wire b_inv280;
  assign b_inv280 = ~b280;
  assign s280  = a280 ^ b280 ^ c280;
  assign sub280 = a280 ^ b_inv280 ^ c280;
  assign and280 = a280 & b280;
  assign or280  = a280 | b280;
  assign c281 = (a280 & b280) | (a280 & c280) | (b280 & c280);
  wire c_sub281;
  assign c_sub281 = (a280 & b_inv280) | (a280 & c280) | (b_inv280 & c280);
  wire s281, sub281, and281, or281;
  wire b_inv281;
  assign b_inv281 = ~b281;
  assign s281  = a281 ^ b281 ^ c281;
  assign sub281 = a281 ^ b_inv281 ^ c281;
  assign and281 = a281 & b281;
  assign or281  = a281 | b281;
  assign c282 = (a281 & b281) | (a281 & c281) | (b281 & c281);
  wire c_sub282;
  assign c_sub282 = (a281 & b_inv281) | (a281 & c281) | (b_inv281 & c281);
  wire s282, sub282, and282, or282;
  wire b_inv282;
  assign b_inv282 = ~b282;
  assign s282  = a282 ^ b282 ^ c282;
  assign sub282 = a282 ^ b_inv282 ^ c282;
  assign and282 = a282 & b282;
  assign or282  = a282 | b282;
  assign c283 = (a282 & b282) | (a282 & c282) | (b282 & c282);
  wire c_sub283;
  assign c_sub283 = (a282 & b_inv282) | (a282 & c282) | (b_inv282 & c282);
  wire s283, sub283, and283, or283;
  wire b_inv283;
  assign b_inv283 = ~b283;
  assign s283  = a283 ^ b283 ^ c283;
  assign sub283 = a283 ^ b_inv283 ^ c283;
  assign and283 = a283 & b283;
  assign or283  = a283 | b283;
  assign c284 = (a283 & b283) | (a283 & c283) | (b283 & c283);
  wire c_sub284;
  assign c_sub284 = (a283 & b_inv283) | (a283 & c283) | (b_inv283 & c283);
  wire s284, sub284, and284, or284;
  wire b_inv284;
  assign b_inv284 = ~b284;
  assign s284  = a284 ^ b284 ^ c284;
  assign sub284 = a284 ^ b_inv284 ^ c284;
  assign and284 = a284 & b284;
  assign or284  = a284 | b284;
  assign c285 = (a284 & b284) | (a284 & c284) | (b284 & c284);
  wire c_sub285;
  assign c_sub285 = (a284 & b_inv284) | (a284 & c284) | (b_inv284 & c284);
  wire s285, sub285, and285, or285;
  wire b_inv285;
  assign b_inv285 = ~b285;
  assign s285  = a285 ^ b285 ^ c285;
  assign sub285 = a285 ^ b_inv285 ^ c285;
  assign and285 = a285 & b285;
  assign or285  = a285 | b285;
  assign c286 = (a285 & b285) | (a285 & c285) | (b285 & c285);
  wire c_sub286;
  assign c_sub286 = (a285 & b_inv285) | (a285 & c285) | (b_inv285 & c285);
  wire s286, sub286, and286, or286;
  wire b_inv286;
  assign b_inv286 = ~b286;
  assign s286  = a286 ^ b286 ^ c286;
  assign sub286 = a286 ^ b_inv286 ^ c286;
  assign and286 = a286 & b286;
  assign or286  = a286 | b286;
  assign c287 = (a286 & b286) | (a286 & c286) | (b286 & c286);
  wire c_sub287;
  assign c_sub287 = (a286 & b_inv286) | (a286 & c286) | (b_inv286 & c286);
  wire s287, sub287, and287, or287;
  wire b_inv287;
  assign b_inv287 = ~b287;
  assign s287  = a287 ^ b287 ^ c287;
  assign sub287 = a287 ^ b_inv287 ^ c287;
  assign and287 = a287 & b287;
  assign or287  = a287 | b287;
  assign c288 = (a287 & b287) | (a287 & c287) | (b287 & c287);
  wire c_sub288;
  assign c_sub288 = (a287 & b_inv287) | (a287 & c287) | (b_inv287 & c287);
  wire s288, sub288, and288, or288;
  wire b_inv288;
  assign b_inv288 = ~b288;
  assign s288  = a288 ^ b288 ^ c288;
  assign sub288 = a288 ^ b_inv288 ^ c288;
  assign and288 = a288 & b288;
  assign or288  = a288 | b288;
  assign c289 = (a288 & b288) | (a288 & c288) | (b288 & c288);
  wire c_sub289;
  assign c_sub289 = (a288 & b_inv288) | (a288 & c288) | (b_inv288 & c288);
  wire s289, sub289, and289, or289;
  wire b_inv289;
  assign b_inv289 = ~b289;
  assign s289  = a289 ^ b289 ^ c289;
  assign sub289 = a289 ^ b_inv289 ^ c289;
  assign and289 = a289 & b289;
  assign or289  = a289 | b289;
  assign c290 = (a289 & b289) | (a289 & c289) | (b289 & c289);
  wire c_sub290;
  assign c_sub290 = (a289 & b_inv289) | (a289 & c289) | (b_inv289 & c289);
  wire s290, sub290, and290, or290;
  wire b_inv290;
  assign b_inv290 = ~b290;
  assign s290  = a290 ^ b290 ^ c290;
  assign sub290 = a290 ^ b_inv290 ^ c290;
  assign and290 = a290 & b290;
  assign or290  = a290 | b290;
  assign c291 = (a290 & b290) | (a290 & c290) | (b290 & c290);
  wire c_sub291;
  assign c_sub291 = (a290 & b_inv290) | (a290 & c290) | (b_inv290 & c290);
  wire s291, sub291, and291, or291;
  wire b_inv291;
  assign b_inv291 = ~b291;
  assign s291  = a291 ^ b291 ^ c291;
  assign sub291 = a291 ^ b_inv291 ^ c291;
  assign and291 = a291 & b291;
  assign or291  = a291 | b291;
  assign c292 = (a291 & b291) | (a291 & c291) | (b291 & c291);
  wire c_sub292;
  assign c_sub292 = (a291 & b_inv291) | (a291 & c291) | (b_inv291 & c291);
  wire s292, sub292, and292, or292;
  wire b_inv292;
  assign b_inv292 = ~b292;
  assign s292  = a292 ^ b292 ^ c292;
  assign sub292 = a292 ^ b_inv292 ^ c292;
  assign and292 = a292 & b292;
  assign or292  = a292 | b292;
  assign c293 = (a292 & b292) | (a292 & c292) | (b292 & c292);
  wire c_sub293;
  assign c_sub293 = (a292 & b_inv292) | (a292 & c292) | (b_inv292 & c292);
  wire s293, sub293, and293, or293;
  wire b_inv293;
  assign b_inv293 = ~b293;
  assign s293  = a293 ^ b293 ^ c293;
  assign sub293 = a293 ^ b_inv293 ^ c293;
  assign and293 = a293 & b293;
  assign or293  = a293 | b293;
  assign c294 = (a293 & b293) | (a293 & c293) | (b293 & c293);
  wire c_sub294;
  assign c_sub294 = (a293 & b_inv293) | (a293 & c293) | (b_inv293 & c293);
  wire s294, sub294, and294, or294;
  wire b_inv294;
  assign b_inv294 = ~b294;
  assign s294  = a294 ^ b294 ^ c294;
  assign sub294 = a294 ^ b_inv294 ^ c294;
  assign and294 = a294 & b294;
  assign or294  = a294 | b294;
  assign c295 = (a294 & b294) | (a294 & c294) | (b294 & c294);
  wire c_sub295;
  assign c_sub295 = (a294 & b_inv294) | (a294 & c294) | (b_inv294 & c294);
  wire s295, sub295, and295, or295;
  wire b_inv295;
  assign b_inv295 = ~b295;
  assign s295  = a295 ^ b295 ^ c295;
  assign sub295 = a295 ^ b_inv295 ^ c295;
  assign and295 = a295 & b295;
  assign or295  = a295 | b295;
  assign c296 = (a295 & b295) | (a295 & c295) | (b295 & c295);
  wire c_sub296;
  assign c_sub296 = (a295 & b_inv295) | (a295 & c295) | (b_inv295 & c295);
  wire s296, sub296, and296, or296;
  wire b_inv296;
  assign b_inv296 = ~b296;
  assign s296  = a296 ^ b296 ^ c296;
  assign sub296 = a296 ^ b_inv296 ^ c296;
  assign and296 = a296 & b296;
  assign or296  = a296 | b296;
  assign c297 = (a296 & b296) | (a296 & c296) | (b296 & c296);
  wire c_sub297;
  assign c_sub297 = (a296 & b_inv296) | (a296 & c296) | (b_inv296 & c296);
  wire s297, sub297, and297, or297;
  wire b_inv297;
  assign b_inv297 = ~b297;
  assign s297  = a297 ^ b297 ^ c297;
  assign sub297 = a297 ^ b_inv297 ^ c297;
  assign and297 = a297 & b297;
  assign or297  = a297 | b297;
  assign c298 = (a297 & b297) | (a297 & c297) | (b297 & c297);
  wire c_sub298;
  assign c_sub298 = (a297 & b_inv297) | (a297 & c297) | (b_inv297 & c297);
  wire s298, sub298, and298, or298;
  wire b_inv298;
  assign b_inv298 = ~b298;
  assign s298  = a298 ^ b298 ^ c298;
  assign sub298 = a298 ^ b_inv298 ^ c298;
  assign and298 = a298 & b298;
  assign or298  = a298 | b298;
  assign c299 = (a298 & b298) | (a298 & c298) | (b298 & c298);
  wire c_sub299;
  assign c_sub299 = (a298 & b_inv298) | (a298 & c298) | (b_inv298 & c298);
  wire s299, sub299, and299, or299;
  wire b_inv299;
  assign b_inv299 = ~b299;
  assign s299  = a299 ^ b299 ^ c299;
  assign sub299 = a299 ^ b_inv299 ^ c299;
  assign and299 = a299 & b299;
  assign or299  = a299 | b299;
  assign c300 = (a299 & b299) | (a299 & c299) | (b299 & c299);
  wire c_sub300;
  assign c_sub300 = (a299 & b_inv299) | (a299 & c299) | (b_inv299 & c299);
  wire s300, sub300, and300, or300;
  wire b_inv300;
  assign b_inv300 = ~b300;
  assign s300  = a300 ^ b300 ^ c300;
  assign sub300 = a300 ^ b_inv300 ^ c300;
  assign and300 = a300 & b300;
  assign or300  = a300 | b300;
  assign c301 = (a300 & b300) | (a300 & c300) | (b300 & c300);
  wire c_sub301;
  assign c_sub301 = (a300 & b_inv300) | (a300 & c300) | (b_inv300 & c300);
  wire s301, sub301, and301, or301;
  wire b_inv301;
  assign b_inv301 = ~b301;
  assign s301  = a301 ^ b301 ^ c301;
  assign sub301 = a301 ^ b_inv301 ^ c301;
  assign and301 = a301 & b301;
  assign or301  = a301 | b301;
  assign c302 = (a301 & b301) | (a301 & c301) | (b301 & c301);
  wire c_sub302;
  assign c_sub302 = (a301 & b_inv301) | (a301 & c301) | (b_inv301 & c301);
  wire s302, sub302, and302, or302;
  wire b_inv302;
  assign b_inv302 = ~b302;
  assign s302  = a302 ^ b302 ^ c302;
  assign sub302 = a302 ^ b_inv302 ^ c302;
  assign and302 = a302 & b302;
  assign or302  = a302 | b302;
  assign c303 = (a302 & b302) | (a302 & c302) | (b302 & c302);
  wire c_sub303;
  assign c_sub303 = (a302 & b_inv302) | (a302 & c302) | (b_inv302 & c302);
  wire s303, sub303, and303, or303;
  wire b_inv303;
  assign b_inv303 = ~b303;
  assign s303  = a303 ^ b303 ^ c303;
  assign sub303 = a303 ^ b_inv303 ^ c303;
  assign and303 = a303 & b303;
  assign or303  = a303 | b303;
  assign c304 = (a303 & b303) | (a303 & c303) | (b303 & c303);
  wire c_sub304;
  assign c_sub304 = (a303 & b_inv303) | (a303 & c303) | (b_inv303 & c303);
  wire s304, sub304, and304, or304;
  wire b_inv304;
  assign b_inv304 = ~b304;
  assign s304  = a304 ^ b304 ^ c304;
  assign sub304 = a304 ^ b_inv304 ^ c304;
  assign and304 = a304 & b304;
  assign or304  = a304 | b304;
  assign c305 = (a304 & b304) | (a304 & c304) | (b304 & c304);
  wire c_sub305;
  assign c_sub305 = (a304 & b_inv304) | (a304 & c304) | (b_inv304 & c304);
  wire s305, sub305, and305, or305;
  wire b_inv305;
  assign b_inv305 = ~b305;
  assign s305  = a305 ^ b305 ^ c305;
  assign sub305 = a305 ^ b_inv305 ^ c305;
  assign and305 = a305 & b305;
  assign or305  = a305 | b305;
  assign c306 = (a305 & b305) | (a305 & c305) | (b305 & c305);
  wire c_sub306;
  assign c_sub306 = (a305 & b_inv305) | (a305 & c305) | (b_inv305 & c305);
  wire s306, sub306, and306, or306;
  wire b_inv306;
  assign b_inv306 = ~b306;
  assign s306  = a306 ^ b306 ^ c306;
  assign sub306 = a306 ^ b_inv306 ^ c306;
  assign and306 = a306 & b306;
  assign or306  = a306 | b306;
  assign c307 = (a306 & b306) | (a306 & c306) | (b306 & c306);
  wire c_sub307;
  assign c_sub307 = (a306 & b_inv306) | (a306 & c306) | (b_inv306 & c306);
  wire s307, sub307, and307, or307;
  wire b_inv307;
  assign b_inv307 = ~b307;
  assign s307  = a307 ^ b307 ^ c307;
  assign sub307 = a307 ^ b_inv307 ^ c307;
  assign and307 = a307 & b307;
  assign or307  = a307 | b307;
  assign c308 = (a307 & b307) | (a307 & c307) | (b307 & c307);
  wire c_sub308;
  assign c_sub308 = (a307 & b_inv307) | (a307 & c307) | (b_inv307 & c307);
  wire s308, sub308, and308, or308;
  wire b_inv308;
  assign b_inv308 = ~b308;
  assign s308  = a308 ^ b308 ^ c308;
  assign sub308 = a308 ^ b_inv308 ^ c308;
  assign and308 = a308 & b308;
  assign or308  = a308 | b308;
  assign c309 = (a308 & b308) | (a308 & c308) | (b308 & c308);
  wire c_sub309;
  assign c_sub309 = (a308 & b_inv308) | (a308 & c308) | (b_inv308 & c308);
  wire s309, sub309, and309, or309;
  wire b_inv309;
  assign b_inv309 = ~b309;
  assign s309  = a309 ^ b309 ^ c309;
  assign sub309 = a309 ^ b_inv309 ^ c309;
  assign and309 = a309 & b309;
  assign or309  = a309 | b309;
  assign c310 = (a309 & b309) | (a309 & c309) | (b309 & c309);
  wire c_sub310;
  assign c_sub310 = (a309 & b_inv309) | (a309 & c309) | (b_inv309 & c309);
  wire s310, sub310, and310, or310;
  wire b_inv310;
  assign b_inv310 = ~b310;
  assign s310  = a310 ^ b310 ^ c310;
  assign sub310 = a310 ^ b_inv310 ^ c310;
  assign and310 = a310 & b310;
  assign or310  = a310 | b310;
  assign c311 = (a310 & b310) | (a310 & c310) | (b310 & c310);
  wire c_sub311;
  assign c_sub311 = (a310 & b_inv310) | (a310 & c310) | (b_inv310 & c310);
  wire s311, sub311, and311, or311;
  wire b_inv311;
  assign b_inv311 = ~b311;
  assign s311  = a311 ^ b311 ^ c311;
  assign sub311 = a311 ^ b_inv311 ^ c311;
  assign and311 = a311 & b311;
  assign or311  = a311 | b311;
  assign c312 = (a311 & b311) | (a311 & c311) | (b311 & c311);
  wire c_sub312;
  assign c_sub312 = (a311 & b_inv311) | (a311 & c311) | (b_inv311 & c311);
  wire s312, sub312, and312, or312;
  wire b_inv312;
  assign b_inv312 = ~b312;
  assign s312  = a312 ^ b312 ^ c312;
  assign sub312 = a312 ^ b_inv312 ^ c312;
  assign and312 = a312 & b312;
  assign or312  = a312 | b312;
  assign c313 = (a312 & b312) | (a312 & c312) | (b312 & c312);
  wire c_sub313;
  assign c_sub313 = (a312 & b_inv312) | (a312 & c312) | (b_inv312 & c312);
  wire s313, sub313, and313, or313;
  wire b_inv313;
  assign b_inv313 = ~b313;
  assign s313  = a313 ^ b313 ^ c313;
  assign sub313 = a313 ^ b_inv313 ^ c313;
  assign and313 = a313 & b313;
  assign or313  = a313 | b313;
  assign c314 = (a313 & b313) | (a313 & c313) | (b313 & c313);
  wire c_sub314;
  assign c_sub314 = (a313 & b_inv313) | (a313 & c313) | (b_inv313 & c313);
  wire s314, sub314, and314, or314;
  wire b_inv314;
  assign b_inv314 = ~b314;
  assign s314  = a314 ^ b314 ^ c314;
  assign sub314 = a314 ^ b_inv314 ^ c314;
  assign and314 = a314 & b314;
  assign or314  = a314 | b314;
  assign c315 = (a314 & b314) | (a314 & c314) | (b314 & c314);
  wire c_sub315;
  assign c_sub315 = (a314 & b_inv314) | (a314 & c314) | (b_inv314 & c314);
  wire s315, sub315, and315, or315;
  wire b_inv315;
  assign b_inv315 = ~b315;
  assign s315  = a315 ^ b315 ^ c315;
  assign sub315 = a315 ^ b_inv315 ^ c315;
  assign and315 = a315 & b315;
  assign or315  = a315 | b315;
  assign c316 = (a315 & b315) | (a315 & c315) | (b315 & c315);
  wire c_sub316;
  assign c_sub316 = (a315 & b_inv315) | (a315 & c315) | (b_inv315 & c315);
  wire s316, sub316, and316, or316;
  wire b_inv316;
  assign b_inv316 = ~b316;
  assign s316  = a316 ^ b316 ^ c316;
  assign sub316 = a316 ^ b_inv316 ^ c316;
  assign and316 = a316 & b316;
  assign or316  = a316 | b316;
  assign c317 = (a316 & b316) | (a316 & c316) | (b316 & c316);
  wire c_sub317;
  assign c_sub317 = (a316 & b_inv316) | (a316 & c316) | (b_inv316 & c316);
  wire s317, sub317, and317, or317;
  wire b_inv317;
  assign b_inv317 = ~b317;
  assign s317  = a317 ^ b317 ^ c317;
  assign sub317 = a317 ^ b_inv317 ^ c317;
  assign and317 = a317 & b317;
  assign or317  = a317 | b317;
  assign c318 = (a317 & b317) | (a317 & c317) | (b317 & c317);
  wire c_sub318;
  assign c_sub318 = (a317 & b_inv317) | (a317 & c317) | (b_inv317 & c317);
  wire s318, sub318, and318, or318;
  wire b_inv318;
  assign b_inv318 = ~b318;
  assign s318  = a318 ^ b318 ^ c318;
  assign sub318 = a318 ^ b_inv318 ^ c318;
  assign and318 = a318 & b318;
  assign or318  = a318 | b318;
  assign c319 = (a318 & b318) | (a318 & c318) | (b318 & c318);
  wire c_sub319;
  assign c_sub319 = (a318 & b_inv318) | (a318 & c318) | (b_inv318 & c318);
  wire s319, sub319, and319, or319;
  wire b_inv319;
  assign b_inv319 = ~b319;
  assign s319  = a319 ^ b319 ^ c319;
  assign sub319 = a319 ^ b_inv319 ^ c319;
  assign and319 = a319 & b319;
  assign or319  = a319 | b319;
  assign c320 = (a319 & b319) | (a319 & c319) | (b319 & c319);
  wire c_sub320;
  assign c_sub320 = (a319 & b_inv319) | (a319 & c319) | (b_inv319 & c319);
  wire s320, sub320, and320, or320;
  wire b_inv320;
  assign b_inv320 = ~b320;
  assign s320  = a320 ^ b320 ^ c320;
  assign sub320 = a320 ^ b_inv320 ^ c320;
  assign and320 = a320 & b320;
  assign or320  = a320 | b320;
  assign c321 = (a320 & b320) | (a320 & c320) | (b320 & c320);
  wire c_sub321;
  assign c_sub321 = (a320 & b_inv320) | (a320 & c320) | (b_inv320 & c320);
  wire s321, sub321, and321, or321;
  wire b_inv321;
  assign b_inv321 = ~b321;
  assign s321  = a321 ^ b321 ^ c321;
  assign sub321 = a321 ^ b_inv321 ^ c321;
  assign and321 = a321 & b321;
  assign or321  = a321 | b321;
  assign c322 = (a321 & b321) | (a321 & c321) | (b321 & c321);
  wire c_sub322;
  assign c_sub322 = (a321 & b_inv321) | (a321 & c321) | (b_inv321 & c321);
  wire s322, sub322, and322, or322;
  wire b_inv322;
  assign b_inv322 = ~b322;
  assign s322  = a322 ^ b322 ^ c322;
  assign sub322 = a322 ^ b_inv322 ^ c322;
  assign and322 = a322 & b322;
  assign or322  = a322 | b322;
  assign c323 = (a322 & b322) | (a322 & c322) | (b322 & c322);
  wire c_sub323;
  assign c_sub323 = (a322 & b_inv322) | (a322 & c322) | (b_inv322 & c322);
  wire s323, sub323, and323, or323;
  wire b_inv323;
  assign b_inv323 = ~b323;
  assign s323  = a323 ^ b323 ^ c323;
  assign sub323 = a323 ^ b_inv323 ^ c323;
  assign and323 = a323 & b323;
  assign or323  = a323 | b323;
  assign c324 = (a323 & b323) | (a323 & c323) | (b323 & c323);
  wire c_sub324;
  assign c_sub324 = (a323 & b_inv323) | (a323 & c323) | (b_inv323 & c323);
  wire s324, sub324, and324, or324;
  wire b_inv324;
  assign b_inv324 = ~b324;
  assign s324  = a324 ^ b324 ^ c324;
  assign sub324 = a324 ^ b_inv324 ^ c324;
  assign and324 = a324 & b324;
  assign or324  = a324 | b324;
  assign c325 = (a324 & b324) | (a324 & c324) | (b324 & c324);
  wire c_sub325;
  assign c_sub325 = (a324 & b_inv324) | (a324 & c324) | (b_inv324 & c324);
  wire s325, sub325, and325, or325;
  wire b_inv325;
  assign b_inv325 = ~b325;
  assign s325  = a325 ^ b325 ^ c325;
  assign sub325 = a325 ^ b_inv325 ^ c325;
  assign and325 = a325 & b325;
  assign or325  = a325 | b325;
  assign c326 = (a325 & b325) | (a325 & c325) | (b325 & c325);
  wire c_sub326;
  assign c_sub326 = (a325 & b_inv325) | (a325 & c325) | (b_inv325 & c325);
  wire s326, sub326, and326, or326;
  wire b_inv326;
  assign b_inv326 = ~b326;
  assign s326  = a326 ^ b326 ^ c326;
  assign sub326 = a326 ^ b_inv326 ^ c326;
  assign and326 = a326 & b326;
  assign or326  = a326 | b326;
  assign c327 = (a326 & b326) | (a326 & c326) | (b326 & c326);
  wire c_sub327;
  assign c_sub327 = (a326 & b_inv326) | (a326 & c326) | (b_inv326 & c326);
  wire s327, sub327, and327, or327;
  wire b_inv327;
  assign b_inv327 = ~b327;
  assign s327  = a327 ^ b327 ^ c327;
  assign sub327 = a327 ^ b_inv327 ^ c327;
  assign and327 = a327 & b327;
  assign or327  = a327 | b327;
  assign c328 = (a327 & b327) | (a327 & c327) | (b327 & c327);
  wire c_sub328;
  assign c_sub328 = (a327 & b_inv327) | (a327 & c327) | (b_inv327 & c327);
  wire s328, sub328, and328, or328;
  wire b_inv328;
  assign b_inv328 = ~b328;
  assign s328  = a328 ^ b328 ^ c328;
  assign sub328 = a328 ^ b_inv328 ^ c328;
  assign and328 = a328 & b328;
  assign or328  = a328 | b328;
  assign c329 = (a328 & b328) | (a328 & c328) | (b328 & c328);
  wire c_sub329;
  assign c_sub329 = (a328 & b_inv328) | (a328 & c328) | (b_inv328 & c328);
  wire s329, sub329, and329, or329;
  wire b_inv329;
  assign b_inv329 = ~b329;
  assign s329  = a329 ^ b329 ^ c329;
  assign sub329 = a329 ^ b_inv329 ^ c329;
  assign and329 = a329 & b329;
  assign or329  = a329 | b329;
  assign c330 = (a329 & b329) | (a329 & c329) | (b329 & c329);
  wire c_sub330;
  assign c_sub330 = (a329 & b_inv329) | (a329 & c329) | (b_inv329 & c329);
  wire s330, sub330, and330, or330;
  wire b_inv330;
  assign b_inv330 = ~b330;
  assign s330  = a330 ^ b330 ^ c330;
  assign sub330 = a330 ^ b_inv330 ^ c330;
  assign and330 = a330 & b330;
  assign or330  = a330 | b330;
  assign c331 = (a330 & b330) | (a330 & c330) | (b330 & c330);
  wire c_sub331;
  assign c_sub331 = (a330 & b_inv330) | (a330 & c330) | (b_inv330 & c330);
  wire s331, sub331, and331, or331;
  wire b_inv331;
  assign b_inv331 = ~b331;
  assign s331  = a331 ^ b331 ^ c331;
  assign sub331 = a331 ^ b_inv331 ^ c331;
  assign and331 = a331 & b331;
  assign or331  = a331 | b331;
  assign c332 = (a331 & b331) | (a331 & c331) | (b331 & c331);
  wire c_sub332;
  assign c_sub332 = (a331 & b_inv331) | (a331 & c331) | (b_inv331 & c331);
  wire s332, sub332, and332, or332;
  wire b_inv332;
  assign b_inv332 = ~b332;
  assign s332  = a332 ^ b332 ^ c332;
  assign sub332 = a332 ^ b_inv332 ^ c332;
  assign and332 = a332 & b332;
  assign or332  = a332 | b332;
  assign c333 = (a332 & b332) | (a332 & c332) | (b332 & c332);
  wire c_sub333;
  assign c_sub333 = (a332 & b_inv332) | (a332 & c332) | (b_inv332 & c332);
  wire s333, sub333, and333, or333;
  wire b_inv333;
  assign b_inv333 = ~b333;
  assign s333  = a333 ^ b333 ^ c333;
  assign sub333 = a333 ^ b_inv333 ^ c333;
  assign and333 = a333 & b333;
  assign or333  = a333 | b333;
  assign c334 = (a333 & b333) | (a333 & c333) | (b333 & c333);
  wire c_sub334;
  assign c_sub334 = (a333 & b_inv333) | (a333 & c333) | (b_inv333 & c333);
  wire s334, sub334, and334, or334;
  wire b_inv334;
  assign b_inv334 = ~b334;
  assign s334  = a334 ^ b334 ^ c334;
  assign sub334 = a334 ^ b_inv334 ^ c334;
  assign and334 = a334 & b334;
  assign or334  = a334 | b334;
  assign c335 = (a334 & b334) | (a334 & c334) | (b334 & c334);
  wire c_sub335;
  assign c_sub335 = (a334 & b_inv334) | (a334 & c334) | (b_inv334 & c334);
  wire s335, sub335, and335, or335;
  wire b_inv335;
  assign b_inv335 = ~b335;
  assign s335  = a335 ^ b335 ^ c335;
  assign sub335 = a335 ^ b_inv335 ^ c335;
  assign and335 = a335 & b335;
  assign or335  = a335 | b335;
  assign c336 = (a335 & b335) | (a335 & c335) | (b335 & c335);
  wire c_sub336;
  assign c_sub336 = (a335 & b_inv335) | (a335 & c335) | (b_inv335 & c335);
  wire s336, sub336, and336, or336;
  wire b_inv336;
  assign b_inv336 = ~b336;
  assign s336  = a336 ^ b336 ^ c336;
  assign sub336 = a336 ^ b_inv336 ^ c336;
  assign and336 = a336 & b336;
  assign or336  = a336 | b336;
  assign c337 = (a336 & b336) | (a336 & c336) | (b336 & c336);
  wire c_sub337;
  assign c_sub337 = (a336 & b_inv336) | (a336 & c336) | (b_inv336 & c336);
  wire s337, sub337, and337, or337;
  wire b_inv337;
  assign b_inv337 = ~b337;
  assign s337  = a337 ^ b337 ^ c337;
  assign sub337 = a337 ^ b_inv337 ^ c337;
  assign and337 = a337 & b337;
  assign or337  = a337 | b337;
  assign c338 = (a337 & b337) | (a337 & c337) | (b337 & c337);
  wire c_sub338;
  assign c_sub338 = (a337 & b_inv337) | (a337 & c337) | (b_inv337 & c337);
  wire s338, sub338, and338, or338;
  wire b_inv338;
  assign b_inv338 = ~b338;
  assign s338  = a338 ^ b338 ^ c338;
  assign sub338 = a338 ^ b_inv338 ^ c338;
  assign and338 = a338 & b338;
  assign or338  = a338 | b338;
  assign c339 = (a338 & b338) | (a338 & c338) | (b338 & c338);
  wire c_sub339;
  assign c_sub339 = (a338 & b_inv338) | (a338 & c338) | (b_inv338 & c338);
  wire s339, sub339, and339, or339;
  wire b_inv339;
  assign b_inv339 = ~b339;
  assign s339  = a339 ^ b339 ^ c339;
  assign sub339 = a339 ^ b_inv339 ^ c339;
  assign and339 = a339 & b339;
  assign or339  = a339 | b339;
  assign c340 = (a339 & b339) | (a339 & c339) | (b339 & c339);
  wire c_sub340;
  assign c_sub340 = (a339 & b_inv339) | (a339 & c339) | (b_inv339 & c339);
  wire s340, sub340, and340, or340;
  wire b_inv340;
  assign b_inv340 = ~b340;
  assign s340  = a340 ^ b340 ^ c340;
  assign sub340 = a340 ^ b_inv340 ^ c340;
  assign and340 = a340 & b340;
  assign or340  = a340 | b340;
  assign c341 = (a340 & b340) | (a340 & c340) | (b340 & c340);
  wire c_sub341;
  assign c_sub341 = (a340 & b_inv340) | (a340 & c340) | (b_inv340 & c340);
  wire s341, sub341, and341, or341;
  wire b_inv341;
  assign b_inv341 = ~b341;
  assign s341  = a341 ^ b341 ^ c341;
  assign sub341 = a341 ^ b_inv341 ^ c341;
  assign and341 = a341 & b341;
  assign or341  = a341 | b341;
  assign c342 = (a341 & b341) | (a341 & c341) | (b341 & c341);
  wire c_sub342;
  assign c_sub342 = (a341 & b_inv341) | (a341 & c341) | (b_inv341 & c341);
  wire s342, sub342, and342, or342;
  wire b_inv342;
  assign b_inv342 = ~b342;
  assign s342  = a342 ^ b342 ^ c342;
  assign sub342 = a342 ^ b_inv342 ^ c342;
  assign and342 = a342 & b342;
  assign or342  = a342 | b342;
  assign c343 = (a342 & b342) | (a342 & c342) | (b342 & c342);
  wire c_sub343;
  assign c_sub343 = (a342 & b_inv342) | (a342 & c342) | (b_inv342 & c342);
  wire s343, sub343, and343, or343;
  wire b_inv343;
  assign b_inv343 = ~b343;
  assign s343  = a343 ^ b343 ^ c343;
  assign sub343 = a343 ^ b_inv343 ^ c343;
  assign and343 = a343 & b343;
  assign or343  = a343 | b343;
  assign c344 = (a343 & b343) | (a343 & c343) | (b343 & c343);
  wire c_sub344;
  assign c_sub344 = (a343 & b_inv343) | (a343 & c343) | (b_inv343 & c343);
  wire s344, sub344, and344, or344;
  wire b_inv344;
  assign b_inv344 = ~b344;
  assign s344  = a344 ^ b344 ^ c344;
  assign sub344 = a344 ^ b_inv344 ^ c344;
  assign and344 = a344 & b344;
  assign or344  = a344 | b344;
  assign c345 = (a344 & b344) | (a344 & c344) | (b344 & c344);
  wire c_sub345;
  assign c_sub345 = (a344 & b_inv344) | (a344 & c344) | (b_inv344 & c344);
  wire s345, sub345, and345, or345;
  wire b_inv345;
  assign b_inv345 = ~b345;
  assign s345  = a345 ^ b345 ^ c345;
  assign sub345 = a345 ^ b_inv345 ^ c345;
  assign and345 = a345 & b345;
  assign or345  = a345 | b345;
  assign c346 = (a345 & b345) | (a345 & c345) | (b345 & c345);
  wire c_sub346;
  assign c_sub346 = (a345 & b_inv345) | (a345 & c345) | (b_inv345 & c345);
  wire s346, sub346, and346, or346;
  wire b_inv346;
  assign b_inv346 = ~b346;
  assign s346  = a346 ^ b346 ^ c346;
  assign sub346 = a346 ^ b_inv346 ^ c346;
  assign and346 = a346 & b346;
  assign or346  = a346 | b346;
  assign c347 = (a346 & b346) | (a346 & c346) | (b346 & c346);
  wire c_sub347;
  assign c_sub347 = (a346 & b_inv346) | (a346 & c346) | (b_inv346 & c346);
  wire s347, sub347, and347, or347;
  wire b_inv347;
  assign b_inv347 = ~b347;
  assign s347  = a347 ^ b347 ^ c347;
  assign sub347 = a347 ^ b_inv347 ^ c347;
  assign and347 = a347 & b347;
  assign or347  = a347 | b347;
  assign c348 = (a347 & b347) | (a347 & c347) | (b347 & c347);
  wire c_sub348;
  assign c_sub348 = (a347 & b_inv347) | (a347 & c347) | (b_inv347 & c347);
  wire s348, sub348, and348, or348;
  wire b_inv348;
  assign b_inv348 = ~b348;
  assign s348  = a348 ^ b348 ^ c348;
  assign sub348 = a348 ^ b_inv348 ^ c348;
  assign and348 = a348 & b348;
  assign or348  = a348 | b348;
  assign c349 = (a348 & b348) | (a348 & c348) | (b348 & c348);
  wire c_sub349;
  assign c_sub349 = (a348 & b_inv348) | (a348 & c348) | (b_inv348 & c348);
  wire s349, sub349, and349, or349;
  wire b_inv349;
  assign b_inv349 = ~b349;
  assign s349  = a349 ^ b349 ^ c349;
  assign sub349 = a349 ^ b_inv349 ^ c349;
  assign and349 = a349 & b349;
  assign or349  = a349 | b349;
  assign c350 = (a349 & b349) | (a349 & c349) | (b349 & c349);
  wire c_sub350;
  assign c_sub350 = (a349 & b_inv349) | (a349 & c349) | (b_inv349 & c349);
  wire s350, sub350, and350, or350;
  wire b_inv350;
  assign b_inv350 = ~b350;
  assign s350  = a350 ^ b350 ^ c350;
  assign sub350 = a350 ^ b_inv350 ^ c350;
  assign and350 = a350 & b350;
  assign or350  = a350 | b350;
  assign c351 = (a350 & b350) | (a350 & c350) | (b350 & c350);
  wire c_sub351;
  assign c_sub351 = (a350 & b_inv350) | (a350 & c350) | (b_inv350 & c350);
  wire s351, sub351, and351, or351;
  wire b_inv351;
  assign b_inv351 = ~b351;
  assign s351  = a351 ^ b351 ^ c351;
  assign sub351 = a351 ^ b_inv351 ^ c351;
  assign and351 = a351 & b351;
  assign or351  = a351 | b351;
  assign c352 = (a351 & b351) | (a351 & c351) | (b351 & c351);
  wire c_sub352;
  assign c_sub352 = (a351 & b_inv351) | (a351 & c351) | (b_inv351 & c351);
  wire s352, sub352, and352, or352;
  wire b_inv352;
  assign b_inv352 = ~b352;
  assign s352  = a352 ^ b352 ^ c352;
  assign sub352 = a352 ^ b_inv352 ^ c352;
  assign and352 = a352 & b352;
  assign or352  = a352 | b352;
  assign c353 = (a352 & b352) | (a352 & c352) | (b352 & c352);
  wire c_sub353;
  assign c_sub353 = (a352 & b_inv352) | (a352 & c352) | (b_inv352 & c352);
  wire s353, sub353, and353, or353;
  wire b_inv353;
  assign b_inv353 = ~b353;
  assign s353  = a353 ^ b353 ^ c353;
  assign sub353 = a353 ^ b_inv353 ^ c353;
  assign and353 = a353 & b353;
  assign or353  = a353 | b353;
  assign c354 = (a353 & b353) | (a353 & c353) | (b353 & c353);
  wire c_sub354;
  assign c_sub354 = (a353 & b_inv353) | (a353 & c353) | (b_inv353 & c353);
  wire s354, sub354, and354, or354;
  wire b_inv354;
  assign b_inv354 = ~b354;
  assign s354  = a354 ^ b354 ^ c354;
  assign sub354 = a354 ^ b_inv354 ^ c354;
  assign and354 = a354 & b354;
  assign or354  = a354 | b354;
  assign c355 = (a354 & b354) | (a354 & c354) | (b354 & c354);
  wire c_sub355;
  assign c_sub355 = (a354 & b_inv354) | (a354 & c354) | (b_inv354 & c354);
  wire s355, sub355, and355, or355;
  wire b_inv355;
  assign b_inv355 = ~b355;
  assign s355  = a355 ^ b355 ^ c355;
  assign sub355 = a355 ^ b_inv355 ^ c355;
  assign and355 = a355 & b355;
  assign or355  = a355 | b355;
  assign c356 = (a355 & b355) | (a355 & c355) | (b355 & c355);
  wire c_sub356;
  assign c_sub356 = (a355 & b_inv355) | (a355 & c355) | (b_inv355 & c355);
  wire s356, sub356, and356, or356;
  wire b_inv356;
  assign b_inv356 = ~b356;
  assign s356  = a356 ^ b356 ^ c356;
  assign sub356 = a356 ^ b_inv356 ^ c356;
  assign and356 = a356 & b356;
  assign or356  = a356 | b356;
  assign c357 = (a356 & b356) | (a356 & c356) | (b356 & c356);
  wire c_sub357;
  assign c_sub357 = (a356 & b_inv356) | (a356 & c356) | (b_inv356 & c356);
  wire s357, sub357, and357, or357;
  wire b_inv357;
  assign b_inv357 = ~b357;
  assign s357  = a357 ^ b357 ^ c357;
  assign sub357 = a357 ^ b_inv357 ^ c357;
  assign and357 = a357 & b357;
  assign or357  = a357 | b357;
  assign c358 = (a357 & b357) | (a357 & c357) | (b357 & c357);
  wire c_sub358;
  assign c_sub358 = (a357 & b_inv357) | (a357 & c357) | (b_inv357 & c357);
  wire s358, sub358, and358, or358;
  wire b_inv358;
  assign b_inv358 = ~b358;
  assign s358  = a358 ^ b358 ^ c358;
  assign sub358 = a358 ^ b_inv358 ^ c358;
  assign and358 = a358 & b358;
  assign or358  = a358 | b358;
  assign c359 = (a358 & b358) | (a358 & c358) | (b358 & c358);
  wire c_sub359;
  assign c_sub359 = (a358 & b_inv358) | (a358 & c358) | (b_inv358 & c358);
  wire s359, sub359, and359, or359;
  wire b_inv359;
  assign b_inv359 = ~b359;
  assign s359  = a359 ^ b359 ^ c359;
  assign sub359 = a359 ^ b_inv359 ^ c359;
  assign and359 = a359 & b359;
  assign or359  = a359 | b359;
  assign c360 = (a359 & b359) | (a359 & c359) | (b359 & c359);
  wire c_sub360;
  assign c_sub360 = (a359 & b_inv359) | (a359 & c359) | (b_inv359 & c359);
  wire s360, sub360, and360, or360;
  wire b_inv360;
  assign b_inv360 = ~b360;
  assign s360  = a360 ^ b360 ^ c360;
  assign sub360 = a360 ^ b_inv360 ^ c360;
  assign and360 = a360 & b360;
  assign or360  = a360 | b360;
  assign c361 = (a360 & b360) | (a360 & c360) | (b360 & c360);
  wire c_sub361;
  assign c_sub361 = (a360 & b_inv360) | (a360 & c360) | (b_inv360 & c360);
  wire s361, sub361, and361, or361;
  wire b_inv361;
  assign b_inv361 = ~b361;
  assign s361  = a361 ^ b361 ^ c361;
  assign sub361 = a361 ^ b_inv361 ^ c361;
  assign and361 = a361 & b361;
  assign or361  = a361 | b361;
  assign c362 = (a361 & b361) | (a361 & c361) | (b361 & c361);
  wire c_sub362;
  assign c_sub362 = (a361 & b_inv361) | (a361 & c361) | (b_inv361 & c361);
  wire s362, sub362, and362, or362;
  wire b_inv362;
  assign b_inv362 = ~b362;
  assign s362  = a362 ^ b362 ^ c362;
  assign sub362 = a362 ^ b_inv362 ^ c362;
  assign and362 = a362 & b362;
  assign or362  = a362 | b362;
  assign c363 = (a362 & b362) | (a362 & c362) | (b362 & c362);
  wire c_sub363;
  assign c_sub363 = (a362 & b_inv362) | (a362 & c362) | (b_inv362 & c362);
  wire s363, sub363, and363, or363;
  wire b_inv363;
  assign b_inv363 = ~b363;
  assign s363  = a363 ^ b363 ^ c363;
  assign sub363 = a363 ^ b_inv363 ^ c363;
  assign and363 = a363 & b363;
  assign or363  = a363 | b363;
  assign c364 = (a363 & b363) | (a363 & c363) | (b363 & c363);
  wire c_sub364;
  assign c_sub364 = (a363 & b_inv363) | (a363 & c363) | (b_inv363 & c363);
  wire s364, sub364, and364, or364;
  wire b_inv364;
  assign b_inv364 = ~b364;
  assign s364  = a364 ^ b364 ^ c364;
  assign sub364 = a364 ^ b_inv364 ^ c364;
  assign and364 = a364 & b364;
  assign or364  = a364 | b364;
  assign c365 = (a364 & b364) | (a364 & c364) | (b364 & c364);
  wire c_sub365;
  assign c_sub365 = (a364 & b_inv364) | (a364 & c364) | (b_inv364 & c364);
  wire s365, sub365, and365, or365;
  wire b_inv365;
  assign b_inv365 = ~b365;
  assign s365  = a365 ^ b365 ^ c365;
  assign sub365 = a365 ^ b_inv365 ^ c365;
  assign and365 = a365 & b365;
  assign or365  = a365 | b365;
  assign c366 = (a365 & b365) | (a365 & c365) | (b365 & c365);
  wire c_sub366;
  assign c_sub366 = (a365 & b_inv365) | (a365 & c365) | (b_inv365 & c365);
  wire s366, sub366, and366, or366;
  wire b_inv366;
  assign b_inv366 = ~b366;
  assign s366  = a366 ^ b366 ^ c366;
  assign sub366 = a366 ^ b_inv366 ^ c366;
  assign and366 = a366 & b366;
  assign or366  = a366 | b366;
  assign c367 = (a366 & b366) | (a366 & c366) | (b366 & c366);
  wire c_sub367;
  assign c_sub367 = (a366 & b_inv366) | (a366 & c366) | (b_inv366 & c366);
  wire s367, sub367, and367, or367;
  wire b_inv367;
  assign b_inv367 = ~b367;
  assign s367  = a367 ^ b367 ^ c367;
  assign sub367 = a367 ^ b_inv367 ^ c367;
  assign and367 = a367 & b367;
  assign or367  = a367 | b367;
  assign c368 = (a367 & b367) | (a367 & c367) | (b367 & c367);
  wire c_sub368;
  assign c_sub368 = (a367 & b_inv367) | (a367 & c367) | (b_inv367 & c367);
  wire s368, sub368, and368, or368;
  wire b_inv368;
  assign b_inv368 = ~b368;
  assign s368  = a368 ^ b368 ^ c368;
  assign sub368 = a368 ^ b_inv368 ^ c368;
  assign and368 = a368 & b368;
  assign or368  = a368 | b368;
  assign c369 = (a368 & b368) | (a368 & c368) | (b368 & c368);
  wire c_sub369;
  assign c_sub369 = (a368 & b_inv368) | (a368 & c368) | (b_inv368 & c368);
  wire s369, sub369, and369, or369;
  wire b_inv369;
  assign b_inv369 = ~b369;
  assign s369  = a369 ^ b369 ^ c369;
  assign sub369 = a369 ^ b_inv369 ^ c369;
  assign and369 = a369 & b369;
  assign or369  = a369 | b369;
  assign c370 = (a369 & b369) | (a369 & c369) | (b369 & c369);
  wire c_sub370;
  assign c_sub370 = (a369 & b_inv369) | (a369 & c369) | (b_inv369 & c369);
  wire s370, sub370, and370, or370;
  wire b_inv370;
  assign b_inv370 = ~b370;
  assign s370  = a370 ^ b370 ^ c370;
  assign sub370 = a370 ^ b_inv370 ^ c370;
  assign and370 = a370 & b370;
  assign or370  = a370 | b370;
  assign c371 = (a370 & b370) | (a370 & c370) | (b370 & c370);
  wire c_sub371;
  assign c_sub371 = (a370 & b_inv370) | (a370 & c370) | (b_inv370 & c370);
  wire s371, sub371, and371, or371;
  wire b_inv371;
  assign b_inv371 = ~b371;
  assign s371  = a371 ^ b371 ^ c371;
  assign sub371 = a371 ^ b_inv371 ^ c371;
  assign and371 = a371 & b371;
  assign or371  = a371 | b371;
  assign c372 = (a371 & b371) | (a371 & c371) | (b371 & c371);
  wire c_sub372;
  assign c_sub372 = (a371 & b_inv371) | (a371 & c371) | (b_inv371 & c371);
  wire s372, sub372, and372, or372;
  wire b_inv372;
  assign b_inv372 = ~b372;
  assign s372  = a372 ^ b372 ^ c372;
  assign sub372 = a372 ^ b_inv372 ^ c372;
  assign and372 = a372 & b372;
  assign or372  = a372 | b372;
  assign c373 = (a372 & b372) | (a372 & c372) | (b372 & c372);
  wire c_sub373;
  assign c_sub373 = (a372 & b_inv372) | (a372 & c372) | (b_inv372 & c372);
  wire s373, sub373, and373, or373;
  wire b_inv373;
  assign b_inv373 = ~b373;
  assign s373  = a373 ^ b373 ^ c373;
  assign sub373 = a373 ^ b_inv373 ^ c373;
  assign and373 = a373 & b373;
  assign or373  = a373 | b373;
  assign c374 = (a373 & b373) | (a373 & c373) | (b373 & c373);
  wire c_sub374;
  assign c_sub374 = (a373 & b_inv373) | (a373 & c373) | (b_inv373 & c373);
  wire s374, sub374, and374, or374;
  wire b_inv374;
  assign b_inv374 = ~b374;
  assign s374  = a374 ^ b374 ^ c374;
  assign sub374 = a374 ^ b_inv374 ^ c374;
  assign and374 = a374 & b374;
  assign or374  = a374 | b374;
  assign c375 = (a374 & b374) | (a374 & c374) | (b374 & c374);
  wire c_sub375;
  assign c_sub375 = (a374 & b_inv374) | (a374 & c374) | (b_inv374 & c374);
  wire s375, sub375, and375, or375;
  wire b_inv375;
  assign b_inv375 = ~b375;
  assign s375  = a375 ^ b375 ^ c375;
  assign sub375 = a375 ^ b_inv375 ^ c375;
  assign and375 = a375 & b375;
  assign or375  = a375 | b375;
  assign c376 = (a375 & b375) | (a375 & c375) | (b375 & c375);
  wire c_sub376;
  assign c_sub376 = (a375 & b_inv375) | (a375 & c375) | (b_inv375 & c375);
  wire s376, sub376, and376, or376;
  wire b_inv376;
  assign b_inv376 = ~b376;
  assign s376  = a376 ^ b376 ^ c376;
  assign sub376 = a376 ^ b_inv376 ^ c376;
  assign and376 = a376 & b376;
  assign or376  = a376 | b376;
  assign c377 = (a376 & b376) | (a376 & c376) | (b376 & c376);
  wire c_sub377;
  assign c_sub377 = (a376 & b_inv376) | (a376 & c376) | (b_inv376 & c376);
  wire s377, sub377, and377, or377;
  wire b_inv377;
  assign b_inv377 = ~b377;
  assign s377  = a377 ^ b377 ^ c377;
  assign sub377 = a377 ^ b_inv377 ^ c377;
  assign and377 = a377 & b377;
  assign or377  = a377 | b377;
  assign c378 = (a377 & b377) | (a377 & c377) | (b377 & c377);
  wire c_sub378;
  assign c_sub378 = (a377 & b_inv377) | (a377 & c377) | (b_inv377 & c377);
  wire s378, sub378, and378, or378;
  wire b_inv378;
  assign b_inv378 = ~b378;
  assign s378  = a378 ^ b378 ^ c378;
  assign sub378 = a378 ^ b_inv378 ^ c378;
  assign and378 = a378 & b378;
  assign or378  = a378 | b378;
  assign c379 = (a378 & b378) | (a378 & c378) | (b378 & c378);
  wire c_sub379;
  assign c_sub379 = (a378 & b_inv378) | (a378 & c378) | (b_inv378 & c378);
  wire s379, sub379, and379, or379;
  wire b_inv379;
  assign b_inv379 = ~b379;
  assign s379  = a379 ^ b379 ^ c379;
  assign sub379 = a379 ^ b_inv379 ^ c379;
  assign and379 = a379 & b379;
  assign or379  = a379 | b379;
  assign c380 = (a379 & b379) | (a379 & c379) | (b379 & c379);
  wire c_sub380;
  assign c_sub380 = (a379 & b_inv379) | (a379 & c379) | (b_inv379 & c379);
  wire s380, sub380, and380, or380;
  wire b_inv380;
  assign b_inv380 = ~b380;
  assign s380  = a380 ^ b380 ^ c380;
  assign sub380 = a380 ^ b_inv380 ^ c380;
  assign and380 = a380 & b380;
  assign or380  = a380 | b380;
  assign c381 = (a380 & b380) | (a380 & c380) | (b380 & c380);
  wire c_sub381;
  assign c_sub381 = (a380 & b_inv380) | (a380 & c380) | (b_inv380 & c380);
  wire s381, sub381, and381, or381;
  wire b_inv381;
  assign b_inv381 = ~b381;
  assign s381  = a381 ^ b381 ^ c381;
  assign sub381 = a381 ^ b_inv381 ^ c381;
  assign and381 = a381 & b381;
  assign or381  = a381 | b381;
  assign c382 = (a381 & b381) | (a381 & c381) | (b381 & c381);
  wire c_sub382;
  assign c_sub382 = (a381 & b_inv381) | (a381 & c381) | (b_inv381 & c381);
  wire s382, sub382, and382, or382;
  wire b_inv382;
  assign b_inv382 = ~b382;
  assign s382  = a382 ^ b382 ^ c382;
  assign sub382 = a382 ^ b_inv382 ^ c382;
  assign and382 = a382 & b382;
  assign or382  = a382 | b382;
  assign c383 = (a382 & b382) | (a382 & c382) | (b382 & c382);
  wire c_sub383;
  assign c_sub383 = (a382 & b_inv382) | (a382 & c382) | (b_inv382 & c382);
  wire s383, sub383, and383, or383;
  wire b_inv383;
  assign b_inv383 = ~b383;
  assign s383  = a383 ^ b383 ^ c383;
  assign sub383 = a383 ^ b_inv383 ^ c383;
  assign and383 = a383 & b383;
  assign or383  = a383 | b383;
  assign c384 = (a383 & b383) | (a383 & c383) | (b383 & c383);
  wire c_sub384;
  assign c_sub384 = (a383 & b_inv383) | (a383 & c383) | (b_inv383 & c383);
  wire s384, sub384, and384, or384;
  wire b_inv384;
  assign b_inv384 = ~b384;
  assign s384  = a384 ^ b384 ^ c384;
  assign sub384 = a384 ^ b_inv384 ^ c384;
  assign and384 = a384 & b384;
  assign or384  = a384 | b384;
  assign c385 = (a384 & b384) | (a384 & c384) | (b384 & c384);
  wire c_sub385;
  assign c_sub385 = (a384 & b_inv384) | (a384 & c384) | (b_inv384 & c384);
  wire s385, sub385, and385, or385;
  wire b_inv385;
  assign b_inv385 = ~b385;
  assign s385  = a385 ^ b385 ^ c385;
  assign sub385 = a385 ^ b_inv385 ^ c385;
  assign and385 = a385 & b385;
  assign or385  = a385 | b385;
  assign c386 = (a385 & b385) | (a385 & c385) | (b385 & c385);
  wire c_sub386;
  assign c_sub386 = (a385 & b_inv385) | (a385 & c385) | (b_inv385 & c385);
  wire s386, sub386, and386, or386;
  wire b_inv386;
  assign b_inv386 = ~b386;
  assign s386  = a386 ^ b386 ^ c386;
  assign sub386 = a386 ^ b_inv386 ^ c386;
  assign and386 = a386 & b386;
  assign or386  = a386 | b386;
  assign c387 = (a386 & b386) | (a386 & c386) | (b386 & c386);
  wire c_sub387;
  assign c_sub387 = (a386 & b_inv386) | (a386 & c386) | (b_inv386 & c386);
  wire s387, sub387, and387, or387;
  wire b_inv387;
  assign b_inv387 = ~b387;
  assign s387  = a387 ^ b387 ^ c387;
  assign sub387 = a387 ^ b_inv387 ^ c387;
  assign and387 = a387 & b387;
  assign or387  = a387 | b387;
  assign c388 = (a387 & b387) | (a387 & c387) | (b387 & c387);
  wire c_sub388;
  assign c_sub388 = (a387 & b_inv387) | (a387 & c387) | (b_inv387 & c387);
  wire s388, sub388, and388, or388;
  wire b_inv388;
  assign b_inv388 = ~b388;
  assign s388  = a388 ^ b388 ^ c388;
  assign sub388 = a388 ^ b_inv388 ^ c388;
  assign and388 = a388 & b388;
  assign or388  = a388 | b388;
  assign c389 = (a388 & b388) | (a388 & c388) | (b388 & c388);
  wire c_sub389;
  assign c_sub389 = (a388 & b_inv388) | (a388 & c388) | (b_inv388 & c388);
  wire s389, sub389, and389, or389;
  wire b_inv389;
  assign b_inv389 = ~b389;
  assign s389  = a389 ^ b389 ^ c389;
  assign sub389 = a389 ^ b_inv389 ^ c389;
  assign and389 = a389 & b389;
  assign or389  = a389 | b389;
  assign c390 = (a389 & b389) | (a389 & c389) | (b389 & c389);
  wire c_sub390;
  assign c_sub390 = (a389 & b_inv389) | (a389 & c389) | (b_inv389 & c389);
  wire s390, sub390, and390, or390;
  wire b_inv390;
  assign b_inv390 = ~b390;
  assign s390  = a390 ^ b390 ^ c390;
  assign sub390 = a390 ^ b_inv390 ^ c390;
  assign and390 = a390 & b390;
  assign or390  = a390 | b390;
  assign c391 = (a390 & b390) | (a390 & c390) | (b390 & c390);
  wire c_sub391;
  assign c_sub391 = (a390 & b_inv390) | (a390 & c390) | (b_inv390 & c390);
  wire s391, sub391, and391, or391;
  wire b_inv391;
  assign b_inv391 = ~b391;
  assign s391  = a391 ^ b391 ^ c391;
  assign sub391 = a391 ^ b_inv391 ^ c391;
  assign and391 = a391 & b391;
  assign or391  = a391 | b391;
  assign c392 = (a391 & b391) | (a391 & c391) | (b391 & c391);
  wire c_sub392;
  assign c_sub392 = (a391 & b_inv391) | (a391 & c391) | (b_inv391 & c391);
  wire s392, sub392, and392, or392;
  wire b_inv392;
  assign b_inv392 = ~b392;
  assign s392  = a392 ^ b392 ^ c392;
  assign sub392 = a392 ^ b_inv392 ^ c392;
  assign and392 = a392 & b392;
  assign or392  = a392 | b392;
  assign c393 = (a392 & b392) | (a392 & c392) | (b392 & c392);
  wire c_sub393;
  assign c_sub393 = (a392 & b_inv392) | (a392 & c392) | (b_inv392 & c392);
  wire s393, sub393, and393, or393;
  wire b_inv393;
  assign b_inv393 = ~b393;
  assign s393  = a393 ^ b393 ^ c393;
  assign sub393 = a393 ^ b_inv393 ^ c393;
  assign and393 = a393 & b393;
  assign or393  = a393 | b393;
  assign c394 = (a393 & b393) | (a393 & c393) | (b393 & c393);
  wire c_sub394;
  assign c_sub394 = (a393 & b_inv393) | (a393 & c393) | (b_inv393 & c393);
  wire s394, sub394, and394, or394;
  wire b_inv394;
  assign b_inv394 = ~b394;
  assign s394  = a394 ^ b394 ^ c394;
  assign sub394 = a394 ^ b_inv394 ^ c394;
  assign and394 = a394 & b394;
  assign or394  = a394 | b394;
  assign c395 = (a394 & b394) | (a394 & c394) | (b394 & c394);
  wire c_sub395;
  assign c_sub395 = (a394 & b_inv394) | (a394 & c394) | (b_inv394 & c394);
  wire s395, sub395, and395, or395;
  wire b_inv395;
  assign b_inv395 = ~b395;
  assign s395  = a395 ^ b395 ^ c395;
  assign sub395 = a395 ^ b_inv395 ^ c395;
  assign and395 = a395 & b395;
  assign or395  = a395 | b395;
  assign c396 = (a395 & b395) | (a395 & c395) | (b395 & c395);
  wire c_sub396;
  assign c_sub396 = (a395 & b_inv395) | (a395 & c395) | (b_inv395 & c395);
  wire s396, sub396, and396, or396;
  wire b_inv396;
  assign b_inv396 = ~b396;
  assign s396  = a396 ^ b396 ^ c396;
  assign sub396 = a396 ^ b_inv396 ^ c396;
  assign and396 = a396 & b396;
  assign or396  = a396 | b396;
  assign c397 = (a396 & b396) | (a396 & c396) | (b396 & c396);
  wire c_sub397;
  assign c_sub397 = (a396 & b_inv396) | (a396 & c396) | (b_inv396 & c396);
  wire s397, sub397, and397, or397;
  wire b_inv397;
  assign b_inv397 = ~b397;
  assign s397  = a397 ^ b397 ^ c397;
  assign sub397 = a397 ^ b_inv397 ^ c397;
  assign and397 = a397 & b397;
  assign or397  = a397 | b397;
  assign c398 = (a397 & b397) | (a397 & c397) | (b397 & c397);
  wire c_sub398;
  assign c_sub398 = (a397 & b_inv397) | (a397 & c397) | (b_inv397 & c397);
  wire s398, sub398, and398, or398;
  wire b_inv398;
  assign b_inv398 = ~b398;
  assign s398  = a398 ^ b398 ^ c398;
  assign sub398 = a398 ^ b_inv398 ^ c398;
  assign and398 = a398 & b398;
  assign or398  = a398 | b398;
  assign c399 = (a398 & b398) | (a398 & c398) | (b398 & c398);
  wire c_sub399;
  assign c_sub399 = (a398 & b_inv398) | (a398 & c398) | (b_inv398 & c398);
  wire s399, sub399, and399, or399;
  wire b_inv399;
  assign b_inv399 = ~b399;
  assign s399  = a399 ^ b399 ^ c399;
  assign sub399 = a399 ^ b_inv399 ^ c399;
  assign and399 = a399 & b399;
  assign or399  = a399 | b399;
  assign c400 = (a399 & b399) | (a399 & c399) | (b399 & c399);
  wire c_sub400;
  assign c_sub400 = (a399 & b_inv399) | (a399 & c399) | (b_inv399 & c399);
  wire s400, sub400, and400, or400;
  wire b_inv400;
  assign b_inv400 = ~b400;
  assign s400  = a400 ^ b400 ^ c400;
  assign sub400 = a400 ^ b_inv400 ^ c400;
  assign and400 = a400 & b400;
  assign or400  = a400 | b400;
  assign c401 = (a400 & b400) | (a400 & c400) | (b400 & c400);
  wire c_sub401;
  assign c_sub401 = (a400 & b_inv400) | (a400 & c400) | (b_inv400 & c400);
  wire s401, sub401, and401, or401;
  wire b_inv401;
  assign b_inv401 = ~b401;
  assign s401  = a401 ^ b401 ^ c401;
  assign sub401 = a401 ^ b_inv401 ^ c401;
  assign and401 = a401 & b401;
  assign or401  = a401 | b401;
  assign c402 = (a401 & b401) | (a401 & c401) | (b401 & c401);
  wire c_sub402;
  assign c_sub402 = (a401 & b_inv401) | (a401 & c401) | (b_inv401 & c401);
  wire s402, sub402, and402, or402;
  wire b_inv402;
  assign b_inv402 = ~b402;
  assign s402  = a402 ^ b402 ^ c402;
  assign sub402 = a402 ^ b_inv402 ^ c402;
  assign and402 = a402 & b402;
  assign or402  = a402 | b402;
  assign c403 = (a402 & b402) | (a402 & c402) | (b402 & c402);
  wire c_sub403;
  assign c_sub403 = (a402 & b_inv402) | (a402 & c402) | (b_inv402 & c402);
  wire s403, sub403, and403, or403;
  wire b_inv403;
  assign b_inv403 = ~b403;
  assign s403  = a403 ^ b403 ^ c403;
  assign sub403 = a403 ^ b_inv403 ^ c403;
  assign and403 = a403 & b403;
  assign or403  = a403 | b403;
  assign c404 = (a403 & b403) | (a403 & c403) | (b403 & c403);
  wire c_sub404;
  assign c_sub404 = (a403 & b_inv403) | (a403 & c403) | (b_inv403 & c403);
  wire s404, sub404, and404, or404;
  wire b_inv404;
  assign b_inv404 = ~b404;
  assign s404  = a404 ^ b404 ^ c404;
  assign sub404 = a404 ^ b_inv404 ^ c404;
  assign and404 = a404 & b404;
  assign or404  = a404 | b404;
  assign c405 = (a404 & b404) | (a404 & c404) | (b404 & c404);
  wire c_sub405;
  assign c_sub405 = (a404 & b_inv404) | (a404 & c404) | (b_inv404 & c404);
  wire s405, sub405, and405, or405;
  wire b_inv405;
  assign b_inv405 = ~b405;
  assign s405  = a405 ^ b405 ^ c405;
  assign sub405 = a405 ^ b_inv405 ^ c405;
  assign and405 = a405 & b405;
  assign or405  = a405 | b405;
  assign c406 = (a405 & b405) | (a405 & c405) | (b405 & c405);
  wire c_sub406;
  assign c_sub406 = (a405 & b_inv405) | (a405 & c405) | (b_inv405 & c405);
  wire s406, sub406, and406, or406;
  wire b_inv406;
  assign b_inv406 = ~b406;
  assign s406  = a406 ^ b406 ^ c406;
  assign sub406 = a406 ^ b_inv406 ^ c406;
  assign and406 = a406 & b406;
  assign or406  = a406 | b406;
  assign c407 = (a406 & b406) | (a406 & c406) | (b406 & c406);
  wire c_sub407;
  assign c_sub407 = (a406 & b_inv406) | (a406 & c406) | (b_inv406 & c406);
  wire s407, sub407, and407, or407;
  wire b_inv407;
  assign b_inv407 = ~b407;
  assign s407  = a407 ^ b407 ^ c407;
  assign sub407 = a407 ^ b_inv407 ^ c407;
  assign and407 = a407 & b407;
  assign or407  = a407 | b407;
  assign c408 = (a407 & b407) | (a407 & c407) | (b407 & c407);
  wire c_sub408;
  assign c_sub408 = (a407 & b_inv407) | (a407 & c407) | (b_inv407 & c407);
  wire s408, sub408, and408, or408;
  wire b_inv408;
  assign b_inv408 = ~b408;
  assign s408  = a408 ^ b408 ^ c408;
  assign sub408 = a408 ^ b_inv408 ^ c408;
  assign and408 = a408 & b408;
  assign or408  = a408 | b408;
  assign c409 = (a408 & b408) | (a408 & c408) | (b408 & c408);
  wire c_sub409;
  assign c_sub409 = (a408 & b_inv408) | (a408 & c408) | (b_inv408 & c408);
  wire s409, sub409, and409, or409;
  wire b_inv409;
  assign b_inv409 = ~b409;
  assign s409  = a409 ^ b409 ^ c409;
  assign sub409 = a409 ^ b_inv409 ^ c409;
  assign and409 = a409 & b409;
  assign or409  = a409 | b409;
  assign c410 = (a409 & b409) | (a409 & c409) | (b409 & c409);
  wire c_sub410;
  assign c_sub410 = (a409 & b_inv409) | (a409 & c409) | (b_inv409 & c409);
  wire s410, sub410, and410, or410;
  wire b_inv410;
  assign b_inv410 = ~b410;
  assign s410  = a410 ^ b410 ^ c410;
  assign sub410 = a410 ^ b_inv410 ^ c410;
  assign and410 = a410 & b410;
  assign or410  = a410 | b410;
  assign c411 = (a410 & b410) | (a410 & c410) | (b410 & c410);
  wire c_sub411;
  assign c_sub411 = (a410 & b_inv410) | (a410 & c410) | (b_inv410 & c410);
  wire s411, sub411, and411, or411;
  wire b_inv411;
  assign b_inv411 = ~b411;
  assign s411  = a411 ^ b411 ^ c411;
  assign sub411 = a411 ^ b_inv411 ^ c411;
  assign and411 = a411 & b411;
  assign or411  = a411 | b411;
  assign c412 = (a411 & b411) | (a411 & c411) | (b411 & c411);
  wire c_sub412;
  assign c_sub412 = (a411 & b_inv411) | (a411 & c411) | (b_inv411 & c411);
  wire s412, sub412, and412, or412;
  wire b_inv412;
  assign b_inv412 = ~b412;
  assign s412  = a412 ^ b412 ^ c412;
  assign sub412 = a412 ^ b_inv412 ^ c412;
  assign and412 = a412 & b412;
  assign or412  = a412 | b412;
  assign c413 = (a412 & b412) | (a412 & c412) | (b412 & c412);
  wire c_sub413;
  assign c_sub413 = (a412 & b_inv412) | (a412 & c412) | (b_inv412 & c412);
  wire s413, sub413, and413, or413;
  wire b_inv413;
  assign b_inv413 = ~b413;
  assign s413  = a413 ^ b413 ^ c413;
  assign sub413 = a413 ^ b_inv413 ^ c413;
  assign and413 = a413 & b413;
  assign or413  = a413 | b413;
  assign c414 = (a413 & b413) | (a413 & c413) | (b413 & c413);
  wire c_sub414;
  assign c_sub414 = (a413 & b_inv413) | (a413 & c413) | (b_inv413 & c413);
  wire s414, sub414, and414, or414;
  wire b_inv414;
  assign b_inv414 = ~b414;
  assign s414  = a414 ^ b414 ^ c414;
  assign sub414 = a414 ^ b_inv414 ^ c414;
  assign and414 = a414 & b414;
  assign or414  = a414 | b414;
  assign c415 = (a414 & b414) | (a414 & c414) | (b414 & c414);
  wire c_sub415;
  assign c_sub415 = (a414 & b_inv414) | (a414 & c414) | (b_inv414 & c414);
  wire s415, sub415, and415, or415;
  wire b_inv415;
  assign b_inv415 = ~b415;
  assign s415  = a415 ^ b415 ^ c415;
  assign sub415 = a415 ^ b_inv415 ^ c415;
  assign and415 = a415 & b415;
  assign or415  = a415 | b415;
  assign c416 = (a415 & b415) | (a415 & c415) | (b415 & c415);
  wire c_sub416;
  assign c_sub416 = (a415 & b_inv415) | (a415 & c415) | (b_inv415 & c415);
  wire s416, sub416, and416, or416;
  wire b_inv416;
  assign b_inv416 = ~b416;
  assign s416  = a416 ^ b416 ^ c416;
  assign sub416 = a416 ^ b_inv416 ^ c416;
  assign and416 = a416 & b416;
  assign or416  = a416 | b416;
  assign c417 = (a416 & b416) | (a416 & c416) | (b416 & c416);
  wire c_sub417;
  assign c_sub417 = (a416 & b_inv416) | (a416 & c416) | (b_inv416 & c416);
  wire s417, sub417, and417, or417;
  wire b_inv417;
  assign b_inv417 = ~b417;
  assign s417  = a417 ^ b417 ^ c417;
  assign sub417 = a417 ^ b_inv417 ^ c417;
  assign and417 = a417 & b417;
  assign or417  = a417 | b417;
  assign c418 = (a417 & b417) | (a417 & c417) | (b417 & c417);
  wire c_sub418;
  assign c_sub418 = (a417 & b_inv417) | (a417 & c417) | (b_inv417 & c417);
  wire s418, sub418, and418, or418;
  wire b_inv418;
  assign b_inv418 = ~b418;
  assign s418  = a418 ^ b418 ^ c418;
  assign sub418 = a418 ^ b_inv418 ^ c418;
  assign and418 = a418 & b418;
  assign or418  = a418 | b418;
  assign c419 = (a418 & b418) | (a418 & c418) | (b418 & c418);
  wire c_sub419;
  assign c_sub419 = (a418 & b_inv418) | (a418 & c418) | (b_inv418 & c418);
  wire s419, sub419, and419, or419;
  wire b_inv419;
  assign b_inv419 = ~b419;
  assign s419  = a419 ^ b419 ^ c419;
  assign sub419 = a419 ^ b_inv419 ^ c419;
  assign and419 = a419 & b419;
  assign or419  = a419 | b419;
  assign c420 = (a419 & b419) | (a419 & c419) | (b419 & c419);
  wire c_sub420;
  assign c_sub420 = (a419 & b_inv419) | (a419 & c419) | (b_inv419 & c419);
  wire s420, sub420, and420, or420;
  wire b_inv420;
  assign b_inv420 = ~b420;
  assign s420  = a420 ^ b420 ^ c420;
  assign sub420 = a420 ^ b_inv420 ^ c420;
  assign and420 = a420 & b420;
  assign or420  = a420 | b420;
  assign c421 = (a420 & b420) | (a420 & c420) | (b420 & c420);
  wire c_sub421;
  assign c_sub421 = (a420 & b_inv420) | (a420 & c420) | (b_inv420 & c420);
  wire s421, sub421, and421, or421;
  wire b_inv421;
  assign b_inv421 = ~b421;
  assign s421  = a421 ^ b421 ^ c421;
  assign sub421 = a421 ^ b_inv421 ^ c421;
  assign and421 = a421 & b421;
  assign or421  = a421 | b421;
  assign c422 = (a421 & b421) | (a421 & c421) | (b421 & c421);
  wire c_sub422;
  assign c_sub422 = (a421 & b_inv421) | (a421 & c421) | (b_inv421 & c421);
  wire s422, sub422, and422, or422;
  wire b_inv422;
  assign b_inv422 = ~b422;
  assign s422  = a422 ^ b422 ^ c422;
  assign sub422 = a422 ^ b_inv422 ^ c422;
  assign and422 = a422 & b422;
  assign or422  = a422 | b422;
  assign c423 = (a422 & b422) | (a422 & c422) | (b422 & c422);
  wire c_sub423;
  assign c_sub423 = (a422 & b_inv422) | (a422 & c422) | (b_inv422 & c422);
  wire s423, sub423, and423, or423;
  wire b_inv423;
  assign b_inv423 = ~b423;
  assign s423  = a423 ^ b423 ^ c423;
  assign sub423 = a423 ^ b_inv423 ^ c423;
  assign and423 = a423 & b423;
  assign or423  = a423 | b423;
  assign c424 = (a423 & b423) | (a423 & c423) | (b423 & c423);
  wire c_sub424;
  assign c_sub424 = (a423 & b_inv423) | (a423 & c423) | (b_inv423 & c423);
  wire s424, sub424, and424, or424;
  wire b_inv424;
  assign b_inv424 = ~b424;
  assign s424  = a424 ^ b424 ^ c424;
  assign sub424 = a424 ^ b_inv424 ^ c424;
  assign and424 = a424 & b424;
  assign or424  = a424 | b424;
  assign c425 = (a424 & b424) | (a424 & c424) | (b424 & c424);
  wire c_sub425;
  assign c_sub425 = (a424 & b_inv424) | (a424 & c424) | (b_inv424 & c424);
  wire s425, sub425, and425, or425;
  wire b_inv425;
  assign b_inv425 = ~b425;
  assign s425  = a425 ^ b425 ^ c425;
  assign sub425 = a425 ^ b_inv425 ^ c425;
  assign and425 = a425 & b425;
  assign or425  = a425 | b425;
  assign c426 = (a425 & b425) | (a425 & c425) | (b425 & c425);
  wire c_sub426;
  assign c_sub426 = (a425 & b_inv425) | (a425 & c425) | (b_inv425 & c425);
  wire s426, sub426, and426, or426;
  wire b_inv426;
  assign b_inv426 = ~b426;
  assign s426  = a426 ^ b426 ^ c426;
  assign sub426 = a426 ^ b_inv426 ^ c426;
  assign and426 = a426 & b426;
  assign or426  = a426 | b426;
  assign c427 = (a426 & b426) | (a426 & c426) | (b426 & c426);
  wire c_sub427;
  assign c_sub427 = (a426 & b_inv426) | (a426 & c426) | (b_inv426 & c426);
  wire s427, sub427, and427, or427;
  wire b_inv427;
  assign b_inv427 = ~b427;
  assign s427  = a427 ^ b427 ^ c427;
  assign sub427 = a427 ^ b_inv427 ^ c427;
  assign and427 = a427 & b427;
  assign or427  = a427 | b427;
  assign c428 = (a427 & b427) | (a427 & c427) | (b427 & c427);
  wire c_sub428;
  assign c_sub428 = (a427 & b_inv427) | (a427 & c427) | (b_inv427 & c427);
  wire s428, sub428, and428, or428;
  wire b_inv428;
  assign b_inv428 = ~b428;
  assign s428  = a428 ^ b428 ^ c428;
  assign sub428 = a428 ^ b_inv428 ^ c428;
  assign and428 = a428 & b428;
  assign or428  = a428 | b428;
  assign c429 = (a428 & b428) | (a428 & c428) | (b428 & c428);
  wire c_sub429;
  assign c_sub429 = (a428 & b_inv428) | (a428 & c428) | (b_inv428 & c428);
  wire s429, sub429, and429, or429;
  wire b_inv429;
  assign b_inv429 = ~b429;
  assign s429  = a429 ^ b429 ^ c429;
  assign sub429 = a429 ^ b_inv429 ^ c429;
  assign and429 = a429 & b429;
  assign or429  = a429 | b429;
  assign c430 = (a429 & b429) | (a429 & c429) | (b429 & c429);
  wire c_sub430;
  assign c_sub430 = (a429 & b_inv429) | (a429 & c429) | (b_inv429 & c429);
  wire s430, sub430, and430, or430;
  wire b_inv430;
  assign b_inv430 = ~b430;
  assign s430  = a430 ^ b430 ^ c430;
  assign sub430 = a430 ^ b_inv430 ^ c430;
  assign and430 = a430 & b430;
  assign or430  = a430 | b430;
  assign c431 = (a430 & b430) | (a430 & c430) | (b430 & c430);
  wire c_sub431;
  assign c_sub431 = (a430 & b_inv430) | (a430 & c430) | (b_inv430 & c430);
  wire s431, sub431, and431, or431;
  wire b_inv431;
  assign b_inv431 = ~b431;
  assign s431  = a431 ^ b431 ^ c431;
  assign sub431 = a431 ^ b_inv431 ^ c431;
  assign and431 = a431 & b431;
  assign or431  = a431 | b431;
  assign c432 = (a431 & b431) | (a431 & c431) | (b431 & c431);
  wire c_sub432;
  assign c_sub432 = (a431 & b_inv431) | (a431 & c431) | (b_inv431 & c431);
  wire s432, sub432, and432, or432;
  wire b_inv432;
  assign b_inv432 = ~b432;
  assign s432  = a432 ^ b432 ^ c432;
  assign sub432 = a432 ^ b_inv432 ^ c432;
  assign and432 = a432 & b432;
  assign or432  = a432 | b432;
  assign c433 = (a432 & b432) | (a432 & c432) | (b432 & c432);
  wire c_sub433;
  assign c_sub433 = (a432 & b_inv432) | (a432 & c432) | (b_inv432 & c432);
  wire s433, sub433, and433, or433;
  wire b_inv433;
  assign b_inv433 = ~b433;
  assign s433  = a433 ^ b433 ^ c433;
  assign sub433 = a433 ^ b_inv433 ^ c433;
  assign and433 = a433 & b433;
  assign or433  = a433 | b433;
  assign c434 = (a433 & b433) | (a433 & c433) | (b433 & c433);
  wire c_sub434;
  assign c_sub434 = (a433 & b_inv433) | (a433 & c433) | (b_inv433 & c433);
  wire s434, sub434, and434, or434;
  wire b_inv434;
  assign b_inv434 = ~b434;
  assign s434  = a434 ^ b434 ^ c434;
  assign sub434 = a434 ^ b_inv434 ^ c434;
  assign and434 = a434 & b434;
  assign or434  = a434 | b434;
  assign c435 = (a434 & b434) | (a434 & c434) | (b434 & c434);
  wire c_sub435;
  assign c_sub435 = (a434 & b_inv434) | (a434 & c434) | (b_inv434 & c434);
  wire s435, sub435, and435, or435;
  wire b_inv435;
  assign b_inv435 = ~b435;
  assign s435  = a435 ^ b435 ^ c435;
  assign sub435 = a435 ^ b_inv435 ^ c435;
  assign and435 = a435 & b435;
  assign or435  = a435 | b435;
  assign c436 = (a435 & b435) | (a435 & c435) | (b435 & c435);
  wire c_sub436;
  assign c_sub436 = (a435 & b_inv435) | (a435 & c435) | (b_inv435 & c435);
  wire s436, sub436, and436, or436;
  wire b_inv436;
  assign b_inv436 = ~b436;
  assign s436  = a436 ^ b436 ^ c436;
  assign sub436 = a436 ^ b_inv436 ^ c436;
  assign and436 = a436 & b436;
  assign or436  = a436 | b436;
  assign c437 = (a436 & b436) | (a436 & c436) | (b436 & c436);
  wire c_sub437;
  assign c_sub437 = (a436 & b_inv436) | (a436 & c436) | (b_inv436 & c436);
  wire s437, sub437, and437, or437;
  wire b_inv437;
  assign b_inv437 = ~b437;
  assign s437  = a437 ^ b437 ^ c437;
  assign sub437 = a437 ^ b_inv437 ^ c437;
  assign and437 = a437 & b437;
  assign or437  = a437 | b437;
  assign c438 = (a437 & b437) | (a437 & c437) | (b437 & c437);
  wire c_sub438;
  assign c_sub438 = (a437 & b_inv437) | (a437 & c437) | (b_inv437 & c437);
  wire s438, sub438, and438, or438;
  wire b_inv438;
  assign b_inv438 = ~b438;
  assign s438  = a438 ^ b438 ^ c438;
  assign sub438 = a438 ^ b_inv438 ^ c438;
  assign and438 = a438 & b438;
  assign or438  = a438 | b438;
  assign c439 = (a438 & b438) | (a438 & c438) | (b438 & c438);
  wire c_sub439;
  assign c_sub439 = (a438 & b_inv438) | (a438 & c438) | (b_inv438 & c438);
  wire s439, sub439, and439, or439;
  wire b_inv439;
  assign b_inv439 = ~b439;
  assign s439  = a439 ^ b439 ^ c439;
  assign sub439 = a439 ^ b_inv439 ^ c439;
  assign and439 = a439 & b439;
  assign or439  = a439 | b439;
  assign c440 = (a439 & b439) | (a439 & c439) | (b439 & c439);
  wire c_sub440;
  assign c_sub440 = (a439 & b_inv439) | (a439 & c439) | (b_inv439 & c439);
  wire s440, sub440, and440, or440;
  wire b_inv440;
  assign b_inv440 = ~b440;
  assign s440  = a440 ^ b440 ^ c440;
  assign sub440 = a440 ^ b_inv440 ^ c440;
  assign and440 = a440 & b440;
  assign or440  = a440 | b440;
  assign c441 = (a440 & b440) | (a440 & c440) | (b440 & c440);
  wire c_sub441;
  assign c_sub441 = (a440 & b_inv440) | (a440 & c440) | (b_inv440 & c440);
  wire s441, sub441, and441, or441;
  wire b_inv441;
  assign b_inv441 = ~b441;
  assign s441  = a441 ^ b441 ^ c441;
  assign sub441 = a441 ^ b_inv441 ^ c441;
  assign and441 = a441 & b441;
  assign or441  = a441 | b441;
  assign c442 = (a441 & b441) | (a441 & c441) | (b441 & c441);
  wire c_sub442;
  assign c_sub442 = (a441 & b_inv441) | (a441 & c441) | (b_inv441 & c441);
  wire s442, sub442, and442, or442;
  wire b_inv442;
  assign b_inv442 = ~b442;
  assign s442  = a442 ^ b442 ^ c442;
  assign sub442 = a442 ^ b_inv442 ^ c442;
  assign and442 = a442 & b442;
  assign or442  = a442 | b442;
  assign c443 = (a442 & b442) | (a442 & c442) | (b442 & c442);
  wire c_sub443;
  assign c_sub443 = (a442 & b_inv442) | (a442 & c442) | (b_inv442 & c442);
  wire s443, sub443, and443, or443;
  wire b_inv443;
  assign b_inv443 = ~b443;
  assign s443  = a443 ^ b443 ^ c443;
  assign sub443 = a443 ^ b_inv443 ^ c443;
  assign and443 = a443 & b443;
  assign or443  = a443 | b443;
  assign c444 = (a443 & b443) | (a443 & c443) | (b443 & c443);
  wire c_sub444;
  assign c_sub444 = (a443 & b_inv443) | (a443 & c443) | (b_inv443 & c443);
  wire s444, sub444, and444, or444;
  wire b_inv444;
  assign b_inv444 = ~b444;
  assign s444  = a444 ^ b444 ^ c444;
  assign sub444 = a444 ^ b_inv444 ^ c444;
  assign and444 = a444 & b444;
  assign or444  = a444 | b444;
  assign c445 = (a444 & b444) | (a444 & c444) | (b444 & c444);
  wire c_sub445;
  assign c_sub445 = (a444 & b_inv444) | (a444 & c444) | (b_inv444 & c444);
  wire s445, sub445, and445, or445;
  wire b_inv445;
  assign b_inv445 = ~b445;
  assign s445  = a445 ^ b445 ^ c445;
  assign sub445 = a445 ^ b_inv445 ^ c445;
  assign and445 = a445 & b445;
  assign or445  = a445 | b445;
  assign c446 = (a445 & b445) | (a445 & c445) | (b445 & c445);
  wire c_sub446;
  assign c_sub446 = (a445 & b_inv445) | (a445 & c445) | (b_inv445 & c445);
  wire s446, sub446, and446, or446;
  wire b_inv446;
  assign b_inv446 = ~b446;
  assign s446  = a446 ^ b446 ^ c446;
  assign sub446 = a446 ^ b_inv446 ^ c446;
  assign and446 = a446 & b446;
  assign or446  = a446 | b446;
  assign c447 = (a446 & b446) | (a446 & c446) | (b446 & c446);
  wire c_sub447;
  assign c_sub447 = (a446 & b_inv446) | (a446 & c446) | (b_inv446 & c446);
  wire s447, sub447, and447, or447;
  wire b_inv447;
  assign b_inv447 = ~b447;
  assign s447  = a447 ^ b447 ^ c447;
  assign sub447 = a447 ^ b_inv447 ^ c447;
  assign and447 = a447 & b447;
  assign or447  = a447 | b447;
  assign c448 = (a447 & b447) | (a447 & c447) | (b447 & c447);
  wire c_sub448;
  assign c_sub448 = (a447 & b_inv447) | (a447 & c447) | (b_inv447 & c447);
  wire s448, sub448, and448, or448;
  wire b_inv448;
  assign b_inv448 = ~b448;
  assign s448  = a448 ^ b448 ^ c448;
  assign sub448 = a448 ^ b_inv448 ^ c448;
  assign and448 = a448 & b448;
  assign or448  = a448 | b448;
  assign c449 = (a448 & b448) | (a448 & c448) | (b448 & c448);
  wire c_sub449;
  assign c_sub449 = (a448 & b_inv448) | (a448 & c448) | (b_inv448 & c448);
  wire s449, sub449, and449, or449;
  wire b_inv449;
  assign b_inv449 = ~b449;
  assign s449  = a449 ^ b449 ^ c449;
  assign sub449 = a449 ^ b_inv449 ^ c449;
  assign and449 = a449 & b449;
  assign or449  = a449 | b449;
  assign c450 = (a449 & b449) | (a449 & c449) | (b449 & c449);
  wire c_sub450;
  assign c_sub450 = (a449 & b_inv449) | (a449 & c449) | (b_inv449 & c449);
  wire s450, sub450, and450, or450;
  wire b_inv450;
  assign b_inv450 = ~b450;
  assign s450  = a450 ^ b450 ^ c450;
  assign sub450 = a450 ^ b_inv450 ^ c450;
  assign and450 = a450 & b450;
  assign or450  = a450 | b450;
  assign c451 = (a450 & b450) | (a450 & c450) | (b450 & c450);
  wire c_sub451;
  assign c_sub451 = (a450 & b_inv450) | (a450 & c450) | (b_inv450 & c450);
  wire s451, sub451, and451, or451;
  wire b_inv451;
  assign b_inv451 = ~b451;
  assign s451  = a451 ^ b451 ^ c451;
  assign sub451 = a451 ^ b_inv451 ^ c451;
  assign and451 = a451 & b451;
  assign or451  = a451 | b451;
  assign c452 = (a451 & b451) | (a451 & c451) | (b451 & c451);
  wire c_sub452;
  assign c_sub452 = (a451 & b_inv451) | (a451 & c451) | (b_inv451 & c451);
  wire s452, sub452, and452, or452;
  wire b_inv452;
  assign b_inv452 = ~b452;
  assign s452  = a452 ^ b452 ^ c452;
  assign sub452 = a452 ^ b_inv452 ^ c452;
  assign and452 = a452 & b452;
  assign or452  = a452 | b452;
  assign c453 = (a452 & b452) | (a452 & c452) | (b452 & c452);
  wire c_sub453;
  assign c_sub453 = (a452 & b_inv452) | (a452 & c452) | (b_inv452 & c452);
  wire s453, sub453, and453, or453;
  wire b_inv453;
  assign b_inv453 = ~b453;
  assign s453  = a453 ^ b453 ^ c453;
  assign sub453 = a453 ^ b_inv453 ^ c453;
  assign and453 = a453 & b453;
  assign or453  = a453 | b453;
  assign c454 = (a453 & b453) | (a453 & c453) | (b453 & c453);
  wire c_sub454;
  assign c_sub454 = (a453 & b_inv453) | (a453 & c453) | (b_inv453 & c453);
  wire s454, sub454, and454, or454;
  wire b_inv454;
  assign b_inv454 = ~b454;
  assign s454  = a454 ^ b454 ^ c454;
  assign sub454 = a454 ^ b_inv454 ^ c454;
  assign and454 = a454 & b454;
  assign or454  = a454 | b454;
  assign c455 = (a454 & b454) | (a454 & c454) | (b454 & c454);
  wire c_sub455;
  assign c_sub455 = (a454 & b_inv454) | (a454 & c454) | (b_inv454 & c454);
  wire s455, sub455, and455, or455;
  wire b_inv455;
  assign b_inv455 = ~b455;
  assign s455  = a455 ^ b455 ^ c455;
  assign sub455 = a455 ^ b_inv455 ^ c455;
  assign and455 = a455 & b455;
  assign or455  = a455 | b455;
  assign c456 = (a455 & b455) | (a455 & c455) | (b455 & c455);
  wire c_sub456;
  assign c_sub456 = (a455 & b_inv455) | (a455 & c455) | (b_inv455 & c455);
  wire s456, sub456, and456, or456;
  wire b_inv456;
  assign b_inv456 = ~b456;
  assign s456  = a456 ^ b456 ^ c456;
  assign sub456 = a456 ^ b_inv456 ^ c456;
  assign and456 = a456 & b456;
  assign or456  = a456 | b456;
  assign c457 = (a456 & b456) | (a456 & c456) | (b456 & c456);
  wire c_sub457;
  assign c_sub457 = (a456 & b_inv456) | (a456 & c456) | (b_inv456 & c456);
  wire s457, sub457, and457, or457;
  wire b_inv457;
  assign b_inv457 = ~b457;
  assign s457  = a457 ^ b457 ^ c457;
  assign sub457 = a457 ^ b_inv457 ^ c457;
  assign and457 = a457 & b457;
  assign or457  = a457 | b457;
  assign c458 = (a457 & b457) | (a457 & c457) | (b457 & c457);
  wire c_sub458;
  assign c_sub458 = (a457 & b_inv457) | (a457 & c457) | (b_inv457 & c457);
  wire s458, sub458, and458, or458;
  wire b_inv458;
  assign b_inv458 = ~b458;
  assign s458  = a458 ^ b458 ^ c458;
  assign sub458 = a458 ^ b_inv458 ^ c458;
  assign and458 = a458 & b458;
  assign or458  = a458 | b458;
  assign c459 = (a458 & b458) | (a458 & c458) | (b458 & c458);
  wire c_sub459;
  assign c_sub459 = (a458 & b_inv458) | (a458 & c458) | (b_inv458 & c458);
  wire s459, sub459, and459, or459;
  wire b_inv459;
  assign b_inv459 = ~b459;
  assign s459  = a459 ^ b459 ^ c459;
  assign sub459 = a459 ^ b_inv459 ^ c459;
  assign and459 = a459 & b459;
  assign or459  = a459 | b459;
  assign c460 = (a459 & b459) | (a459 & c459) | (b459 & c459);
  wire c_sub460;
  assign c_sub460 = (a459 & b_inv459) | (a459 & c459) | (b_inv459 & c459);
  wire s460, sub460, and460, or460;
  wire b_inv460;
  assign b_inv460 = ~b460;
  assign s460  = a460 ^ b460 ^ c460;
  assign sub460 = a460 ^ b_inv460 ^ c460;
  assign and460 = a460 & b460;
  assign or460  = a460 | b460;
  assign c461 = (a460 & b460) | (a460 & c460) | (b460 & c460);
  wire c_sub461;
  assign c_sub461 = (a460 & b_inv460) | (a460 & c460) | (b_inv460 & c460);
  wire s461, sub461, and461, or461;
  wire b_inv461;
  assign b_inv461 = ~b461;
  assign s461  = a461 ^ b461 ^ c461;
  assign sub461 = a461 ^ b_inv461 ^ c461;
  assign and461 = a461 & b461;
  assign or461  = a461 | b461;
  assign c462 = (a461 & b461) | (a461 & c461) | (b461 & c461);
  wire c_sub462;
  assign c_sub462 = (a461 & b_inv461) | (a461 & c461) | (b_inv461 & c461);
  wire s462, sub462, and462, or462;
  wire b_inv462;
  assign b_inv462 = ~b462;
  assign s462  = a462 ^ b462 ^ c462;
  assign sub462 = a462 ^ b_inv462 ^ c462;
  assign and462 = a462 & b462;
  assign or462  = a462 | b462;
  assign c463 = (a462 & b462) | (a462 & c462) | (b462 & c462);
  wire c_sub463;
  assign c_sub463 = (a462 & b_inv462) | (a462 & c462) | (b_inv462 & c462);
  wire s463, sub463, and463, or463;
  wire b_inv463;
  assign b_inv463 = ~b463;
  assign s463  = a463 ^ b463 ^ c463;
  assign sub463 = a463 ^ b_inv463 ^ c463;
  assign and463 = a463 & b463;
  assign or463  = a463 | b463;
  assign c464 = (a463 & b463) | (a463 & c463) | (b463 & c463);
  wire c_sub464;
  assign c_sub464 = (a463 & b_inv463) | (a463 & c463) | (b_inv463 & c463);
  wire s464, sub464, and464, or464;
  wire b_inv464;
  assign b_inv464 = ~b464;
  assign s464  = a464 ^ b464 ^ c464;
  assign sub464 = a464 ^ b_inv464 ^ c464;
  assign and464 = a464 & b464;
  assign or464  = a464 | b464;
  assign c465 = (a464 & b464) | (a464 & c464) | (b464 & c464);
  wire c_sub465;
  assign c_sub465 = (a464 & b_inv464) | (a464 & c464) | (b_inv464 & c464);
  wire s465, sub465, and465, or465;
  wire b_inv465;
  assign b_inv465 = ~b465;
  assign s465  = a465 ^ b465 ^ c465;
  assign sub465 = a465 ^ b_inv465 ^ c465;
  assign and465 = a465 & b465;
  assign or465  = a465 | b465;
  assign c466 = (a465 & b465) | (a465 & c465) | (b465 & c465);
  wire c_sub466;
  assign c_sub466 = (a465 & b_inv465) | (a465 & c465) | (b_inv465 & c465);
  wire s466, sub466, and466, or466;
  wire b_inv466;
  assign b_inv466 = ~b466;
  assign s466  = a466 ^ b466 ^ c466;
  assign sub466 = a466 ^ b_inv466 ^ c466;
  assign and466 = a466 & b466;
  assign or466  = a466 | b466;
  assign c467 = (a466 & b466) | (a466 & c466) | (b466 & c466);
  wire c_sub467;
  assign c_sub467 = (a466 & b_inv466) | (a466 & c466) | (b_inv466 & c466);
  wire s467, sub467, and467, or467;
  wire b_inv467;
  assign b_inv467 = ~b467;
  assign s467  = a467 ^ b467 ^ c467;
  assign sub467 = a467 ^ b_inv467 ^ c467;
  assign and467 = a467 & b467;
  assign or467  = a467 | b467;
  assign c468 = (a467 & b467) | (a467 & c467) | (b467 & c467);
  wire c_sub468;
  assign c_sub468 = (a467 & b_inv467) | (a467 & c467) | (b_inv467 & c467);
  wire s468, sub468, and468, or468;
  wire b_inv468;
  assign b_inv468 = ~b468;
  assign s468  = a468 ^ b468 ^ c468;
  assign sub468 = a468 ^ b_inv468 ^ c468;
  assign and468 = a468 & b468;
  assign or468  = a468 | b468;
  assign c469 = (a468 & b468) | (a468 & c468) | (b468 & c468);
  wire c_sub469;
  assign c_sub469 = (a468 & b_inv468) | (a468 & c468) | (b_inv468 & c468);
  wire s469, sub469, and469, or469;
  wire b_inv469;
  assign b_inv469 = ~b469;
  assign s469  = a469 ^ b469 ^ c469;
  assign sub469 = a469 ^ b_inv469 ^ c469;
  assign and469 = a469 & b469;
  assign or469  = a469 | b469;
  assign c470 = (a469 & b469) | (a469 & c469) | (b469 & c469);
  wire c_sub470;
  assign c_sub470 = (a469 & b_inv469) | (a469 & c469) | (b_inv469 & c469);
  wire s470, sub470, and470, or470;
  wire b_inv470;
  assign b_inv470 = ~b470;
  assign s470  = a470 ^ b470 ^ c470;
  assign sub470 = a470 ^ b_inv470 ^ c470;
  assign and470 = a470 & b470;
  assign or470  = a470 | b470;
  assign c471 = (a470 & b470) | (a470 & c470) | (b470 & c470);
  wire c_sub471;
  assign c_sub471 = (a470 & b_inv470) | (a470 & c470) | (b_inv470 & c470);
  wire s471, sub471, and471, or471;
  wire b_inv471;
  assign b_inv471 = ~b471;
  assign s471  = a471 ^ b471 ^ c471;
  assign sub471 = a471 ^ b_inv471 ^ c471;
  assign and471 = a471 & b471;
  assign or471  = a471 | b471;
  assign c472 = (a471 & b471) | (a471 & c471) | (b471 & c471);
  wire c_sub472;
  assign c_sub472 = (a471 & b_inv471) | (a471 & c471) | (b_inv471 & c471);
  wire s472, sub472, and472, or472;
  wire b_inv472;
  assign b_inv472 = ~b472;
  assign s472  = a472 ^ b472 ^ c472;
  assign sub472 = a472 ^ b_inv472 ^ c472;
  assign and472 = a472 & b472;
  assign or472  = a472 | b472;
  assign c473 = (a472 & b472) | (a472 & c472) | (b472 & c472);
  wire c_sub473;
  assign c_sub473 = (a472 & b_inv472) | (a472 & c472) | (b_inv472 & c472);
  wire s473, sub473, and473, or473;
  wire b_inv473;
  assign b_inv473 = ~b473;
  assign s473  = a473 ^ b473 ^ c473;
  assign sub473 = a473 ^ b_inv473 ^ c473;
  assign and473 = a473 & b473;
  assign or473  = a473 | b473;
  assign c474 = (a473 & b473) | (a473 & c473) | (b473 & c473);
  wire c_sub474;
  assign c_sub474 = (a473 & b_inv473) | (a473 & c473) | (b_inv473 & c473);
  wire s474, sub474, and474, or474;
  wire b_inv474;
  assign b_inv474 = ~b474;
  assign s474  = a474 ^ b474 ^ c474;
  assign sub474 = a474 ^ b_inv474 ^ c474;
  assign and474 = a474 & b474;
  assign or474  = a474 | b474;
  assign c475 = (a474 & b474) | (a474 & c474) | (b474 & c474);
  wire c_sub475;
  assign c_sub475 = (a474 & b_inv474) | (a474 & c474) | (b_inv474 & c474);
  wire s475, sub475, and475, or475;
  wire b_inv475;
  assign b_inv475 = ~b475;
  assign s475  = a475 ^ b475 ^ c475;
  assign sub475 = a475 ^ b_inv475 ^ c475;
  assign and475 = a475 & b475;
  assign or475  = a475 | b475;
  assign c476 = (a475 & b475) | (a475 & c475) | (b475 & c475);
  wire c_sub476;
  assign c_sub476 = (a475 & b_inv475) | (a475 & c475) | (b_inv475 & c475);
  wire s476, sub476, and476, or476;
  wire b_inv476;
  assign b_inv476 = ~b476;
  assign s476  = a476 ^ b476 ^ c476;
  assign sub476 = a476 ^ b_inv476 ^ c476;
  assign and476 = a476 & b476;
  assign or476  = a476 | b476;
  assign c477 = (a476 & b476) | (a476 & c476) | (b476 & c476);
  wire c_sub477;
  assign c_sub477 = (a476 & b_inv476) | (a476 & c476) | (b_inv476 & c476);
  wire s477, sub477, and477, or477;
  wire b_inv477;
  assign b_inv477 = ~b477;
  assign s477  = a477 ^ b477 ^ c477;
  assign sub477 = a477 ^ b_inv477 ^ c477;
  assign and477 = a477 & b477;
  assign or477  = a477 | b477;
  assign c478 = (a477 & b477) | (a477 & c477) | (b477 & c477);
  wire c_sub478;
  assign c_sub478 = (a477 & b_inv477) | (a477 & c477) | (b_inv477 & c477);
  wire s478, sub478, and478, or478;
  wire b_inv478;
  assign b_inv478 = ~b478;
  assign s478  = a478 ^ b478 ^ c478;
  assign sub478 = a478 ^ b_inv478 ^ c478;
  assign and478 = a478 & b478;
  assign or478  = a478 | b478;
  assign c479 = (a478 & b478) | (a478 & c478) | (b478 & c478);
  wire c_sub479;
  assign c_sub479 = (a478 & b_inv478) | (a478 & c478) | (b_inv478 & c478);
  wire s479, sub479, and479, or479;
  wire b_inv479;
  assign b_inv479 = ~b479;
  assign s479  = a479 ^ b479 ^ c479;
  assign sub479 = a479 ^ b_inv479 ^ c479;
  assign and479 = a479 & b479;
  assign or479  = a479 | b479;
  assign c480 = (a479 & b479) | (a479 & c479) | (b479 & c479);
  wire c_sub480;
  assign c_sub480 = (a479 & b_inv479) | (a479 & c479) | (b_inv479 & c479);
  wire s480, sub480, and480, or480;
  wire b_inv480;
  assign b_inv480 = ~b480;
  assign s480  = a480 ^ b480 ^ c480;
  assign sub480 = a480 ^ b_inv480 ^ c480;
  assign and480 = a480 & b480;
  assign or480  = a480 | b480;
  assign c481 = (a480 & b480) | (a480 & c480) | (b480 & c480);
  wire c_sub481;
  assign c_sub481 = (a480 & b_inv480) | (a480 & c480) | (b_inv480 & c480);
  wire s481, sub481, and481, or481;
  wire b_inv481;
  assign b_inv481 = ~b481;
  assign s481  = a481 ^ b481 ^ c481;
  assign sub481 = a481 ^ b_inv481 ^ c481;
  assign and481 = a481 & b481;
  assign or481  = a481 | b481;
  assign c482 = (a481 & b481) | (a481 & c481) | (b481 & c481);
  wire c_sub482;
  assign c_sub482 = (a481 & b_inv481) | (a481 & c481) | (b_inv481 & c481);
  wire s482, sub482, and482, or482;
  wire b_inv482;
  assign b_inv482 = ~b482;
  assign s482  = a482 ^ b482 ^ c482;
  assign sub482 = a482 ^ b_inv482 ^ c482;
  assign and482 = a482 & b482;
  assign or482  = a482 | b482;
  assign c483 = (a482 & b482) | (a482 & c482) | (b482 & c482);
  wire c_sub483;
  assign c_sub483 = (a482 & b_inv482) | (a482 & c482) | (b_inv482 & c482);
  wire s483, sub483, and483, or483;
  wire b_inv483;
  assign b_inv483 = ~b483;
  assign s483  = a483 ^ b483 ^ c483;
  assign sub483 = a483 ^ b_inv483 ^ c483;
  assign and483 = a483 & b483;
  assign or483  = a483 | b483;
  assign c484 = (a483 & b483) | (a483 & c483) | (b483 & c483);
  wire c_sub484;
  assign c_sub484 = (a483 & b_inv483) | (a483 & c483) | (b_inv483 & c483);
  wire s484, sub484, and484, or484;
  wire b_inv484;
  assign b_inv484 = ~b484;
  assign s484  = a484 ^ b484 ^ c484;
  assign sub484 = a484 ^ b_inv484 ^ c484;
  assign and484 = a484 & b484;
  assign or484  = a484 | b484;
  assign c485 = (a484 & b484) | (a484 & c484) | (b484 & c484);
  wire c_sub485;
  assign c_sub485 = (a484 & b_inv484) | (a484 & c484) | (b_inv484 & c484);
  wire s485, sub485, and485, or485;
  wire b_inv485;
  assign b_inv485 = ~b485;
  assign s485  = a485 ^ b485 ^ c485;
  assign sub485 = a485 ^ b_inv485 ^ c485;
  assign and485 = a485 & b485;
  assign or485  = a485 | b485;
  assign c486 = (a485 & b485) | (a485 & c485) | (b485 & c485);
  wire c_sub486;
  assign c_sub486 = (a485 & b_inv485) | (a485 & c485) | (b_inv485 & c485);
  wire s486, sub486, and486, or486;
  wire b_inv486;
  assign b_inv486 = ~b486;
  assign s486  = a486 ^ b486 ^ c486;
  assign sub486 = a486 ^ b_inv486 ^ c486;
  assign and486 = a486 & b486;
  assign or486  = a486 | b486;
  assign c487 = (a486 & b486) | (a486 & c486) | (b486 & c486);
  wire c_sub487;
  assign c_sub487 = (a486 & b_inv486) | (a486 & c486) | (b_inv486 & c486);
  wire s487, sub487, and487, or487;
  wire b_inv487;
  assign b_inv487 = ~b487;
  assign s487  = a487 ^ b487 ^ c487;
  assign sub487 = a487 ^ b_inv487 ^ c487;
  assign and487 = a487 & b487;
  assign or487  = a487 | b487;
  assign c488 = (a487 & b487) | (a487 & c487) | (b487 & c487);
  wire c_sub488;
  assign c_sub488 = (a487 & b_inv487) | (a487 & c487) | (b_inv487 & c487);
  wire s488, sub488, and488, or488;
  wire b_inv488;
  assign b_inv488 = ~b488;
  assign s488  = a488 ^ b488 ^ c488;
  assign sub488 = a488 ^ b_inv488 ^ c488;
  assign and488 = a488 & b488;
  assign or488  = a488 | b488;
  assign c489 = (a488 & b488) | (a488 & c488) | (b488 & c488);
  wire c_sub489;
  assign c_sub489 = (a488 & b_inv488) | (a488 & c488) | (b_inv488 & c488);
  wire s489, sub489, and489, or489;
  wire b_inv489;
  assign b_inv489 = ~b489;
  assign s489  = a489 ^ b489 ^ c489;
  assign sub489 = a489 ^ b_inv489 ^ c489;
  assign and489 = a489 & b489;
  assign or489  = a489 | b489;
  assign c490 = (a489 & b489) | (a489 & c489) | (b489 & c489);
  wire c_sub490;
  assign c_sub490 = (a489 & b_inv489) | (a489 & c489) | (b_inv489 & c489);
  wire s490, sub490, and490, or490;
  wire b_inv490;
  assign b_inv490 = ~b490;
  assign s490  = a490 ^ b490 ^ c490;
  assign sub490 = a490 ^ b_inv490 ^ c490;
  assign and490 = a490 & b490;
  assign or490  = a490 | b490;
  assign c491 = (a490 & b490) | (a490 & c490) | (b490 & c490);
  wire c_sub491;
  assign c_sub491 = (a490 & b_inv490) | (a490 & c490) | (b_inv490 & c490);
  wire s491, sub491, and491, or491;
  wire b_inv491;
  assign b_inv491 = ~b491;
  assign s491  = a491 ^ b491 ^ c491;
  assign sub491 = a491 ^ b_inv491 ^ c491;
  assign and491 = a491 & b491;
  assign or491  = a491 | b491;
  assign c492 = (a491 & b491) | (a491 & c491) | (b491 & c491);
  wire c_sub492;
  assign c_sub492 = (a491 & b_inv491) | (a491 & c491) | (b_inv491 & c491);
  wire s492, sub492, and492, or492;
  wire b_inv492;
  assign b_inv492 = ~b492;
  assign s492  = a492 ^ b492 ^ c492;
  assign sub492 = a492 ^ b_inv492 ^ c492;
  assign and492 = a492 & b492;
  assign or492  = a492 | b492;
  assign c493 = (a492 & b492) | (a492 & c492) | (b492 & c492);
  wire c_sub493;
  assign c_sub493 = (a492 & b_inv492) | (a492 & c492) | (b_inv492 & c492);
  wire s493, sub493, and493, or493;
  wire b_inv493;
  assign b_inv493 = ~b493;
  assign s493  = a493 ^ b493 ^ c493;
  assign sub493 = a493 ^ b_inv493 ^ c493;
  assign and493 = a493 & b493;
  assign or493  = a493 | b493;
  assign c494 = (a493 & b493) | (a493 & c493) | (b493 & c493);
  wire c_sub494;
  assign c_sub494 = (a493 & b_inv493) | (a493 & c493) | (b_inv493 & c493);
  wire s494, sub494, and494, or494;
  wire b_inv494;
  assign b_inv494 = ~b494;
  assign s494  = a494 ^ b494 ^ c494;
  assign sub494 = a494 ^ b_inv494 ^ c494;
  assign and494 = a494 & b494;
  assign or494  = a494 | b494;
  assign c495 = (a494 & b494) | (a494 & c494) | (b494 & c494);
  wire c_sub495;
  assign c_sub495 = (a494 & b_inv494) | (a494 & c494) | (b_inv494 & c494);
  wire s495, sub495, and495, or495;
  wire b_inv495;
  assign b_inv495 = ~b495;
  assign s495  = a495 ^ b495 ^ c495;
  assign sub495 = a495 ^ b_inv495 ^ c495;
  assign and495 = a495 & b495;
  assign or495  = a495 | b495;
  assign c496 = (a495 & b495) | (a495 & c495) | (b495 & c495);
  wire c_sub496;
  assign c_sub496 = (a495 & b_inv495) | (a495 & c495) | (b_inv495 & c495);
  wire s496, sub496, and496, or496;
  wire b_inv496;
  assign b_inv496 = ~b496;
  assign s496  = a496 ^ b496 ^ c496;
  assign sub496 = a496 ^ b_inv496 ^ c496;
  assign and496 = a496 & b496;
  assign or496  = a496 | b496;
  assign c497 = (a496 & b496) | (a496 & c496) | (b496 & c496);
  wire c_sub497;
  assign c_sub497 = (a496 & b_inv496) | (a496 & c496) | (b_inv496 & c496);
  wire s497, sub497, and497, or497;
  wire b_inv497;
  assign b_inv497 = ~b497;
  assign s497  = a497 ^ b497 ^ c497;
  assign sub497 = a497 ^ b_inv497 ^ c497;
  assign and497 = a497 & b497;
  assign or497  = a497 | b497;
  assign c498 = (a497 & b497) | (a497 & c497) | (b497 & c497);
  wire c_sub498;
  assign c_sub498 = (a497 & b_inv497) | (a497 & c497) | (b_inv497 & c497);
  wire s498, sub498, and498, or498;
  wire b_inv498;
  assign b_inv498 = ~b498;
  assign s498  = a498 ^ b498 ^ c498;
  assign sub498 = a498 ^ b_inv498 ^ c498;
  assign and498 = a498 & b498;
  assign or498  = a498 | b498;
  assign c499 = (a498 & b498) | (a498 & c498) | (b498 & c498);
  wire c_sub499;
  assign c_sub499 = (a498 & b_inv498) | (a498 & c498) | (b_inv498 & c498);
  wire s499, sub499, and499, or499;
  wire b_inv499;
  assign b_inv499 = ~b499;
  assign s499  = a499 ^ b499 ^ c499;
  assign sub499 = a499 ^ b_inv499 ^ c499;
  assign and499 = a499 & b499;
  assign or499  = a499 | b499;
  assign c500 = (a499 & b499) | (a499 & c499) | (b499 & c499);
  wire c_sub500;
  assign c_sub500 = (a499 & b_inv499) | (a499 & c499) | (b_inv499 & c499);
  wire s500, sub500, and500, or500;
  wire b_inv500;
  assign b_inv500 = ~b500;
  assign s500  = a500 ^ b500 ^ c500;
  assign sub500 = a500 ^ b_inv500 ^ c500;
  assign and500 = a500 & b500;
  assign or500  = a500 | b500;
  assign c501 = (a500 & b500) | (a500 & c500) | (b500 & c500);
  wire c_sub501;
  assign c_sub501 = (a500 & b_inv500) | (a500 & c500) | (b_inv500 & c500);
  wire s501, sub501, and501, or501;
  wire b_inv501;
  assign b_inv501 = ~b501;
  assign s501  = a501 ^ b501 ^ c501;
  assign sub501 = a501 ^ b_inv501 ^ c501;
  assign and501 = a501 & b501;
  assign or501  = a501 | b501;
  assign c502 = (a501 & b501) | (a501 & c501) | (b501 & c501);
  wire c_sub502;
  assign c_sub502 = (a501 & b_inv501) | (a501 & c501) | (b_inv501 & c501);
  wire s502, sub502, and502, or502;
  wire b_inv502;
  assign b_inv502 = ~b502;
  assign s502  = a502 ^ b502 ^ c502;
  assign sub502 = a502 ^ b_inv502 ^ c502;
  assign and502 = a502 & b502;
  assign or502  = a502 | b502;
  assign c503 = (a502 & b502) | (a502 & c502) | (b502 & c502);
  wire c_sub503;
  assign c_sub503 = (a502 & b_inv502) | (a502 & c502) | (b_inv502 & c502);
  wire s503, sub503, and503, or503;
  wire b_inv503;
  assign b_inv503 = ~b503;
  assign s503  = a503 ^ b503 ^ c503;
  assign sub503 = a503 ^ b_inv503 ^ c503;
  assign and503 = a503 & b503;
  assign or503  = a503 | b503;
  assign c504 = (a503 & b503) | (a503 & c503) | (b503 & c503);
  wire c_sub504;
  assign c_sub504 = (a503 & b_inv503) | (a503 & c503) | (b_inv503 & c503);
  wire s504, sub504, and504, or504;
  wire b_inv504;
  assign b_inv504 = ~b504;
  assign s504  = a504 ^ b504 ^ c504;
  assign sub504 = a504 ^ b_inv504 ^ c504;
  assign and504 = a504 & b504;
  assign or504  = a504 | b504;
  assign c505 = (a504 & b504) | (a504 & c504) | (b504 & c504);
  wire c_sub505;
  assign c_sub505 = (a504 & b_inv504) | (a504 & c504) | (b_inv504 & c504);
  wire s505, sub505, and505, or505;
  wire b_inv505;
  assign b_inv505 = ~b505;
  assign s505  = a505 ^ b505 ^ c505;
  assign sub505 = a505 ^ b_inv505 ^ c505;
  assign and505 = a505 & b505;
  assign or505  = a505 | b505;
  assign c506 = (a505 & b505) | (a505 & c505) | (b505 & c505);
  wire c_sub506;
  assign c_sub506 = (a505 & b_inv505) | (a505 & c505) | (b_inv505 & c505);
  wire s506, sub506, and506, or506;
  wire b_inv506;
  assign b_inv506 = ~b506;
  assign s506  = a506 ^ b506 ^ c506;
  assign sub506 = a506 ^ b_inv506 ^ c506;
  assign and506 = a506 & b506;
  assign or506  = a506 | b506;
  assign c507 = (a506 & b506) | (a506 & c506) | (b506 & c506);
  wire c_sub507;
  assign c_sub507 = (a506 & b_inv506) | (a506 & c506) | (b_inv506 & c506);
  wire s507, sub507, and507, or507;
  wire b_inv507;
  assign b_inv507 = ~b507;
  assign s507  = a507 ^ b507 ^ c507;
  assign sub507 = a507 ^ b_inv507 ^ c507;
  assign and507 = a507 & b507;
  assign or507  = a507 | b507;
  assign c508 = (a507 & b507) | (a507 & c507) | (b507 & c507);
  wire c_sub508;
  assign c_sub508 = (a507 & b_inv507) | (a507 & c507) | (b_inv507 & c507);
  wire s508, sub508, and508, or508;
  wire b_inv508;
  assign b_inv508 = ~b508;
  assign s508  = a508 ^ b508 ^ c508;
  assign sub508 = a508 ^ b_inv508 ^ c508;
  assign and508 = a508 & b508;
  assign or508  = a508 | b508;
  assign c509 = (a508 & b508) | (a508 & c508) | (b508 & c508);
  wire c_sub509;
  assign c_sub509 = (a508 & b_inv508) | (a508 & c508) | (b_inv508 & c508);
  wire s509, sub509, and509, or509;
  wire b_inv509;
  assign b_inv509 = ~b509;
  assign s509  = a509 ^ b509 ^ c509;
  assign sub509 = a509 ^ b_inv509 ^ c509;
  assign and509 = a509 & b509;
  assign or509  = a509 | b509;
  assign c510 = (a509 & b509) | (a509 & c509) | (b509 & c509);
  wire c_sub510;
  assign c_sub510 = (a509 & b_inv509) | (a509 & c509) | (b_inv509 & c509);
  wire s510, sub510, and510, or510;
  wire b_inv510;
  assign b_inv510 = ~b510;
  assign s510  = a510 ^ b510 ^ c510;
  assign sub510 = a510 ^ b_inv510 ^ c510;
  assign and510 = a510 & b510;
  assign or510  = a510 | b510;
  assign c511 = (a510 & b510) | (a510 & c510) | (b510 & c510);
  wire c_sub511;
  assign c_sub511 = (a510 & b_inv510) | (a510 & c510) | (b_inv510 & c510);
  wire s511, sub511, and511, or511;
  wire b_inv511;
  assign b_inv511 = ~b511;
  assign s511  = a511 ^ b511 ^ c511;
  assign sub511 = a511 ^ b_inv511 ^ c511;
  assign and511 = a511 & b511;
  assign or511  = a511 | b511;
  assign c512 = (a511 & b511) | (a511 & c511) | (b511 & c511);
  wire c_sub512;
  assign c_sub512 = (a511 & b_inv511) | (a511 & c511) | (b_inv511 & c511);
  wire s512, sub512, and512, or512;
  wire b_inv512;
  assign b_inv512 = ~b512;
  assign s512  = a512 ^ b512 ^ c512;
  assign sub512 = a512 ^ b_inv512 ^ c512;
  assign and512 = a512 & b512;
  assign or512  = a512 | b512;
  assign c513 = (a512 & b512) | (a512 & c512) | (b512 & c512);
  wire c_sub513;
  assign c_sub513 = (a512 & b_inv512) | (a512 & c512) | (b_inv512 & c512);
  wire s513, sub513, and513, or513;
  wire b_inv513;
  assign b_inv513 = ~b513;
  assign s513  = a513 ^ b513 ^ c513;
  assign sub513 = a513 ^ b_inv513 ^ c513;
  assign and513 = a513 & b513;
  assign or513  = a513 | b513;
  assign c514 = (a513 & b513) | (a513 & c513) | (b513 & c513);
  wire c_sub514;
  assign c_sub514 = (a513 & b_inv513) | (a513 & c513) | (b_inv513 & c513);
  wire s514, sub514, and514, or514;
  wire b_inv514;
  assign b_inv514 = ~b514;
  assign s514  = a514 ^ b514 ^ c514;
  assign sub514 = a514 ^ b_inv514 ^ c514;
  assign and514 = a514 & b514;
  assign or514  = a514 | b514;
  assign c515 = (a514 & b514) | (a514 & c514) | (b514 & c514);
  wire c_sub515;
  assign c_sub515 = (a514 & b_inv514) | (a514 & c514) | (b_inv514 & c514);
  wire s515, sub515, and515, or515;
  wire b_inv515;
  assign b_inv515 = ~b515;
  assign s515  = a515 ^ b515 ^ c515;
  assign sub515 = a515 ^ b_inv515 ^ c515;
  assign and515 = a515 & b515;
  assign or515  = a515 | b515;
  assign c516 = (a515 & b515) | (a515 & c515) | (b515 & c515);
  wire c_sub516;
  assign c_sub516 = (a515 & b_inv515) | (a515 & c515) | (b_inv515 & c515);
  wire s516, sub516, and516, or516;
  wire b_inv516;
  assign b_inv516 = ~b516;
  assign s516  = a516 ^ b516 ^ c516;
  assign sub516 = a516 ^ b_inv516 ^ c516;
  assign and516 = a516 & b516;
  assign or516  = a516 | b516;
  assign c517 = (a516 & b516) | (a516 & c516) | (b516 & c516);
  wire c_sub517;
  assign c_sub517 = (a516 & b_inv516) | (a516 & c516) | (b_inv516 & c516);
  wire s517, sub517, and517, or517;
  wire b_inv517;
  assign b_inv517 = ~b517;
  assign s517  = a517 ^ b517 ^ c517;
  assign sub517 = a517 ^ b_inv517 ^ c517;
  assign and517 = a517 & b517;
  assign or517  = a517 | b517;
  assign c518 = (a517 & b517) | (a517 & c517) | (b517 & c517);
  wire c_sub518;
  assign c_sub518 = (a517 & b_inv517) | (a517 & c517) | (b_inv517 & c517);
  wire s518, sub518, and518, or518;
  wire b_inv518;
  assign b_inv518 = ~b518;
  assign s518  = a518 ^ b518 ^ c518;
  assign sub518 = a518 ^ b_inv518 ^ c518;
  assign and518 = a518 & b518;
  assign or518  = a518 | b518;
  assign c519 = (a518 & b518) | (a518 & c518) | (b518 & c518);
  wire c_sub519;
  assign c_sub519 = (a518 & b_inv518) | (a518 & c518) | (b_inv518 & c518);
  wire s519, sub519, and519, or519;
  wire b_inv519;
  assign b_inv519 = ~b519;
  assign s519  = a519 ^ b519 ^ c519;
  assign sub519 = a519 ^ b_inv519 ^ c519;
  assign and519 = a519 & b519;
  assign or519  = a519 | b519;
  assign c520 = (a519 & b519) | (a519 & c519) | (b519 & c519);
  wire c_sub520;
  assign c_sub520 = (a519 & b_inv519) | (a519 & c519) | (b_inv519 & c519);
  wire s520, sub520, and520, or520;
  wire b_inv520;
  assign b_inv520 = ~b520;
  assign s520  = a520 ^ b520 ^ c520;
  assign sub520 = a520 ^ b_inv520 ^ c520;
  assign and520 = a520 & b520;
  assign or520  = a520 | b520;
  assign c521 = (a520 & b520) | (a520 & c520) | (b520 & c520);
  wire c_sub521;
  assign c_sub521 = (a520 & b_inv520) | (a520 & c520) | (b_inv520 & c520);
  wire s521, sub521, and521, or521;
  wire b_inv521;
  assign b_inv521 = ~b521;
  assign s521  = a521 ^ b521 ^ c521;
  assign sub521 = a521 ^ b_inv521 ^ c521;
  assign and521 = a521 & b521;
  assign or521  = a521 | b521;
  assign c522 = (a521 & b521) | (a521 & c521) | (b521 & c521);
  wire c_sub522;
  assign c_sub522 = (a521 & b_inv521) | (a521 & c521) | (b_inv521 & c521);
  wire s522, sub522, and522, or522;
  wire b_inv522;
  assign b_inv522 = ~b522;
  assign s522  = a522 ^ b522 ^ c522;
  assign sub522 = a522 ^ b_inv522 ^ c522;
  assign and522 = a522 & b522;
  assign or522  = a522 | b522;
  assign c523 = (a522 & b522) | (a522 & c522) | (b522 & c522);
  wire c_sub523;
  assign c_sub523 = (a522 & b_inv522) | (a522 & c522) | (b_inv522 & c522);
  wire s523, sub523, and523, or523;
  wire b_inv523;
  assign b_inv523 = ~b523;
  assign s523  = a523 ^ b523 ^ c523;
  assign sub523 = a523 ^ b_inv523 ^ c523;
  assign and523 = a523 & b523;
  assign or523  = a523 | b523;
  assign c524 = (a523 & b523) | (a523 & c523) | (b523 & c523);
  wire c_sub524;
  assign c_sub524 = (a523 & b_inv523) | (a523 & c523) | (b_inv523 & c523);
  wire s524, sub524, and524, or524;
  wire b_inv524;
  assign b_inv524 = ~b524;
  assign s524  = a524 ^ b524 ^ c524;
  assign sub524 = a524 ^ b_inv524 ^ c524;
  assign and524 = a524 & b524;
  assign or524  = a524 | b524;
  assign c525 = (a524 & b524) | (a524 & c524) | (b524 & c524);
  wire c_sub525;
  assign c_sub525 = (a524 & b_inv524) | (a524 & c524) | (b_inv524 & c524);
  wire s525, sub525, and525, or525;
  wire b_inv525;
  assign b_inv525 = ~b525;
  assign s525  = a525 ^ b525 ^ c525;
  assign sub525 = a525 ^ b_inv525 ^ c525;
  assign and525 = a525 & b525;
  assign or525  = a525 | b525;
  assign c526 = (a525 & b525) | (a525 & c525) | (b525 & c525);
  wire c_sub526;
  assign c_sub526 = (a525 & b_inv525) | (a525 & c525) | (b_inv525 & c525);
  wire s526, sub526, and526, or526;
  wire b_inv526;
  assign b_inv526 = ~b526;
  assign s526  = a526 ^ b526 ^ c526;
  assign sub526 = a526 ^ b_inv526 ^ c526;
  assign and526 = a526 & b526;
  assign or526  = a526 | b526;
  assign c527 = (a526 & b526) | (a526 & c526) | (b526 & c526);
  wire c_sub527;
  assign c_sub527 = (a526 & b_inv526) | (a526 & c526) | (b_inv526 & c526);
  wire s527, sub527, and527, or527;
  wire b_inv527;
  assign b_inv527 = ~b527;
  assign s527  = a527 ^ b527 ^ c527;
  assign sub527 = a527 ^ b_inv527 ^ c527;
  assign and527 = a527 & b527;
  assign or527  = a527 | b527;
  assign c528 = (a527 & b527) | (a527 & c527) | (b527 & c527);
  wire c_sub528;
  assign c_sub528 = (a527 & b_inv527) | (a527 & c527) | (b_inv527 & c527);
  wire s528, sub528, and528, or528;
  wire b_inv528;
  assign b_inv528 = ~b528;
  assign s528  = a528 ^ b528 ^ c528;
  assign sub528 = a528 ^ b_inv528 ^ c528;
  assign and528 = a528 & b528;
  assign or528  = a528 | b528;
  assign c529 = (a528 & b528) | (a528 & c528) | (b528 & c528);
  wire c_sub529;
  assign c_sub529 = (a528 & b_inv528) | (a528 & c528) | (b_inv528 & c528);
  wire s529, sub529, and529, or529;
  wire b_inv529;
  assign b_inv529 = ~b529;
  assign s529  = a529 ^ b529 ^ c529;
  assign sub529 = a529 ^ b_inv529 ^ c529;
  assign and529 = a529 & b529;
  assign or529  = a529 | b529;
  assign c530 = (a529 & b529) | (a529 & c529) | (b529 & c529);
  wire c_sub530;
  assign c_sub530 = (a529 & b_inv529) | (a529 & c529) | (b_inv529 & c529);
  wire s530, sub530, and530, or530;
  wire b_inv530;
  assign b_inv530 = ~b530;
  assign s530  = a530 ^ b530 ^ c530;
  assign sub530 = a530 ^ b_inv530 ^ c530;
  assign and530 = a530 & b530;
  assign or530  = a530 | b530;
  assign c531 = (a530 & b530) | (a530 & c530) | (b530 & c530);
  wire c_sub531;
  assign c_sub531 = (a530 & b_inv530) | (a530 & c530) | (b_inv530 & c530);
  wire s531, sub531, and531, or531;
  wire b_inv531;
  assign b_inv531 = ~b531;
  assign s531  = a531 ^ b531 ^ c531;
  assign sub531 = a531 ^ b_inv531 ^ c531;
  assign and531 = a531 & b531;
  assign or531  = a531 | b531;
  assign c532 = (a531 & b531) | (a531 & c531) | (b531 & c531);
  wire c_sub532;
  assign c_sub532 = (a531 & b_inv531) | (a531 & c531) | (b_inv531 & c531);
  wire s532, sub532, and532, or532;
  wire b_inv532;
  assign b_inv532 = ~b532;
  assign s532  = a532 ^ b532 ^ c532;
  assign sub532 = a532 ^ b_inv532 ^ c532;
  assign and532 = a532 & b532;
  assign or532  = a532 | b532;
  assign c533 = (a532 & b532) | (a532 & c532) | (b532 & c532);
  wire c_sub533;
  assign c_sub533 = (a532 & b_inv532) | (a532 & c532) | (b_inv532 & c532);
  wire s533, sub533, and533, or533;
  wire b_inv533;
  assign b_inv533 = ~b533;
  assign s533  = a533 ^ b533 ^ c533;
  assign sub533 = a533 ^ b_inv533 ^ c533;
  assign and533 = a533 & b533;
  assign or533  = a533 | b533;
  assign c534 = (a533 & b533) | (a533 & c533) | (b533 & c533);
  wire c_sub534;
  assign c_sub534 = (a533 & b_inv533) | (a533 & c533) | (b_inv533 & c533);
  wire s534, sub534, and534, or534;
  wire b_inv534;
  assign b_inv534 = ~b534;
  assign s534  = a534 ^ b534 ^ c534;
  assign sub534 = a534 ^ b_inv534 ^ c534;
  assign and534 = a534 & b534;
  assign or534  = a534 | b534;
  assign c535 = (a534 & b534) | (a534 & c534) | (b534 & c534);
  wire c_sub535;
  assign c_sub535 = (a534 & b_inv534) | (a534 & c534) | (b_inv534 & c534);
  wire s535, sub535, and535, or535;
  wire b_inv535;
  assign b_inv535 = ~b535;
  assign s535  = a535 ^ b535 ^ c535;
  assign sub535 = a535 ^ b_inv535 ^ c535;
  assign and535 = a535 & b535;
  assign or535  = a535 | b535;
  assign c536 = (a535 & b535) | (a535 & c535) | (b535 & c535);
  wire c_sub536;
  assign c_sub536 = (a535 & b_inv535) | (a535 & c535) | (b_inv535 & c535);
  wire s536, sub536, and536, or536;
  wire b_inv536;
  assign b_inv536 = ~b536;
  assign s536  = a536 ^ b536 ^ c536;
  assign sub536 = a536 ^ b_inv536 ^ c536;
  assign and536 = a536 & b536;
  assign or536  = a536 | b536;
  assign c537 = (a536 & b536) | (a536 & c536) | (b536 & c536);
  wire c_sub537;
  assign c_sub537 = (a536 & b_inv536) | (a536 & c536) | (b_inv536 & c536);
  wire s537, sub537, and537, or537;
  wire b_inv537;
  assign b_inv537 = ~b537;
  assign s537  = a537 ^ b537 ^ c537;
  assign sub537 = a537 ^ b_inv537 ^ c537;
  assign and537 = a537 & b537;
  assign or537  = a537 | b537;
  assign c538 = (a537 & b537) | (a537 & c537) | (b537 & c537);
  wire c_sub538;
  assign c_sub538 = (a537 & b_inv537) | (a537 & c537) | (b_inv537 & c537);
  wire s538, sub538, and538, or538;
  wire b_inv538;
  assign b_inv538 = ~b538;
  assign s538  = a538 ^ b538 ^ c538;
  assign sub538 = a538 ^ b_inv538 ^ c538;
  assign and538 = a538 & b538;
  assign or538  = a538 | b538;
  assign c539 = (a538 & b538) | (a538 & c538) | (b538 & c538);
  wire c_sub539;
  assign c_sub539 = (a538 & b_inv538) | (a538 & c538) | (b_inv538 & c538);
  wire s539, sub539, and539, or539;
  wire b_inv539;
  assign b_inv539 = ~b539;
  assign s539  = a539 ^ b539 ^ c539;
  assign sub539 = a539 ^ b_inv539 ^ c539;
  assign and539 = a539 & b539;
  assign or539  = a539 | b539;
  assign c540 = (a539 & b539) | (a539 & c539) | (b539 & c539);
  wire c_sub540;
  assign c_sub540 = (a539 & b_inv539) | (a539 & c539) | (b_inv539 & c539);
  wire s540, sub540, and540, or540;
  wire b_inv540;
  assign b_inv540 = ~b540;
  assign s540  = a540 ^ b540 ^ c540;
  assign sub540 = a540 ^ b_inv540 ^ c540;
  assign and540 = a540 & b540;
  assign or540  = a540 | b540;
  assign c541 = (a540 & b540) | (a540 & c540) | (b540 & c540);
  wire c_sub541;
  assign c_sub541 = (a540 & b_inv540) | (a540 & c540) | (b_inv540 & c540);
  wire s541, sub541, and541, or541;
  wire b_inv541;
  assign b_inv541 = ~b541;
  assign s541  = a541 ^ b541 ^ c541;
  assign sub541 = a541 ^ b_inv541 ^ c541;
  assign and541 = a541 & b541;
  assign or541  = a541 | b541;
  assign c542 = (a541 & b541) | (a541 & c541) | (b541 & c541);
  wire c_sub542;
  assign c_sub542 = (a541 & b_inv541) | (a541 & c541) | (b_inv541 & c541);
  wire s542, sub542, and542, or542;
  wire b_inv542;
  assign b_inv542 = ~b542;
  assign s542  = a542 ^ b542 ^ c542;
  assign sub542 = a542 ^ b_inv542 ^ c542;
  assign and542 = a542 & b542;
  assign or542  = a542 | b542;
  assign c543 = (a542 & b542) | (a542 & c542) | (b542 & c542);
  wire c_sub543;
  assign c_sub543 = (a542 & b_inv542) | (a542 & c542) | (b_inv542 & c542);
  wire s543, sub543, and543, or543;
  wire b_inv543;
  assign b_inv543 = ~b543;
  assign s543  = a543 ^ b543 ^ c543;
  assign sub543 = a543 ^ b_inv543 ^ c543;
  assign and543 = a543 & b543;
  assign or543  = a543 | b543;
  assign c544 = (a543 & b543) | (a543 & c543) | (b543 & c543);
  wire c_sub544;
  assign c_sub544 = (a543 & b_inv543) | (a543 & c543) | (b_inv543 & c543);
  wire s544, sub544, and544, or544;
  wire b_inv544;
  assign b_inv544 = ~b544;
  assign s544  = a544 ^ b544 ^ c544;
  assign sub544 = a544 ^ b_inv544 ^ c544;
  assign and544 = a544 & b544;
  assign or544  = a544 | b544;
  assign c545 = (a544 & b544) | (a544 & c544) | (b544 & c544);
  wire c_sub545;
  assign c_sub545 = (a544 & b_inv544) | (a544 & c544) | (b_inv544 & c544);
  wire s545, sub545, and545, or545;
  wire b_inv545;
  assign b_inv545 = ~b545;
  assign s545  = a545 ^ b545 ^ c545;
  assign sub545 = a545 ^ b_inv545 ^ c545;
  assign and545 = a545 & b545;
  assign or545  = a545 | b545;
  assign c546 = (a545 & b545) | (a545 & c545) | (b545 & c545);
  wire c_sub546;
  assign c_sub546 = (a545 & b_inv545) | (a545 & c545) | (b_inv545 & c545);
  wire s546, sub546, and546, or546;
  wire b_inv546;
  assign b_inv546 = ~b546;
  assign s546  = a546 ^ b546 ^ c546;
  assign sub546 = a546 ^ b_inv546 ^ c546;
  assign and546 = a546 & b546;
  assign or546  = a546 | b546;
  assign c547 = (a546 & b546) | (a546 & c546) | (b546 & c546);
  wire c_sub547;
  assign c_sub547 = (a546 & b_inv546) | (a546 & c546) | (b_inv546 & c546);
  wire s547, sub547, and547, or547;
  wire b_inv547;
  assign b_inv547 = ~b547;
  assign s547  = a547 ^ b547 ^ c547;
  assign sub547 = a547 ^ b_inv547 ^ c547;
  assign and547 = a547 & b547;
  assign or547  = a547 | b547;
  assign c548 = (a547 & b547) | (a547 & c547) | (b547 & c547);
  wire c_sub548;
  assign c_sub548 = (a547 & b_inv547) | (a547 & c547) | (b_inv547 & c547);
  wire s548, sub548, and548, or548;
  wire b_inv548;
  assign b_inv548 = ~b548;
  assign s548  = a548 ^ b548 ^ c548;
  assign sub548 = a548 ^ b_inv548 ^ c548;
  assign and548 = a548 & b548;
  assign or548  = a548 | b548;
  assign c549 = (a548 & b548) | (a548 & c548) | (b548 & c548);
  wire c_sub549;
  assign c_sub549 = (a548 & b_inv548) | (a548 & c548) | (b_inv548 & c548);
  wire s549, sub549, and549, or549;
  wire b_inv549;
  assign b_inv549 = ~b549;
  assign s549  = a549 ^ b549 ^ c549;
  assign sub549 = a549 ^ b_inv549 ^ c549;
  assign and549 = a549 & b549;
  assign or549  = a549 | b549;
  assign c550 = (a549 & b549) | (a549 & c549) | (b549 & c549);
  wire c_sub550;
  assign c_sub550 = (a549 & b_inv549) | (a549 & c549) | (b_inv549 & c549);
  wire s550, sub550, and550, or550;
  wire b_inv550;
  assign b_inv550 = ~b550;
  assign s550  = a550 ^ b550 ^ c550;
  assign sub550 = a550 ^ b_inv550 ^ c550;
  assign and550 = a550 & b550;
  assign or550  = a550 | b550;
  assign c551 = (a550 & b550) | (a550 & c550) | (b550 & c550);
  wire c_sub551;
  assign c_sub551 = (a550 & b_inv550) | (a550 & c550) | (b_inv550 & c550);
  wire s551, sub551, and551, or551;
  wire b_inv551;
  assign b_inv551 = ~b551;
  assign s551  = a551 ^ b551 ^ c551;
  assign sub551 = a551 ^ b_inv551 ^ c551;
  assign and551 = a551 & b551;
  assign or551  = a551 | b551;
  assign c552 = (a551 & b551) | (a551 & c551) | (b551 & c551);
  wire c_sub552;
  assign c_sub552 = (a551 & b_inv551) | (a551 & c551) | (b_inv551 & c551);
  wire s552, sub552, and552, or552;
  wire b_inv552;
  assign b_inv552 = ~b552;
  assign s552  = a552 ^ b552 ^ c552;
  assign sub552 = a552 ^ b_inv552 ^ c552;
  assign and552 = a552 & b552;
  assign or552  = a552 | b552;
  assign c553 = (a552 & b552) | (a552 & c552) | (b552 & c552);
  wire c_sub553;
  assign c_sub553 = (a552 & b_inv552) | (a552 & c552) | (b_inv552 & c552);
  wire s553, sub553, and553, or553;
  wire b_inv553;
  assign b_inv553 = ~b553;
  assign s553  = a553 ^ b553 ^ c553;
  assign sub553 = a553 ^ b_inv553 ^ c553;
  assign and553 = a553 & b553;
  assign or553  = a553 | b553;
  assign c554 = (a553 & b553) | (a553 & c553) | (b553 & c553);
  wire c_sub554;
  assign c_sub554 = (a553 & b_inv553) | (a553 & c553) | (b_inv553 & c553);
  wire s554, sub554, and554, or554;
  wire b_inv554;
  assign b_inv554 = ~b554;
  assign s554  = a554 ^ b554 ^ c554;
  assign sub554 = a554 ^ b_inv554 ^ c554;
  assign and554 = a554 & b554;
  assign or554  = a554 | b554;
  assign c555 = (a554 & b554) | (a554 & c554) | (b554 & c554);
  wire c_sub555;
  assign c_sub555 = (a554 & b_inv554) | (a554 & c554) | (b_inv554 & c554);
  wire s555, sub555, and555, or555;
  wire b_inv555;
  assign b_inv555 = ~b555;
  assign s555  = a555 ^ b555 ^ c555;
  assign sub555 = a555 ^ b_inv555 ^ c555;
  assign and555 = a555 & b555;
  assign or555  = a555 | b555;
  assign c556 = (a555 & b555) | (a555 & c555) | (b555 & c555);
  wire c_sub556;
  assign c_sub556 = (a555 & b_inv555) | (a555 & c555) | (b_inv555 & c555);
  wire s556, sub556, and556, or556;
  wire b_inv556;
  assign b_inv556 = ~b556;
  assign s556  = a556 ^ b556 ^ c556;
  assign sub556 = a556 ^ b_inv556 ^ c556;
  assign and556 = a556 & b556;
  assign or556  = a556 | b556;
  assign c557 = (a556 & b556) | (a556 & c556) | (b556 & c556);
  wire c_sub557;
  assign c_sub557 = (a556 & b_inv556) | (a556 & c556) | (b_inv556 & c556);
  wire s557, sub557, and557, or557;
  wire b_inv557;
  assign b_inv557 = ~b557;
  assign s557  = a557 ^ b557 ^ c557;
  assign sub557 = a557 ^ b_inv557 ^ c557;
  assign and557 = a557 & b557;
  assign or557  = a557 | b557;
  assign c558 = (a557 & b557) | (a557 & c557) | (b557 & c557);
  wire c_sub558;
  assign c_sub558 = (a557 & b_inv557) | (a557 & c557) | (b_inv557 & c557);
  wire s558, sub558, and558, or558;
  wire b_inv558;
  assign b_inv558 = ~b558;
  assign s558  = a558 ^ b558 ^ c558;
  assign sub558 = a558 ^ b_inv558 ^ c558;
  assign and558 = a558 & b558;
  assign or558  = a558 | b558;
  assign c559 = (a558 & b558) | (a558 & c558) | (b558 & c558);
  wire c_sub559;
  assign c_sub559 = (a558 & b_inv558) | (a558 & c558) | (b_inv558 & c558);
  wire s559, sub559, and559, or559;
  wire b_inv559;
  assign b_inv559 = ~b559;
  assign s559  = a559 ^ b559 ^ c559;
  assign sub559 = a559 ^ b_inv559 ^ c559;
  assign and559 = a559 & b559;
  assign or559  = a559 | b559;
  assign c560 = (a559 & b559) | (a559 & c559) | (b559 & c559);
  wire c_sub560;
  assign c_sub560 = (a559 & b_inv559) | (a559 & c559) | (b_inv559 & c559);
  wire s560, sub560, and560, or560;
  wire b_inv560;
  assign b_inv560 = ~b560;
  assign s560  = a560 ^ b560 ^ c560;
  assign sub560 = a560 ^ b_inv560 ^ c560;
  assign and560 = a560 & b560;
  assign or560  = a560 | b560;
  assign c561 = (a560 & b560) | (a560 & c560) | (b560 & c560);
  wire c_sub561;
  assign c_sub561 = (a560 & b_inv560) | (a560 & c560) | (b_inv560 & c560);
  wire s561, sub561, and561, or561;
  wire b_inv561;
  assign b_inv561 = ~b561;
  assign s561  = a561 ^ b561 ^ c561;
  assign sub561 = a561 ^ b_inv561 ^ c561;
  assign and561 = a561 & b561;
  assign or561  = a561 | b561;
  assign c562 = (a561 & b561) | (a561 & c561) | (b561 & c561);
  wire c_sub562;
  assign c_sub562 = (a561 & b_inv561) | (a561 & c561) | (b_inv561 & c561);
  wire s562, sub562, and562, or562;
  wire b_inv562;
  assign b_inv562 = ~b562;
  assign s562  = a562 ^ b562 ^ c562;
  assign sub562 = a562 ^ b_inv562 ^ c562;
  assign and562 = a562 & b562;
  assign or562  = a562 | b562;
  assign c563 = (a562 & b562) | (a562 & c562) | (b562 & c562);
  wire c_sub563;
  assign c_sub563 = (a562 & b_inv562) | (a562 & c562) | (b_inv562 & c562);
  wire s563, sub563, and563, or563;
  wire b_inv563;
  assign b_inv563 = ~b563;
  assign s563  = a563 ^ b563 ^ c563;
  assign sub563 = a563 ^ b_inv563 ^ c563;
  assign and563 = a563 & b563;
  assign or563  = a563 | b563;
  assign c564 = (a563 & b563) | (a563 & c563) | (b563 & c563);
  wire c_sub564;
  assign c_sub564 = (a563 & b_inv563) | (a563 & c563) | (b_inv563 & c563);
  wire s564, sub564, and564, or564;
  wire b_inv564;
  assign b_inv564 = ~b564;
  assign s564  = a564 ^ b564 ^ c564;
  assign sub564 = a564 ^ b_inv564 ^ c564;
  assign and564 = a564 & b564;
  assign or564  = a564 | b564;
  assign c565 = (a564 & b564) | (a564 & c564) | (b564 & c564);
  wire c_sub565;
  assign c_sub565 = (a564 & b_inv564) | (a564 & c564) | (b_inv564 & c564);
  wire s565, sub565, and565, or565;
  wire b_inv565;
  assign b_inv565 = ~b565;
  assign s565  = a565 ^ b565 ^ c565;
  assign sub565 = a565 ^ b_inv565 ^ c565;
  assign and565 = a565 & b565;
  assign or565  = a565 | b565;
  assign c566 = (a565 & b565) | (a565 & c565) | (b565 & c565);
  wire c_sub566;
  assign c_sub566 = (a565 & b_inv565) | (a565 & c565) | (b_inv565 & c565);
  wire s566, sub566, and566, or566;
  wire b_inv566;
  assign b_inv566 = ~b566;
  assign s566  = a566 ^ b566 ^ c566;
  assign sub566 = a566 ^ b_inv566 ^ c566;
  assign and566 = a566 & b566;
  assign or566  = a566 | b566;
  assign c567 = (a566 & b566) | (a566 & c566) | (b566 & c566);
  wire c_sub567;
  assign c_sub567 = (a566 & b_inv566) | (a566 & c566) | (b_inv566 & c566);
  wire s567, sub567, and567, or567;
  wire b_inv567;
  assign b_inv567 = ~b567;
  assign s567  = a567 ^ b567 ^ c567;
  assign sub567 = a567 ^ b_inv567 ^ c567;
  assign and567 = a567 & b567;
  assign or567  = a567 | b567;
  assign c568 = (a567 & b567) | (a567 & c567) | (b567 & c567);
  wire c_sub568;
  assign c_sub568 = (a567 & b_inv567) | (a567 & c567) | (b_inv567 & c567);
  wire s568, sub568, and568, or568;
  wire b_inv568;
  assign b_inv568 = ~b568;
  assign s568  = a568 ^ b568 ^ c568;
  assign sub568 = a568 ^ b_inv568 ^ c568;
  assign and568 = a568 & b568;
  assign or568  = a568 | b568;
  assign c569 = (a568 & b568) | (a568 & c568) | (b568 & c568);
  wire c_sub569;
  assign c_sub569 = (a568 & b_inv568) | (a568 & c568) | (b_inv568 & c568);
  wire s569, sub569, and569, or569;
  wire b_inv569;
  assign b_inv569 = ~b569;
  assign s569  = a569 ^ b569 ^ c569;
  assign sub569 = a569 ^ b_inv569 ^ c569;
  assign and569 = a569 & b569;
  assign or569  = a569 | b569;
  assign c570 = (a569 & b569) | (a569 & c569) | (b569 & c569);
  wire c_sub570;
  assign c_sub570 = (a569 & b_inv569) | (a569 & c569) | (b_inv569 & c569);
  wire s570, sub570, and570, or570;
  wire b_inv570;
  assign b_inv570 = ~b570;
  assign s570  = a570 ^ b570 ^ c570;
  assign sub570 = a570 ^ b_inv570 ^ c570;
  assign and570 = a570 & b570;
  assign or570  = a570 | b570;
  assign c571 = (a570 & b570) | (a570 & c570) | (b570 & c570);
  wire c_sub571;
  assign c_sub571 = (a570 & b_inv570) | (a570 & c570) | (b_inv570 & c570);
  wire s571, sub571, and571, or571;
  wire b_inv571;
  assign b_inv571 = ~b571;
  assign s571  = a571 ^ b571 ^ c571;
  assign sub571 = a571 ^ b_inv571 ^ c571;
  assign and571 = a571 & b571;
  assign or571  = a571 | b571;
  assign c572 = (a571 & b571) | (a571 & c571) | (b571 & c571);
  wire c_sub572;
  assign c_sub572 = (a571 & b_inv571) | (a571 & c571) | (b_inv571 & c571);
  wire s572, sub572, and572, or572;
  wire b_inv572;
  assign b_inv572 = ~b572;
  assign s572  = a572 ^ b572 ^ c572;
  assign sub572 = a572 ^ b_inv572 ^ c572;
  assign and572 = a572 & b572;
  assign or572  = a572 | b572;
  assign c573 = (a572 & b572) | (a572 & c572) | (b572 & c572);
  wire c_sub573;
  assign c_sub573 = (a572 & b_inv572) | (a572 & c572) | (b_inv572 & c572);
  wire s573, sub573, and573, or573;
  wire b_inv573;
  assign b_inv573 = ~b573;
  assign s573  = a573 ^ b573 ^ c573;
  assign sub573 = a573 ^ b_inv573 ^ c573;
  assign and573 = a573 & b573;
  assign or573  = a573 | b573;
  assign c574 = (a573 & b573) | (a573 & c573) | (b573 & c573);
  wire c_sub574;
  assign c_sub574 = (a573 & b_inv573) | (a573 & c573) | (b_inv573 & c573);
  wire s574, sub574, and574, or574;
  wire b_inv574;
  assign b_inv574 = ~b574;
  assign s574  = a574 ^ b574 ^ c574;
  assign sub574 = a574 ^ b_inv574 ^ c574;
  assign and574 = a574 & b574;
  assign or574  = a574 | b574;
  assign c575 = (a574 & b574) | (a574 & c574) | (b574 & c574);
  wire c_sub575;
  assign c_sub575 = (a574 & b_inv574) | (a574 & c574) | (b_inv574 & c574);
  wire s575, sub575, and575, or575;
  wire b_inv575;
  assign b_inv575 = ~b575;
  assign s575  = a575 ^ b575 ^ c575;
  assign sub575 = a575 ^ b_inv575 ^ c575;
  assign and575 = a575 & b575;
  assign or575  = a575 | b575;
  assign c576 = (a575 & b575) | (a575 & c575) | (b575 & c575);
  wire c_sub576;
  assign c_sub576 = (a575 & b_inv575) | (a575 & c575) | (b_inv575 & c575);
  wire s576, sub576, and576, or576;
  wire b_inv576;
  assign b_inv576 = ~b576;
  assign s576  = a576 ^ b576 ^ c576;
  assign sub576 = a576 ^ b_inv576 ^ c576;
  assign and576 = a576 & b576;
  assign or576  = a576 | b576;
  assign c577 = (a576 & b576) | (a576 & c576) | (b576 & c576);
  wire c_sub577;
  assign c_sub577 = (a576 & b_inv576) | (a576 & c576) | (b_inv576 & c576);
  wire s577, sub577, and577, or577;
  wire b_inv577;
  assign b_inv577 = ~b577;
  assign s577  = a577 ^ b577 ^ c577;
  assign sub577 = a577 ^ b_inv577 ^ c577;
  assign and577 = a577 & b577;
  assign or577  = a577 | b577;
  assign c578 = (a577 & b577) | (a577 & c577) | (b577 & c577);
  wire c_sub578;
  assign c_sub578 = (a577 & b_inv577) | (a577 & c577) | (b_inv577 & c577);
  wire s578, sub578, and578, or578;
  wire b_inv578;
  assign b_inv578 = ~b578;
  assign s578  = a578 ^ b578 ^ c578;
  assign sub578 = a578 ^ b_inv578 ^ c578;
  assign and578 = a578 & b578;
  assign or578  = a578 | b578;
  assign c579 = (a578 & b578) | (a578 & c578) | (b578 & c578);
  wire c_sub579;
  assign c_sub579 = (a578 & b_inv578) | (a578 & c578) | (b_inv578 & c578);
  wire s579, sub579, and579, or579;
  wire b_inv579;
  assign b_inv579 = ~b579;
  assign s579  = a579 ^ b579 ^ c579;
  assign sub579 = a579 ^ b_inv579 ^ c579;
  assign and579 = a579 & b579;
  assign or579  = a579 | b579;
  assign c580 = (a579 & b579) | (a579 & c579) | (b579 & c579);
  wire c_sub580;
  assign c_sub580 = (a579 & b_inv579) | (a579 & c579) | (b_inv579 & c579);
  wire s580, sub580, and580, or580;
  wire b_inv580;
  assign b_inv580 = ~b580;
  assign s580  = a580 ^ b580 ^ c580;
  assign sub580 = a580 ^ b_inv580 ^ c580;
  assign and580 = a580 & b580;
  assign or580  = a580 | b580;
  assign c581 = (a580 & b580) | (a580 & c580) | (b580 & c580);
  wire c_sub581;
  assign c_sub581 = (a580 & b_inv580) | (a580 & c580) | (b_inv580 & c580);
  wire s581, sub581, and581, or581;
  wire b_inv581;
  assign b_inv581 = ~b581;
  assign s581  = a581 ^ b581 ^ c581;
  assign sub581 = a581 ^ b_inv581 ^ c581;
  assign and581 = a581 & b581;
  assign or581  = a581 | b581;
  assign c582 = (a581 & b581) | (a581 & c581) | (b581 & c581);
  wire c_sub582;
  assign c_sub582 = (a581 & b_inv581) | (a581 & c581) | (b_inv581 & c581);
  wire s582, sub582, and582, or582;
  wire b_inv582;
  assign b_inv582 = ~b582;
  assign s582  = a582 ^ b582 ^ c582;
  assign sub582 = a582 ^ b_inv582 ^ c582;
  assign and582 = a582 & b582;
  assign or582  = a582 | b582;
  assign c583 = (a582 & b582) | (a582 & c582) | (b582 & c582);
  wire c_sub583;
  assign c_sub583 = (a582 & b_inv582) | (a582 & c582) | (b_inv582 & c582);
  wire s583, sub583, and583, or583;
  wire b_inv583;
  assign b_inv583 = ~b583;
  assign s583  = a583 ^ b583 ^ c583;
  assign sub583 = a583 ^ b_inv583 ^ c583;
  assign and583 = a583 & b583;
  assign or583  = a583 | b583;
  assign c584 = (a583 & b583) | (a583 & c583) | (b583 & c583);
  wire c_sub584;
  assign c_sub584 = (a583 & b_inv583) | (a583 & c583) | (b_inv583 & c583);
  wire s584, sub584, and584, or584;
  wire b_inv584;
  assign b_inv584 = ~b584;
  assign s584  = a584 ^ b584 ^ c584;
  assign sub584 = a584 ^ b_inv584 ^ c584;
  assign and584 = a584 & b584;
  assign or584  = a584 | b584;
  assign c585 = (a584 & b584) | (a584 & c584) | (b584 & c584);
  wire c_sub585;
  assign c_sub585 = (a584 & b_inv584) | (a584 & c584) | (b_inv584 & c584);
  wire s585, sub585, and585, or585;
  wire b_inv585;
  assign b_inv585 = ~b585;
  assign s585  = a585 ^ b585 ^ c585;
  assign sub585 = a585 ^ b_inv585 ^ c585;
  assign and585 = a585 & b585;
  assign or585  = a585 | b585;
  assign c586 = (a585 & b585) | (a585 & c585) | (b585 & c585);
  wire c_sub586;
  assign c_sub586 = (a585 & b_inv585) | (a585 & c585) | (b_inv585 & c585);
  wire s586, sub586, and586, or586;
  wire b_inv586;
  assign b_inv586 = ~b586;
  assign s586  = a586 ^ b586 ^ c586;
  assign sub586 = a586 ^ b_inv586 ^ c586;
  assign and586 = a586 & b586;
  assign or586  = a586 | b586;
  assign c587 = (a586 & b586) | (a586 & c586) | (b586 & c586);
  wire c_sub587;
  assign c_sub587 = (a586 & b_inv586) | (a586 & c586) | (b_inv586 & c586);
  wire s587, sub587, and587, or587;
  wire b_inv587;
  assign b_inv587 = ~b587;
  assign s587  = a587 ^ b587 ^ c587;
  assign sub587 = a587 ^ b_inv587 ^ c587;
  assign and587 = a587 & b587;
  assign or587  = a587 | b587;
  assign c588 = (a587 & b587) | (a587 & c587) | (b587 & c587);
  wire c_sub588;
  assign c_sub588 = (a587 & b_inv587) | (a587 & c587) | (b_inv587 & c587);
  wire s588, sub588, and588, or588;
  wire b_inv588;
  assign b_inv588 = ~b588;
  assign s588  = a588 ^ b588 ^ c588;
  assign sub588 = a588 ^ b_inv588 ^ c588;
  assign and588 = a588 & b588;
  assign or588  = a588 | b588;
  assign c589 = (a588 & b588) | (a588 & c588) | (b588 & c588);
  wire c_sub589;
  assign c_sub589 = (a588 & b_inv588) | (a588 & c588) | (b_inv588 & c588);
  wire s589, sub589, and589, or589;
  wire b_inv589;
  assign b_inv589 = ~b589;
  assign s589  = a589 ^ b589 ^ c589;
  assign sub589 = a589 ^ b_inv589 ^ c589;
  assign and589 = a589 & b589;
  assign or589  = a589 | b589;
  assign c590 = (a589 & b589) | (a589 & c589) | (b589 & c589);
  wire c_sub590;
  assign c_sub590 = (a589 & b_inv589) | (a589 & c589) | (b_inv589 & c589);
  wire s590, sub590, and590, or590;
  wire b_inv590;
  assign b_inv590 = ~b590;
  assign s590  = a590 ^ b590 ^ c590;
  assign sub590 = a590 ^ b_inv590 ^ c590;
  assign and590 = a590 & b590;
  assign or590  = a590 | b590;
  assign c591 = (a590 & b590) | (a590 & c590) | (b590 & c590);
  wire c_sub591;
  assign c_sub591 = (a590 & b_inv590) | (a590 & c590) | (b_inv590 & c590);
  wire s591, sub591, and591, or591;
  wire b_inv591;
  assign b_inv591 = ~b591;
  assign s591  = a591 ^ b591 ^ c591;
  assign sub591 = a591 ^ b_inv591 ^ c591;
  assign and591 = a591 & b591;
  assign or591  = a591 | b591;
  assign c592 = (a591 & b591) | (a591 & c591) | (b591 & c591);
  wire c_sub592;
  assign c_sub592 = (a591 & b_inv591) | (a591 & c591) | (b_inv591 & c591);
  wire s592, sub592, and592, or592;
  wire b_inv592;
  assign b_inv592 = ~b592;
  assign s592  = a592 ^ b592 ^ c592;
  assign sub592 = a592 ^ b_inv592 ^ c592;
  assign and592 = a592 & b592;
  assign or592  = a592 | b592;
  assign c593 = (a592 & b592) | (a592 & c592) | (b592 & c592);
  wire c_sub593;
  assign c_sub593 = (a592 & b_inv592) | (a592 & c592) | (b_inv592 & c592);
  wire s593, sub593, and593, or593;
  wire b_inv593;
  assign b_inv593 = ~b593;
  assign s593  = a593 ^ b593 ^ c593;
  assign sub593 = a593 ^ b_inv593 ^ c593;
  assign and593 = a593 & b593;
  assign or593  = a593 | b593;
  assign c594 = (a593 & b593) | (a593 & c593) | (b593 & c593);
  wire c_sub594;
  assign c_sub594 = (a593 & b_inv593) | (a593 & c593) | (b_inv593 & c593);
  wire s594, sub594, and594, or594;
  wire b_inv594;
  assign b_inv594 = ~b594;
  assign s594  = a594 ^ b594 ^ c594;
  assign sub594 = a594 ^ b_inv594 ^ c594;
  assign and594 = a594 & b594;
  assign or594  = a594 | b594;
  assign c595 = (a594 & b594) | (a594 & c594) | (b594 & c594);
  wire c_sub595;
  assign c_sub595 = (a594 & b_inv594) | (a594 & c594) | (b_inv594 & c594);
  wire s595, sub595, and595, or595;
  wire b_inv595;
  assign b_inv595 = ~b595;
  assign s595  = a595 ^ b595 ^ c595;
  assign sub595 = a595 ^ b_inv595 ^ c595;
  assign and595 = a595 & b595;
  assign or595  = a595 | b595;
  assign c596 = (a595 & b595) | (a595 & c595) | (b595 & c595);
  wire c_sub596;
  assign c_sub596 = (a595 & b_inv595) | (a595 & c595) | (b_inv595 & c595);
  wire s596, sub596, and596, or596;
  wire b_inv596;
  assign b_inv596 = ~b596;
  assign s596  = a596 ^ b596 ^ c596;
  assign sub596 = a596 ^ b_inv596 ^ c596;
  assign and596 = a596 & b596;
  assign or596  = a596 | b596;
  assign c597 = (a596 & b596) | (a596 & c596) | (b596 & c596);
  wire c_sub597;
  assign c_sub597 = (a596 & b_inv596) | (a596 & c596) | (b_inv596 & c596);
  wire s597, sub597, and597, or597;
  wire b_inv597;
  assign b_inv597 = ~b597;
  assign s597  = a597 ^ b597 ^ c597;
  assign sub597 = a597 ^ b_inv597 ^ c597;
  assign and597 = a597 & b597;
  assign or597  = a597 | b597;
  assign c598 = (a597 & b597) | (a597 & c597) | (b597 & c597);
  wire c_sub598;
  assign c_sub598 = (a597 & b_inv597) | (a597 & c597) | (b_inv597 & c597);
  wire s598, sub598, and598, or598;
  wire b_inv598;
  assign b_inv598 = ~b598;
  assign s598  = a598 ^ b598 ^ c598;
  assign sub598 = a598 ^ b_inv598 ^ c598;
  assign and598 = a598 & b598;
  assign or598  = a598 | b598;
  assign c599 = (a598 & b598) | (a598 & c598) | (b598 & c598);
  wire c_sub599;
  assign c_sub599 = (a598 & b_inv598) | (a598 & c598) | (b_inv598 & c598);
  wire s599, sub599, and599, or599;
  wire b_inv599;
  assign b_inv599 = ~b599;
  assign s599  = a599 ^ b599 ^ c599;
  assign sub599 = a599 ^ b_inv599 ^ c599;
  assign and599 = a599 & b599;
  assign or599  = a599 | b599;
  assign c600 = (a599 & b599) | (a599 & c599) | (b599 & c599);
  wire c_sub600;
  assign c_sub600 = (a599 & b_inv599) | (a599 & c599) | (b_inv599 & c599);
  wire s600, sub600, and600, or600;
  wire b_inv600;
  assign b_inv600 = ~b600;
  assign s600  = a600 ^ b600 ^ c600;
  assign sub600 = a600 ^ b_inv600 ^ c600;
  assign and600 = a600 & b600;
  assign or600  = a600 | b600;
  assign c601 = (a600 & b600) | (a600 & c600) | (b600 & c600);
  wire c_sub601;
  assign c_sub601 = (a600 & b_inv600) | (a600 & c600) | (b_inv600 & c600);
  wire s601, sub601, and601, or601;
  wire b_inv601;
  assign b_inv601 = ~b601;
  assign s601  = a601 ^ b601 ^ c601;
  assign sub601 = a601 ^ b_inv601 ^ c601;
  assign and601 = a601 & b601;
  assign or601  = a601 | b601;
  assign c602 = (a601 & b601) | (a601 & c601) | (b601 & c601);
  wire c_sub602;
  assign c_sub602 = (a601 & b_inv601) | (a601 & c601) | (b_inv601 & c601);
  wire s602, sub602, and602, or602;
  wire b_inv602;
  assign b_inv602 = ~b602;
  assign s602  = a602 ^ b602 ^ c602;
  assign sub602 = a602 ^ b_inv602 ^ c602;
  assign and602 = a602 & b602;
  assign or602  = a602 | b602;
  assign c603 = (a602 & b602) | (a602 & c602) | (b602 & c602);
  wire c_sub603;
  assign c_sub603 = (a602 & b_inv602) | (a602 & c602) | (b_inv602 & c602);
  wire s603, sub603, and603, or603;
  wire b_inv603;
  assign b_inv603 = ~b603;
  assign s603  = a603 ^ b603 ^ c603;
  assign sub603 = a603 ^ b_inv603 ^ c603;
  assign and603 = a603 & b603;
  assign or603  = a603 | b603;
  assign c604 = (a603 & b603) | (a603 & c603) | (b603 & c603);
  wire c_sub604;
  assign c_sub604 = (a603 & b_inv603) | (a603 & c603) | (b_inv603 & c603);
  wire s604, sub604, and604, or604;
  wire b_inv604;
  assign b_inv604 = ~b604;
  assign s604  = a604 ^ b604 ^ c604;
  assign sub604 = a604 ^ b_inv604 ^ c604;
  assign and604 = a604 & b604;
  assign or604  = a604 | b604;
  assign c605 = (a604 & b604) | (a604 & c604) | (b604 & c604);
  wire c_sub605;
  assign c_sub605 = (a604 & b_inv604) | (a604 & c604) | (b_inv604 & c604);
  wire s605, sub605, and605, or605;
  wire b_inv605;
  assign b_inv605 = ~b605;
  assign s605  = a605 ^ b605 ^ c605;
  assign sub605 = a605 ^ b_inv605 ^ c605;
  assign and605 = a605 & b605;
  assign or605  = a605 | b605;
  assign c606 = (a605 & b605) | (a605 & c605) | (b605 & c605);
  wire c_sub606;
  assign c_sub606 = (a605 & b_inv605) | (a605 & c605) | (b_inv605 & c605);
  wire s606, sub606, and606, or606;
  wire b_inv606;
  assign b_inv606 = ~b606;
  assign s606  = a606 ^ b606 ^ c606;
  assign sub606 = a606 ^ b_inv606 ^ c606;
  assign and606 = a606 & b606;
  assign or606  = a606 | b606;
  assign c607 = (a606 & b606) | (a606 & c606) | (b606 & c606);
  wire c_sub607;
  assign c_sub607 = (a606 & b_inv606) | (a606 & c606) | (b_inv606 & c606);
  wire s607, sub607, and607, or607;
  wire b_inv607;
  assign b_inv607 = ~b607;
  assign s607  = a607 ^ b607 ^ c607;
  assign sub607 = a607 ^ b_inv607 ^ c607;
  assign and607 = a607 & b607;
  assign or607  = a607 | b607;
  assign c608 = (a607 & b607) | (a607 & c607) | (b607 & c607);
  wire c_sub608;
  assign c_sub608 = (a607 & b_inv607) | (a607 & c607) | (b_inv607 & c607);
  wire s608, sub608, and608, or608;
  wire b_inv608;
  assign b_inv608 = ~b608;
  assign s608  = a608 ^ b608 ^ c608;
  assign sub608 = a608 ^ b_inv608 ^ c608;
  assign and608 = a608 & b608;
  assign or608  = a608 | b608;
  assign c609 = (a608 & b608) | (a608 & c608) | (b608 & c608);
  wire c_sub609;
  assign c_sub609 = (a608 & b_inv608) | (a608 & c608) | (b_inv608 & c608);
  wire s609, sub609, and609, or609;
  wire b_inv609;
  assign b_inv609 = ~b609;
  assign s609  = a609 ^ b609 ^ c609;
  assign sub609 = a609 ^ b_inv609 ^ c609;
  assign and609 = a609 & b609;
  assign or609  = a609 | b609;
  assign c610 = (a609 & b609) | (a609 & c609) | (b609 & c609);
  wire c_sub610;
  assign c_sub610 = (a609 & b_inv609) | (a609 & c609) | (b_inv609 & c609);
  wire s610, sub610, and610, or610;
  wire b_inv610;
  assign b_inv610 = ~b610;
  assign s610  = a610 ^ b610 ^ c610;
  assign sub610 = a610 ^ b_inv610 ^ c610;
  assign and610 = a610 & b610;
  assign or610  = a610 | b610;
  assign c611 = (a610 & b610) | (a610 & c610) | (b610 & c610);
  wire c_sub611;
  assign c_sub611 = (a610 & b_inv610) | (a610 & c610) | (b_inv610 & c610);
  wire s611, sub611, and611, or611;
  wire b_inv611;
  assign b_inv611 = ~b611;
  assign s611  = a611 ^ b611 ^ c611;
  assign sub611 = a611 ^ b_inv611 ^ c611;
  assign and611 = a611 & b611;
  assign or611  = a611 | b611;
  assign c612 = (a611 & b611) | (a611 & c611) | (b611 & c611);
  wire c_sub612;
  assign c_sub612 = (a611 & b_inv611) | (a611 & c611) | (b_inv611 & c611);
  wire s612, sub612, and612, or612;
  wire b_inv612;
  assign b_inv612 = ~b612;
  assign s612  = a612 ^ b612 ^ c612;
  assign sub612 = a612 ^ b_inv612 ^ c612;
  assign and612 = a612 & b612;
  assign or612  = a612 | b612;
  assign c613 = (a612 & b612) | (a612 & c612) | (b612 & c612);
  wire c_sub613;
  assign c_sub613 = (a612 & b_inv612) | (a612 & c612) | (b_inv612 & c612);
  wire s613, sub613, and613, or613;
  wire b_inv613;
  assign b_inv613 = ~b613;
  assign s613  = a613 ^ b613 ^ c613;
  assign sub613 = a613 ^ b_inv613 ^ c613;
  assign and613 = a613 & b613;
  assign or613  = a613 | b613;
  assign c614 = (a613 & b613) | (a613 & c613) | (b613 & c613);
  wire c_sub614;
  assign c_sub614 = (a613 & b_inv613) | (a613 & c613) | (b_inv613 & c613);
  wire s614, sub614, and614, or614;
  wire b_inv614;
  assign b_inv614 = ~b614;
  assign s614  = a614 ^ b614 ^ c614;
  assign sub614 = a614 ^ b_inv614 ^ c614;
  assign and614 = a614 & b614;
  assign or614  = a614 | b614;
  assign c615 = (a614 & b614) | (a614 & c614) | (b614 & c614);
  wire c_sub615;
  assign c_sub615 = (a614 & b_inv614) | (a614 & c614) | (b_inv614 & c614);
  wire s615, sub615, and615, or615;
  wire b_inv615;
  assign b_inv615 = ~b615;
  assign s615  = a615 ^ b615 ^ c615;
  assign sub615 = a615 ^ b_inv615 ^ c615;
  assign and615 = a615 & b615;
  assign or615  = a615 | b615;
  assign c616 = (a615 & b615) | (a615 & c615) | (b615 & c615);
  wire c_sub616;
  assign c_sub616 = (a615 & b_inv615) | (a615 & c615) | (b_inv615 & c615);
  wire s616, sub616, and616, or616;
  wire b_inv616;
  assign b_inv616 = ~b616;
  assign s616  = a616 ^ b616 ^ c616;
  assign sub616 = a616 ^ b_inv616 ^ c616;
  assign and616 = a616 & b616;
  assign or616  = a616 | b616;
  assign c617 = (a616 & b616) | (a616 & c616) | (b616 & c616);
  wire c_sub617;
  assign c_sub617 = (a616 & b_inv616) | (a616 & c616) | (b_inv616 & c616);
  wire s617, sub617, and617, or617;
  wire b_inv617;
  assign b_inv617 = ~b617;
  assign s617  = a617 ^ b617 ^ c617;
  assign sub617 = a617 ^ b_inv617 ^ c617;
  assign and617 = a617 & b617;
  assign or617  = a617 | b617;
  assign c618 = (a617 & b617) | (a617 & c617) | (b617 & c617);
  wire c_sub618;
  assign c_sub618 = (a617 & b_inv617) | (a617 & c617) | (b_inv617 & c617);
  wire s618, sub618, and618, or618;
  wire b_inv618;
  assign b_inv618 = ~b618;
  assign s618  = a618 ^ b618 ^ c618;
  assign sub618 = a618 ^ b_inv618 ^ c618;
  assign and618 = a618 & b618;
  assign or618  = a618 | b618;
  assign c619 = (a618 & b618) | (a618 & c618) | (b618 & c618);
  wire c_sub619;
  assign c_sub619 = (a618 & b_inv618) | (a618 & c618) | (b_inv618 & c618);
  wire s619, sub619, and619, or619;
  wire b_inv619;
  assign b_inv619 = ~b619;
  assign s619  = a619 ^ b619 ^ c619;
  assign sub619 = a619 ^ b_inv619 ^ c619;
  assign and619 = a619 & b619;
  assign or619  = a619 | b619;
  assign c620 = (a619 & b619) | (a619 & c619) | (b619 & c619);
  wire c_sub620;
  assign c_sub620 = (a619 & b_inv619) | (a619 & c619) | (b_inv619 & c619);
  wire s620, sub620, and620, or620;
  wire b_inv620;
  assign b_inv620 = ~b620;
  assign s620  = a620 ^ b620 ^ c620;
  assign sub620 = a620 ^ b_inv620 ^ c620;
  assign and620 = a620 & b620;
  assign or620  = a620 | b620;
  assign c621 = (a620 & b620) | (a620 & c620) | (b620 & c620);
  wire c_sub621;
  assign c_sub621 = (a620 & b_inv620) | (a620 & c620) | (b_inv620 & c620);
  wire s621, sub621, and621, or621;
  wire b_inv621;
  assign b_inv621 = ~b621;
  assign s621  = a621 ^ b621 ^ c621;
  assign sub621 = a621 ^ b_inv621 ^ c621;
  assign and621 = a621 & b621;
  assign or621  = a621 | b621;
  assign c622 = (a621 & b621) | (a621 & c621) | (b621 & c621);
  wire c_sub622;
  assign c_sub622 = (a621 & b_inv621) | (a621 & c621) | (b_inv621 & c621);
  wire s622, sub622, and622, or622;
  wire b_inv622;
  assign b_inv622 = ~b622;
  assign s622  = a622 ^ b622 ^ c622;
  assign sub622 = a622 ^ b_inv622 ^ c622;
  assign and622 = a622 & b622;
  assign or622  = a622 | b622;
  assign c623 = (a622 & b622) | (a622 & c622) | (b622 & c622);
  wire c_sub623;
  assign c_sub623 = (a622 & b_inv622) | (a622 & c622) | (b_inv622 & c622);
  wire s623, sub623, and623, or623;
  wire b_inv623;
  assign b_inv623 = ~b623;
  assign s623  = a623 ^ b623 ^ c623;
  assign sub623 = a623 ^ b_inv623 ^ c623;
  assign and623 = a623 & b623;
  assign or623  = a623 | b623;
  assign c624 = (a623 & b623) | (a623 & c623) | (b623 & c623);
  wire c_sub624;
  assign c_sub624 = (a623 & b_inv623) | (a623 & c623) | (b_inv623 & c623);
  wire s624, sub624, and624, or624;
  wire b_inv624;
  assign b_inv624 = ~b624;
  assign s624  = a624 ^ b624 ^ c624;
  assign sub624 = a624 ^ b_inv624 ^ c624;
  assign and624 = a624 & b624;
  assign or624  = a624 | b624;
  assign c625 = (a624 & b624) | (a624 & c624) | (b624 & c624);
  wire c_sub625;
  assign c_sub625 = (a624 & b_inv624) | (a624 & c624) | (b_inv624 & c624);
  wire s625, sub625, and625, or625;
  wire b_inv625;
  assign b_inv625 = ~b625;
  assign s625  = a625 ^ b625 ^ c625;
  assign sub625 = a625 ^ b_inv625 ^ c625;
  assign and625 = a625 & b625;
  assign or625  = a625 | b625;
  assign c626 = (a625 & b625) | (a625 & c625) | (b625 & c625);
  wire c_sub626;
  assign c_sub626 = (a625 & b_inv625) | (a625 & c625) | (b_inv625 & c625);
  wire s626, sub626, and626, or626;
  wire b_inv626;
  assign b_inv626 = ~b626;
  assign s626  = a626 ^ b626 ^ c626;
  assign sub626 = a626 ^ b_inv626 ^ c626;
  assign and626 = a626 & b626;
  assign or626  = a626 | b626;
  assign c627 = (a626 & b626) | (a626 & c626) | (b626 & c626);
  wire c_sub627;
  assign c_sub627 = (a626 & b_inv626) | (a626 & c626) | (b_inv626 & c626);
  wire s627, sub627, and627, or627;
  wire b_inv627;
  assign b_inv627 = ~b627;
  assign s627  = a627 ^ b627 ^ c627;
  assign sub627 = a627 ^ b_inv627 ^ c627;
  assign and627 = a627 & b627;
  assign or627  = a627 | b627;
  assign c628 = (a627 & b627) | (a627 & c627) | (b627 & c627);
  wire c_sub628;
  assign c_sub628 = (a627 & b_inv627) | (a627 & c627) | (b_inv627 & c627);
  wire s628, sub628, and628, or628;
  wire b_inv628;
  assign b_inv628 = ~b628;
  assign s628  = a628 ^ b628 ^ c628;
  assign sub628 = a628 ^ b_inv628 ^ c628;
  assign and628 = a628 & b628;
  assign or628  = a628 | b628;
  assign c629 = (a628 & b628) | (a628 & c628) | (b628 & c628);
  wire c_sub629;
  assign c_sub629 = (a628 & b_inv628) | (a628 & c628) | (b_inv628 & c628);
  wire s629, sub629, and629, or629;
  wire b_inv629;
  assign b_inv629 = ~b629;
  assign s629  = a629 ^ b629 ^ c629;
  assign sub629 = a629 ^ b_inv629 ^ c629;
  assign and629 = a629 & b629;
  assign or629  = a629 | b629;
  assign c630 = (a629 & b629) | (a629 & c629) | (b629 & c629);
  wire c_sub630;
  assign c_sub630 = (a629 & b_inv629) | (a629 & c629) | (b_inv629 & c629);
  wire s630, sub630, and630, or630;
  wire b_inv630;
  assign b_inv630 = ~b630;
  assign s630  = a630 ^ b630 ^ c630;
  assign sub630 = a630 ^ b_inv630 ^ c630;
  assign and630 = a630 & b630;
  assign or630  = a630 | b630;
  assign c631 = (a630 & b630) | (a630 & c630) | (b630 & c630);
  wire c_sub631;
  assign c_sub631 = (a630 & b_inv630) | (a630 & c630) | (b_inv630 & c630);
  wire s631, sub631, and631, or631;
  wire b_inv631;
  assign b_inv631 = ~b631;
  assign s631  = a631 ^ b631 ^ c631;
  assign sub631 = a631 ^ b_inv631 ^ c631;
  assign and631 = a631 & b631;
  assign or631  = a631 | b631;
  assign c632 = (a631 & b631) | (a631 & c631) | (b631 & c631);
  wire c_sub632;
  assign c_sub632 = (a631 & b_inv631) | (a631 & c631) | (b_inv631 & c631);
  wire s632, sub632, and632, or632;
  wire b_inv632;
  assign b_inv632 = ~b632;
  assign s632  = a632 ^ b632 ^ c632;
  assign sub632 = a632 ^ b_inv632 ^ c632;
  assign and632 = a632 & b632;
  assign or632  = a632 | b632;
  assign c633 = (a632 & b632) | (a632 & c632) | (b632 & c632);
  wire c_sub633;
  assign c_sub633 = (a632 & b_inv632) | (a632 & c632) | (b_inv632 & c632);
  wire s633, sub633, and633, or633;
  wire b_inv633;
  assign b_inv633 = ~b633;
  assign s633  = a633 ^ b633 ^ c633;
  assign sub633 = a633 ^ b_inv633 ^ c633;
  assign and633 = a633 & b633;
  assign or633  = a633 | b633;
  assign c634 = (a633 & b633) | (a633 & c633) | (b633 & c633);
  wire c_sub634;
  assign c_sub634 = (a633 & b_inv633) | (a633 & c633) | (b_inv633 & c633);
  wire s634, sub634, and634, or634;
  wire b_inv634;
  assign b_inv634 = ~b634;
  assign s634  = a634 ^ b634 ^ c634;
  assign sub634 = a634 ^ b_inv634 ^ c634;
  assign and634 = a634 & b634;
  assign or634  = a634 | b634;
  assign c635 = (a634 & b634) | (a634 & c634) | (b634 & c634);
  wire c_sub635;
  assign c_sub635 = (a634 & b_inv634) | (a634 & c634) | (b_inv634 & c634);
  wire s635, sub635, and635, or635;
  wire b_inv635;
  assign b_inv635 = ~b635;
  assign s635  = a635 ^ b635 ^ c635;
  assign sub635 = a635 ^ b_inv635 ^ c635;
  assign and635 = a635 & b635;
  assign or635  = a635 | b635;
  assign c636 = (a635 & b635) | (a635 & c635) | (b635 & c635);
  wire c_sub636;
  assign c_sub636 = (a635 & b_inv635) | (a635 & c635) | (b_inv635 & c635);
  wire s636, sub636, and636, or636;
  wire b_inv636;
  assign b_inv636 = ~b636;
  assign s636  = a636 ^ b636 ^ c636;
  assign sub636 = a636 ^ b_inv636 ^ c636;
  assign and636 = a636 & b636;
  assign or636  = a636 | b636;
  assign c637 = (a636 & b636) | (a636 & c636) | (b636 & c636);
  wire c_sub637;
  assign c_sub637 = (a636 & b_inv636) | (a636 & c636) | (b_inv636 & c636);
  wire s637, sub637, and637, or637;
  wire b_inv637;
  assign b_inv637 = ~b637;
  assign s637  = a637 ^ b637 ^ c637;
  assign sub637 = a637 ^ b_inv637 ^ c637;
  assign and637 = a637 & b637;
  assign or637  = a637 | b637;
  assign c638 = (a637 & b637) | (a637 & c637) | (b637 & c637);
  wire c_sub638;
  assign c_sub638 = (a637 & b_inv637) | (a637 & c637) | (b_inv637 & c637);
  wire s638, sub638, and638, or638;
  wire b_inv638;
  assign b_inv638 = ~b638;
  assign s638  = a638 ^ b638 ^ c638;
  assign sub638 = a638 ^ b_inv638 ^ c638;
  assign and638 = a638 & b638;
  assign or638  = a638 | b638;
  assign c639 = (a638 & b638) | (a638 & c638) | (b638 & c638);
  wire c_sub639;
  assign c_sub639 = (a638 & b_inv638) | (a638 & c638) | (b_inv638 & c638);
  wire s639, sub639, and639, or639;
  wire b_inv639;
  assign b_inv639 = ~b639;
  assign s639  = a639 ^ b639 ^ c639;
  assign sub639 = a639 ^ b_inv639 ^ c639;
  assign and639 = a639 & b639;
  assign or639  = a639 | b639;
  assign c640 = (a639 & b639) | (a639 & c639) | (b639 & c639);
  wire c_sub640;
  assign c_sub640 = (a639 & b_inv639) | (a639 & c639) | (b_inv639 & c639);
  wire s640, sub640, and640, or640;
  wire b_inv640;
  assign b_inv640 = ~b640;
  assign s640  = a640 ^ b640 ^ c640;
  assign sub640 = a640 ^ b_inv640 ^ c640;
  assign and640 = a640 & b640;
  assign or640  = a640 | b640;
  assign c641 = (a640 & b640) | (a640 & c640) | (b640 & c640);
  wire c_sub641;
  assign c_sub641 = (a640 & b_inv640) | (a640 & c640) | (b_inv640 & c640);
  wire s641, sub641, and641, or641;
  wire b_inv641;
  assign b_inv641 = ~b641;
  assign s641  = a641 ^ b641 ^ c641;
  assign sub641 = a641 ^ b_inv641 ^ c641;
  assign and641 = a641 & b641;
  assign or641  = a641 | b641;
  assign c642 = (a641 & b641) | (a641 & c641) | (b641 & c641);
  wire c_sub642;
  assign c_sub642 = (a641 & b_inv641) | (a641 & c641) | (b_inv641 & c641);
  wire s642, sub642, and642, or642;
  wire b_inv642;
  assign b_inv642 = ~b642;
  assign s642  = a642 ^ b642 ^ c642;
  assign sub642 = a642 ^ b_inv642 ^ c642;
  assign and642 = a642 & b642;
  assign or642  = a642 | b642;
  assign c643 = (a642 & b642) | (a642 & c642) | (b642 & c642);
  wire c_sub643;
  assign c_sub643 = (a642 & b_inv642) | (a642 & c642) | (b_inv642 & c642);
  wire s643, sub643, and643, or643;
  wire b_inv643;
  assign b_inv643 = ~b643;
  assign s643  = a643 ^ b643 ^ c643;
  assign sub643 = a643 ^ b_inv643 ^ c643;
  assign and643 = a643 & b643;
  assign or643  = a643 | b643;
  assign c644 = (a643 & b643) | (a643 & c643) | (b643 & c643);
  wire c_sub644;
  assign c_sub644 = (a643 & b_inv643) | (a643 & c643) | (b_inv643 & c643);
  wire s644, sub644, and644, or644;
  wire b_inv644;
  assign b_inv644 = ~b644;
  assign s644  = a644 ^ b644 ^ c644;
  assign sub644 = a644 ^ b_inv644 ^ c644;
  assign and644 = a644 & b644;
  assign or644  = a644 | b644;
  assign c645 = (a644 & b644) | (a644 & c644) | (b644 & c644);
  wire c_sub645;
  assign c_sub645 = (a644 & b_inv644) | (a644 & c644) | (b_inv644 & c644);
  wire s645, sub645, and645, or645;
  wire b_inv645;
  assign b_inv645 = ~b645;
  assign s645  = a645 ^ b645 ^ c645;
  assign sub645 = a645 ^ b_inv645 ^ c645;
  assign and645 = a645 & b645;
  assign or645  = a645 | b645;
  assign c646 = (a645 & b645) | (a645 & c645) | (b645 & c645);
  wire c_sub646;
  assign c_sub646 = (a645 & b_inv645) | (a645 & c645) | (b_inv645 & c645);
  wire s646, sub646, and646, or646;
  wire b_inv646;
  assign b_inv646 = ~b646;
  assign s646  = a646 ^ b646 ^ c646;
  assign sub646 = a646 ^ b_inv646 ^ c646;
  assign and646 = a646 & b646;
  assign or646  = a646 | b646;
  assign c647 = (a646 & b646) | (a646 & c646) | (b646 & c646);
  wire c_sub647;
  assign c_sub647 = (a646 & b_inv646) | (a646 & c646) | (b_inv646 & c646);
  wire s647, sub647, and647, or647;
  wire b_inv647;
  assign b_inv647 = ~b647;
  assign s647  = a647 ^ b647 ^ c647;
  assign sub647 = a647 ^ b_inv647 ^ c647;
  assign and647 = a647 & b647;
  assign or647  = a647 | b647;
  assign c648 = (a647 & b647) | (a647 & c647) | (b647 & c647);
  wire c_sub648;
  assign c_sub648 = (a647 & b_inv647) | (a647 & c647) | (b_inv647 & c647);
  wire s648, sub648, and648, or648;
  wire b_inv648;
  assign b_inv648 = ~b648;
  assign s648  = a648 ^ b648 ^ c648;
  assign sub648 = a648 ^ b_inv648 ^ c648;
  assign and648 = a648 & b648;
  assign or648  = a648 | b648;
  assign c649 = (a648 & b648) | (a648 & c648) | (b648 & c648);
  wire c_sub649;
  assign c_sub649 = (a648 & b_inv648) | (a648 & c648) | (b_inv648 & c648);
  wire s649, sub649, and649, or649;
  wire b_inv649;
  assign b_inv649 = ~b649;
  assign s649  = a649 ^ b649 ^ c649;
  assign sub649 = a649 ^ b_inv649 ^ c649;
  assign and649 = a649 & b649;
  assign or649  = a649 | b649;
  assign c650 = (a649 & b649) | (a649 & c649) | (b649 & c649);
  wire c_sub650;
  assign c_sub650 = (a649 & b_inv649) | (a649 & c649) | (b_inv649 & c649);
  wire s650, sub650, and650, or650;
  wire b_inv650;
  assign b_inv650 = ~b650;
  assign s650  = a650 ^ b650 ^ c650;
  assign sub650 = a650 ^ b_inv650 ^ c650;
  assign and650 = a650 & b650;
  assign or650  = a650 | b650;
  assign c651 = (a650 & b650) | (a650 & c650) | (b650 & c650);
  wire c_sub651;
  assign c_sub651 = (a650 & b_inv650) | (a650 & c650) | (b_inv650 & c650);
  wire s651, sub651, and651, or651;
  wire b_inv651;
  assign b_inv651 = ~b651;
  assign s651  = a651 ^ b651 ^ c651;
  assign sub651 = a651 ^ b_inv651 ^ c651;
  assign and651 = a651 & b651;
  assign or651  = a651 | b651;
  assign c652 = (a651 & b651) | (a651 & c651) | (b651 & c651);
  wire c_sub652;
  assign c_sub652 = (a651 & b_inv651) | (a651 & c651) | (b_inv651 & c651);
  wire s652, sub652, and652, or652;
  wire b_inv652;
  assign b_inv652 = ~b652;
  assign s652  = a652 ^ b652 ^ c652;
  assign sub652 = a652 ^ b_inv652 ^ c652;
  assign and652 = a652 & b652;
  assign or652  = a652 | b652;
  assign c653 = (a652 & b652) | (a652 & c652) | (b652 & c652);
  wire c_sub653;
  assign c_sub653 = (a652 & b_inv652) | (a652 & c652) | (b_inv652 & c652);
  wire s653, sub653, and653, or653;
  wire b_inv653;
  assign b_inv653 = ~b653;
  assign s653  = a653 ^ b653 ^ c653;
  assign sub653 = a653 ^ b_inv653 ^ c653;
  assign and653 = a653 & b653;
  assign or653  = a653 | b653;
  assign c654 = (a653 & b653) | (a653 & c653) | (b653 & c653);
  wire c_sub654;
  assign c_sub654 = (a653 & b_inv653) | (a653 & c653) | (b_inv653 & c653);
  wire s654, sub654, and654, or654;
  wire b_inv654;
  assign b_inv654 = ~b654;
  assign s654  = a654 ^ b654 ^ c654;
  assign sub654 = a654 ^ b_inv654 ^ c654;
  assign and654 = a654 & b654;
  assign or654  = a654 | b654;
  assign c655 = (a654 & b654) | (a654 & c654) | (b654 & c654);
  wire c_sub655;
  assign c_sub655 = (a654 & b_inv654) | (a654 & c654) | (b_inv654 & c654);
  wire s655, sub655, and655, or655;
  wire b_inv655;
  assign b_inv655 = ~b655;
  assign s655  = a655 ^ b655 ^ c655;
  assign sub655 = a655 ^ b_inv655 ^ c655;
  assign and655 = a655 & b655;
  assign or655  = a655 | b655;
  assign c656 = (a655 & b655) | (a655 & c655) | (b655 & c655);
  wire c_sub656;
  assign c_sub656 = (a655 & b_inv655) | (a655 & c655) | (b_inv655 & c655);
  wire s656, sub656, and656, or656;
  wire b_inv656;
  assign b_inv656 = ~b656;
  assign s656  = a656 ^ b656 ^ c656;
  assign sub656 = a656 ^ b_inv656 ^ c656;
  assign and656 = a656 & b656;
  assign or656  = a656 | b656;
  assign c657 = (a656 & b656) | (a656 & c656) | (b656 & c656);
  wire c_sub657;
  assign c_sub657 = (a656 & b_inv656) | (a656 & c656) | (b_inv656 & c656);
  wire s657, sub657, and657, or657;
  wire b_inv657;
  assign b_inv657 = ~b657;
  assign s657  = a657 ^ b657 ^ c657;
  assign sub657 = a657 ^ b_inv657 ^ c657;
  assign and657 = a657 & b657;
  assign or657  = a657 | b657;
  assign c658 = (a657 & b657) | (a657 & c657) | (b657 & c657);
  wire c_sub658;
  assign c_sub658 = (a657 & b_inv657) | (a657 & c657) | (b_inv657 & c657);
  wire s658, sub658, and658, or658;
  wire b_inv658;
  assign b_inv658 = ~b658;
  assign s658  = a658 ^ b658 ^ c658;
  assign sub658 = a658 ^ b_inv658 ^ c658;
  assign and658 = a658 & b658;
  assign or658  = a658 | b658;
  assign c659 = (a658 & b658) | (a658 & c658) | (b658 & c658);
  wire c_sub659;
  assign c_sub659 = (a658 & b_inv658) | (a658 & c658) | (b_inv658 & c658);
  wire s659, sub659, and659, or659;
  wire b_inv659;
  assign b_inv659 = ~b659;
  assign s659  = a659 ^ b659 ^ c659;
  assign sub659 = a659 ^ b_inv659 ^ c659;
  assign and659 = a659 & b659;
  assign or659  = a659 | b659;
  assign c660 = (a659 & b659) | (a659 & c659) | (b659 & c659);
  wire c_sub660;
  assign c_sub660 = (a659 & b_inv659) | (a659 & c659) | (b_inv659 & c659);
  wire s660, sub660, and660, or660;
  wire b_inv660;
  assign b_inv660 = ~b660;
  assign s660  = a660 ^ b660 ^ c660;
  assign sub660 = a660 ^ b_inv660 ^ c660;
  assign and660 = a660 & b660;
  assign or660  = a660 | b660;
  assign c661 = (a660 & b660) | (a660 & c660) | (b660 & c660);
  wire c_sub661;
  assign c_sub661 = (a660 & b_inv660) | (a660 & c660) | (b_inv660 & c660);
  wire s661, sub661, and661, or661;
  wire b_inv661;
  assign b_inv661 = ~b661;
  assign s661  = a661 ^ b661 ^ c661;
  assign sub661 = a661 ^ b_inv661 ^ c661;
  assign and661 = a661 & b661;
  assign or661  = a661 | b661;
  assign c662 = (a661 & b661) | (a661 & c661) | (b661 & c661);
  wire c_sub662;
  assign c_sub662 = (a661 & b_inv661) | (a661 & c661) | (b_inv661 & c661);
  wire s662, sub662, and662, or662;
  wire b_inv662;
  assign b_inv662 = ~b662;
  assign s662  = a662 ^ b662 ^ c662;
  assign sub662 = a662 ^ b_inv662 ^ c662;
  assign and662 = a662 & b662;
  assign or662  = a662 | b662;
  assign c663 = (a662 & b662) | (a662 & c662) | (b662 & c662);
  wire c_sub663;
  assign c_sub663 = (a662 & b_inv662) | (a662 & c662) | (b_inv662 & c662);
  wire s663, sub663, and663, or663;
  wire b_inv663;
  assign b_inv663 = ~b663;
  assign s663  = a663 ^ b663 ^ c663;
  assign sub663 = a663 ^ b_inv663 ^ c663;
  assign and663 = a663 & b663;
  assign or663  = a663 | b663;
  assign c664 = (a663 & b663) | (a663 & c663) | (b663 & c663);
  wire c_sub664;
  assign c_sub664 = (a663 & b_inv663) | (a663 & c663) | (b_inv663 & c663);
  wire s664, sub664, and664, or664;
  wire b_inv664;
  assign b_inv664 = ~b664;
  assign s664  = a664 ^ b664 ^ c664;
  assign sub664 = a664 ^ b_inv664 ^ c664;
  assign and664 = a664 & b664;
  assign or664  = a664 | b664;
  assign c665 = (a664 & b664) | (a664 & c664) | (b664 & c664);
  wire c_sub665;
  assign c_sub665 = (a664 & b_inv664) | (a664 & c664) | (b_inv664 & c664);
  wire s665, sub665, and665, or665;
  wire b_inv665;
  assign b_inv665 = ~b665;
  assign s665  = a665 ^ b665 ^ c665;
  assign sub665 = a665 ^ b_inv665 ^ c665;
  assign and665 = a665 & b665;
  assign or665  = a665 | b665;
  assign c666 = (a665 & b665) | (a665 & c665) | (b665 & c665);
  wire c_sub666;
  assign c_sub666 = (a665 & b_inv665) | (a665 & c665) | (b_inv665 & c665);
  wire s666, sub666, and666, or666;
  wire b_inv666;
  assign b_inv666 = ~b666;
  assign s666  = a666 ^ b666 ^ c666;
  assign sub666 = a666 ^ b_inv666 ^ c666;
  assign and666 = a666 & b666;
  assign or666  = a666 | b666;
  assign c667 = (a666 & b666) | (a666 & c666) | (b666 & c666);
  wire c_sub667;
  assign c_sub667 = (a666 & b_inv666) | (a666 & c666) | (b_inv666 & c666);
  wire s667, sub667, and667, or667;
  wire b_inv667;
  assign b_inv667 = ~b667;
  assign s667  = a667 ^ b667 ^ c667;
  assign sub667 = a667 ^ b_inv667 ^ c667;
  assign and667 = a667 & b667;
  assign or667  = a667 | b667;
  assign c668 = (a667 & b667) | (a667 & c667) | (b667 & c667);
  wire c_sub668;
  assign c_sub668 = (a667 & b_inv667) | (a667 & c667) | (b_inv667 & c667);
  wire s668, sub668, and668, or668;
  wire b_inv668;
  assign b_inv668 = ~b668;
  assign s668  = a668 ^ b668 ^ c668;
  assign sub668 = a668 ^ b_inv668 ^ c668;
  assign and668 = a668 & b668;
  assign or668  = a668 | b668;
  assign c669 = (a668 & b668) | (a668 & c668) | (b668 & c668);
  wire c_sub669;
  assign c_sub669 = (a668 & b_inv668) | (a668 & c668) | (b_inv668 & c668);
  wire s669, sub669, and669, or669;
  wire b_inv669;
  assign b_inv669 = ~b669;
  assign s669  = a669 ^ b669 ^ c669;
  assign sub669 = a669 ^ b_inv669 ^ c669;
  assign and669 = a669 & b669;
  assign or669  = a669 | b669;
  assign c670 = (a669 & b669) | (a669 & c669) | (b669 & c669);
  wire c_sub670;
  assign c_sub670 = (a669 & b_inv669) | (a669 & c669) | (b_inv669 & c669);
  wire s670, sub670, and670, or670;
  wire b_inv670;
  assign b_inv670 = ~b670;
  assign s670  = a670 ^ b670 ^ c670;
  assign sub670 = a670 ^ b_inv670 ^ c670;
  assign and670 = a670 & b670;
  assign or670  = a670 | b670;
  assign c671 = (a670 & b670) | (a670 & c670) | (b670 & c670);
  wire c_sub671;
  assign c_sub671 = (a670 & b_inv670) | (a670 & c670) | (b_inv670 & c670);
  wire s671, sub671, and671, or671;
  wire b_inv671;
  assign b_inv671 = ~b671;
  assign s671  = a671 ^ b671 ^ c671;
  assign sub671 = a671 ^ b_inv671 ^ c671;
  assign and671 = a671 & b671;
  assign or671  = a671 | b671;
  assign c672 = (a671 & b671) | (a671 & c671) | (b671 & c671);
  wire c_sub672;
  assign c_sub672 = (a671 & b_inv671) | (a671 & c671) | (b_inv671 & c671);
  wire s672, sub672, and672, or672;
  wire b_inv672;
  assign b_inv672 = ~b672;
  assign s672  = a672 ^ b672 ^ c672;
  assign sub672 = a672 ^ b_inv672 ^ c672;
  assign and672 = a672 & b672;
  assign or672  = a672 | b672;
  assign c673 = (a672 & b672) | (a672 & c672) | (b672 & c672);
  wire c_sub673;
  assign c_sub673 = (a672 & b_inv672) | (a672 & c672) | (b_inv672 & c672);
  wire s673, sub673, and673, or673;
  wire b_inv673;
  assign b_inv673 = ~b673;
  assign s673  = a673 ^ b673 ^ c673;
  assign sub673 = a673 ^ b_inv673 ^ c673;
  assign and673 = a673 & b673;
  assign or673  = a673 | b673;
  assign c674 = (a673 & b673) | (a673 & c673) | (b673 & c673);
  wire c_sub674;
  assign c_sub674 = (a673 & b_inv673) | (a673 & c673) | (b_inv673 & c673);
  wire s674, sub674, and674, or674;
  wire b_inv674;
  assign b_inv674 = ~b674;
  assign s674  = a674 ^ b674 ^ c674;
  assign sub674 = a674 ^ b_inv674 ^ c674;
  assign and674 = a674 & b674;
  assign or674  = a674 | b674;
  assign c675 = (a674 & b674) | (a674 & c674) | (b674 & c674);
  wire c_sub675;
  assign c_sub675 = (a674 & b_inv674) | (a674 & c674) | (b_inv674 & c674);
  wire s675, sub675, and675, or675;
  wire b_inv675;
  assign b_inv675 = ~b675;
  assign s675  = a675 ^ b675 ^ c675;
  assign sub675 = a675 ^ b_inv675 ^ c675;
  assign and675 = a675 & b675;
  assign or675  = a675 | b675;
  assign c676 = (a675 & b675) | (a675 & c675) | (b675 & c675);
  wire c_sub676;
  assign c_sub676 = (a675 & b_inv675) | (a675 & c675) | (b_inv675 & c675);
  wire s676, sub676, and676, or676;
  wire b_inv676;
  assign b_inv676 = ~b676;
  assign s676  = a676 ^ b676 ^ c676;
  assign sub676 = a676 ^ b_inv676 ^ c676;
  assign and676 = a676 & b676;
  assign or676  = a676 | b676;
  assign c677 = (a676 & b676) | (a676 & c676) | (b676 & c676);
  wire c_sub677;
  assign c_sub677 = (a676 & b_inv676) | (a676 & c676) | (b_inv676 & c676);
  wire s677, sub677, and677, or677;
  wire b_inv677;
  assign b_inv677 = ~b677;
  assign s677  = a677 ^ b677 ^ c677;
  assign sub677 = a677 ^ b_inv677 ^ c677;
  assign and677 = a677 & b677;
  assign or677  = a677 | b677;
  assign c678 = (a677 & b677) | (a677 & c677) | (b677 & c677);
  wire c_sub678;
  assign c_sub678 = (a677 & b_inv677) | (a677 & c677) | (b_inv677 & c677);
  wire s678, sub678, and678, or678;
  wire b_inv678;
  assign b_inv678 = ~b678;
  assign s678  = a678 ^ b678 ^ c678;
  assign sub678 = a678 ^ b_inv678 ^ c678;
  assign and678 = a678 & b678;
  assign or678  = a678 | b678;
  assign c679 = (a678 & b678) | (a678 & c678) | (b678 & c678);
  wire c_sub679;
  assign c_sub679 = (a678 & b_inv678) | (a678 & c678) | (b_inv678 & c678);
  wire s679, sub679, and679, or679;
  wire b_inv679;
  assign b_inv679 = ~b679;
  assign s679  = a679 ^ b679 ^ c679;
  assign sub679 = a679 ^ b_inv679 ^ c679;
  assign and679 = a679 & b679;
  assign or679  = a679 | b679;
  assign c680 = (a679 & b679) | (a679 & c679) | (b679 & c679);
  wire c_sub680;
  assign c_sub680 = (a679 & b_inv679) | (a679 & c679) | (b_inv679 & c679);
  wire s680, sub680, and680, or680;
  wire b_inv680;
  assign b_inv680 = ~b680;
  assign s680  = a680 ^ b680 ^ c680;
  assign sub680 = a680 ^ b_inv680 ^ c680;
  assign and680 = a680 & b680;
  assign or680  = a680 | b680;
  assign c681 = (a680 & b680) | (a680 & c680) | (b680 & c680);
  wire c_sub681;
  assign c_sub681 = (a680 & b_inv680) | (a680 & c680) | (b_inv680 & c680);
  wire s681, sub681, and681, or681;
  wire b_inv681;
  assign b_inv681 = ~b681;
  assign s681  = a681 ^ b681 ^ c681;
  assign sub681 = a681 ^ b_inv681 ^ c681;
  assign and681 = a681 & b681;
  assign or681  = a681 | b681;
  assign c682 = (a681 & b681) | (a681 & c681) | (b681 & c681);
  wire c_sub682;
  assign c_sub682 = (a681 & b_inv681) | (a681 & c681) | (b_inv681 & c681);
  wire s682, sub682, and682, or682;
  wire b_inv682;
  assign b_inv682 = ~b682;
  assign s682  = a682 ^ b682 ^ c682;
  assign sub682 = a682 ^ b_inv682 ^ c682;
  assign and682 = a682 & b682;
  assign or682  = a682 | b682;
  assign c683 = (a682 & b682) | (a682 & c682) | (b682 & c682);
  wire c_sub683;
  assign c_sub683 = (a682 & b_inv682) | (a682 & c682) | (b_inv682 & c682);
  wire s683, sub683, and683, or683;
  wire b_inv683;
  assign b_inv683 = ~b683;
  assign s683  = a683 ^ b683 ^ c683;
  assign sub683 = a683 ^ b_inv683 ^ c683;
  assign and683 = a683 & b683;
  assign or683  = a683 | b683;
  assign c684 = (a683 & b683) | (a683 & c683) | (b683 & c683);
  wire c_sub684;
  assign c_sub684 = (a683 & b_inv683) | (a683 & c683) | (b_inv683 & c683);
  wire s684, sub684, and684, or684;
  wire b_inv684;
  assign b_inv684 = ~b684;
  assign s684  = a684 ^ b684 ^ c684;
  assign sub684 = a684 ^ b_inv684 ^ c684;
  assign and684 = a684 & b684;
  assign or684  = a684 | b684;
  assign c685 = (a684 & b684) | (a684 & c684) | (b684 & c684);
  wire c_sub685;
  assign c_sub685 = (a684 & b_inv684) | (a684 & c684) | (b_inv684 & c684);
  wire s685, sub685, and685, or685;
  wire b_inv685;
  assign b_inv685 = ~b685;
  assign s685  = a685 ^ b685 ^ c685;
  assign sub685 = a685 ^ b_inv685 ^ c685;
  assign and685 = a685 & b685;
  assign or685  = a685 | b685;
  assign c686 = (a685 & b685) | (a685 & c685) | (b685 & c685);
  wire c_sub686;
  assign c_sub686 = (a685 & b_inv685) | (a685 & c685) | (b_inv685 & c685);
  wire s686, sub686, and686, or686;
  wire b_inv686;
  assign b_inv686 = ~b686;
  assign s686  = a686 ^ b686 ^ c686;
  assign sub686 = a686 ^ b_inv686 ^ c686;
  assign and686 = a686 & b686;
  assign or686  = a686 | b686;
  assign c687 = (a686 & b686) | (a686 & c686) | (b686 & c686);
  wire c_sub687;
  assign c_sub687 = (a686 & b_inv686) | (a686 & c686) | (b_inv686 & c686);
  wire s687, sub687, and687, or687;
  wire b_inv687;
  assign b_inv687 = ~b687;
  assign s687  = a687 ^ b687 ^ c687;
  assign sub687 = a687 ^ b_inv687 ^ c687;
  assign and687 = a687 & b687;
  assign or687  = a687 | b687;
  assign c688 = (a687 & b687) | (a687 & c687) | (b687 & c687);
  wire c_sub688;
  assign c_sub688 = (a687 & b_inv687) | (a687 & c687) | (b_inv687 & c687);
  wire s688, sub688, and688, or688;
  wire b_inv688;
  assign b_inv688 = ~b688;
  assign s688  = a688 ^ b688 ^ c688;
  assign sub688 = a688 ^ b_inv688 ^ c688;
  assign and688 = a688 & b688;
  assign or688  = a688 | b688;
  assign c689 = (a688 & b688) | (a688 & c688) | (b688 & c688);
  wire c_sub689;
  assign c_sub689 = (a688 & b_inv688) | (a688 & c688) | (b_inv688 & c688);
  wire s689, sub689, and689, or689;
  wire b_inv689;
  assign b_inv689 = ~b689;
  assign s689  = a689 ^ b689 ^ c689;
  assign sub689 = a689 ^ b_inv689 ^ c689;
  assign and689 = a689 & b689;
  assign or689  = a689 | b689;
  assign c690 = (a689 & b689) | (a689 & c689) | (b689 & c689);
  wire c_sub690;
  assign c_sub690 = (a689 & b_inv689) | (a689 & c689) | (b_inv689 & c689);
  wire s690, sub690, and690, or690;
  wire b_inv690;
  assign b_inv690 = ~b690;
  assign s690  = a690 ^ b690 ^ c690;
  assign sub690 = a690 ^ b_inv690 ^ c690;
  assign and690 = a690 & b690;
  assign or690  = a690 | b690;
  assign c691 = (a690 & b690) | (a690 & c690) | (b690 & c690);
  wire c_sub691;
  assign c_sub691 = (a690 & b_inv690) | (a690 & c690) | (b_inv690 & c690);
  wire s691, sub691, and691, or691;
  wire b_inv691;
  assign b_inv691 = ~b691;
  assign s691  = a691 ^ b691 ^ c691;
  assign sub691 = a691 ^ b_inv691 ^ c691;
  assign and691 = a691 & b691;
  assign or691  = a691 | b691;
  assign c692 = (a691 & b691) | (a691 & c691) | (b691 & c691);
  wire c_sub692;
  assign c_sub692 = (a691 & b_inv691) | (a691 & c691) | (b_inv691 & c691);
  wire s692, sub692, and692, or692;
  wire b_inv692;
  assign b_inv692 = ~b692;
  assign s692  = a692 ^ b692 ^ c692;
  assign sub692 = a692 ^ b_inv692 ^ c692;
  assign and692 = a692 & b692;
  assign or692  = a692 | b692;
  assign c693 = (a692 & b692) | (a692 & c692) | (b692 & c692);
  wire c_sub693;
  assign c_sub693 = (a692 & b_inv692) | (a692 & c692) | (b_inv692 & c692);
  wire s693, sub693, and693, or693;
  wire b_inv693;
  assign b_inv693 = ~b693;
  assign s693  = a693 ^ b693 ^ c693;
  assign sub693 = a693 ^ b_inv693 ^ c693;
  assign and693 = a693 & b693;
  assign or693  = a693 | b693;
  assign c694 = (a693 & b693) | (a693 & c693) | (b693 & c693);
  wire c_sub694;
  assign c_sub694 = (a693 & b_inv693) | (a693 & c693) | (b_inv693 & c693);
  wire s694, sub694, and694, or694;
  wire b_inv694;
  assign b_inv694 = ~b694;
  assign s694  = a694 ^ b694 ^ c694;
  assign sub694 = a694 ^ b_inv694 ^ c694;
  assign and694 = a694 & b694;
  assign or694  = a694 | b694;
  assign c695 = (a694 & b694) | (a694 & c694) | (b694 & c694);
  wire c_sub695;
  assign c_sub695 = (a694 & b_inv694) | (a694 & c694) | (b_inv694 & c694);
  wire s695, sub695, and695, or695;
  wire b_inv695;
  assign b_inv695 = ~b695;
  assign s695  = a695 ^ b695 ^ c695;
  assign sub695 = a695 ^ b_inv695 ^ c695;
  assign and695 = a695 & b695;
  assign or695  = a695 | b695;
  assign c696 = (a695 & b695) | (a695 & c695) | (b695 & c695);
  wire c_sub696;
  assign c_sub696 = (a695 & b_inv695) | (a695 & c695) | (b_inv695 & c695);
  wire s696, sub696, and696, or696;
  wire b_inv696;
  assign b_inv696 = ~b696;
  assign s696  = a696 ^ b696 ^ c696;
  assign sub696 = a696 ^ b_inv696 ^ c696;
  assign and696 = a696 & b696;
  assign or696  = a696 | b696;
  assign c697 = (a696 & b696) | (a696 & c696) | (b696 & c696);
  wire c_sub697;
  assign c_sub697 = (a696 & b_inv696) | (a696 & c696) | (b_inv696 & c696);
  wire s697, sub697, and697, or697;
  wire b_inv697;
  assign b_inv697 = ~b697;
  assign s697  = a697 ^ b697 ^ c697;
  assign sub697 = a697 ^ b_inv697 ^ c697;
  assign and697 = a697 & b697;
  assign or697  = a697 | b697;
  assign c698 = (a697 & b697) | (a697 & c697) | (b697 & c697);
  wire c_sub698;
  assign c_sub698 = (a697 & b_inv697) | (a697 & c697) | (b_inv697 & c697);
  wire s698, sub698, and698, or698;
  wire b_inv698;
  assign b_inv698 = ~b698;
  assign s698  = a698 ^ b698 ^ c698;
  assign sub698 = a698 ^ b_inv698 ^ c698;
  assign and698 = a698 & b698;
  assign or698  = a698 | b698;
  assign c699 = (a698 & b698) | (a698 & c698) | (b698 & c698);
  wire c_sub699;
  assign c_sub699 = (a698 & b_inv698) | (a698 & c698) | (b_inv698 & c698);
  wire s699, sub699, and699, or699;
  wire b_inv699;
  assign b_inv699 = ~b699;
  assign s699  = a699 ^ b699 ^ c699;
  assign sub699 = a699 ^ b_inv699 ^ c699;
  assign and699 = a699 & b699;
  assign or699  = a699 | b699;
  assign c700 = (a699 & b699) | (a699 & c699) | (b699 & c699);
  wire c_sub700;
  assign c_sub700 = (a699 & b_inv699) | (a699 & c699) | (b_inv699 & c699);
  wire s700, sub700, and700, or700;
  wire b_inv700;
  assign b_inv700 = ~b700;
  assign s700  = a700 ^ b700 ^ c700;
  assign sub700 = a700 ^ b_inv700 ^ c700;
  assign and700 = a700 & b700;
  assign or700  = a700 | b700;
  assign c701 = (a700 & b700) | (a700 & c700) | (b700 & c700);
  wire c_sub701;
  assign c_sub701 = (a700 & b_inv700) | (a700 & c700) | (b_inv700 & c700);
  wire s701, sub701, and701, or701;
  wire b_inv701;
  assign b_inv701 = ~b701;
  assign s701  = a701 ^ b701 ^ c701;
  assign sub701 = a701 ^ b_inv701 ^ c701;
  assign and701 = a701 & b701;
  assign or701  = a701 | b701;
  assign c702 = (a701 & b701) | (a701 & c701) | (b701 & c701);
  wire c_sub702;
  assign c_sub702 = (a701 & b_inv701) | (a701 & c701) | (b_inv701 & c701);
  wire s702, sub702, and702, or702;
  wire b_inv702;
  assign b_inv702 = ~b702;
  assign s702  = a702 ^ b702 ^ c702;
  assign sub702 = a702 ^ b_inv702 ^ c702;
  assign and702 = a702 & b702;
  assign or702  = a702 | b702;
  assign c703 = (a702 & b702) | (a702 & c702) | (b702 & c702);
  wire c_sub703;
  assign c_sub703 = (a702 & b_inv702) | (a702 & c702) | (b_inv702 & c702);
  wire s703, sub703, and703, or703;
  wire b_inv703;
  assign b_inv703 = ~b703;
  assign s703  = a703 ^ b703 ^ c703;
  assign sub703 = a703 ^ b_inv703 ^ c703;
  assign and703 = a703 & b703;
  assign or703  = a703 | b703;
  assign c704 = (a703 & b703) | (a703 & c703) | (b703 & c703);
  wire c_sub704;
  assign c_sub704 = (a703 & b_inv703) | (a703 & c703) | (b_inv703 & c703);
  wire s704, sub704, and704, or704;
  wire b_inv704;
  assign b_inv704 = ~b704;
  assign s704  = a704 ^ b704 ^ c704;
  assign sub704 = a704 ^ b_inv704 ^ c704;
  assign and704 = a704 & b704;
  assign or704  = a704 | b704;
  assign c705 = (a704 & b704) | (a704 & c704) | (b704 & c704);
  wire c_sub705;
  assign c_sub705 = (a704 & b_inv704) | (a704 & c704) | (b_inv704 & c704);
  wire s705, sub705, and705, or705;
  wire b_inv705;
  assign b_inv705 = ~b705;
  assign s705  = a705 ^ b705 ^ c705;
  assign sub705 = a705 ^ b_inv705 ^ c705;
  assign and705 = a705 & b705;
  assign or705  = a705 | b705;
  assign c706 = (a705 & b705) | (a705 & c705) | (b705 & c705);
  wire c_sub706;
  assign c_sub706 = (a705 & b_inv705) | (a705 & c705) | (b_inv705 & c705);
  wire s706, sub706, and706, or706;
  wire b_inv706;
  assign b_inv706 = ~b706;
  assign s706  = a706 ^ b706 ^ c706;
  assign sub706 = a706 ^ b_inv706 ^ c706;
  assign and706 = a706 & b706;
  assign or706  = a706 | b706;
  assign c707 = (a706 & b706) | (a706 & c706) | (b706 & c706);
  wire c_sub707;
  assign c_sub707 = (a706 & b_inv706) | (a706 & c706) | (b_inv706 & c706);
  wire s707, sub707, and707, or707;
  wire b_inv707;
  assign b_inv707 = ~b707;
  assign s707  = a707 ^ b707 ^ c707;
  assign sub707 = a707 ^ b_inv707 ^ c707;
  assign and707 = a707 & b707;
  assign or707  = a707 | b707;
  assign c708 = (a707 & b707) | (a707 & c707) | (b707 & c707);
  wire c_sub708;
  assign c_sub708 = (a707 & b_inv707) | (a707 & c707) | (b_inv707 & c707);
  wire s708, sub708, and708, or708;
  wire b_inv708;
  assign b_inv708 = ~b708;
  assign s708  = a708 ^ b708 ^ c708;
  assign sub708 = a708 ^ b_inv708 ^ c708;
  assign and708 = a708 & b708;
  assign or708  = a708 | b708;
  assign c709 = (a708 & b708) | (a708 & c708) | (b708 & c708);
  wire c_sub709;
  assign c_sub709 = (a708 & b_inv708) | (a708 & c708) | (b_inv708 & c708);
  wire s709, sub709, and709, or709;
  wire b_inv709;
  assign b_inv709 = ~b709;
  assign s709  = a709 ^ b709 ^ c709;
  assign sub709 = a709 ^ b_inv709 ^ c709;
  assign and709 = a709 & b709;
  assign or709  = a709 | b709;
  assign c710 = (a709 & b709) | (a709 & c709) | (b709 & c709);
  wire c_sub710;
  assign c_sub710 = (a709 & b_inv709) | (a709 & c709) | (b_inv709 & c709);
  wire s710, sub710, and710, or710;
  wire b_inv710;
  assign b_inv710 = ~b710;
  assign s710  = a710 ^ b710 ^ c710;
  assign sub710 = a710 ^ b_inv710 ^ c710;
  assign and710 = a710 & b710;
  assign or710  = a710 | b710;
  assign c711 = (a710 & b710) | (a710 & c710) | (b710 & c710);
  wire c_sub711;
  assign c_sub711 = (a710 & b_inv710) | (a710 & c710) | (b_inv710 & c710);
  wire s711, sub711, and711, or711;
  wire b_inv711;
  assign b_inv711 = ~b711;
  assign s711  = a711 ^ b711 ^ c711;
  assign sub711 = a711 ^ b_inv711 ^ c711;
  assign and711 = a711 & b711;
  assign or711  = a711 | b711;
  assign c712 = (a711 & b711) | (a711 & c711) | (b711 & c711);
  wire c_sub712;
  assign c_sub712 = (a711 & b_inv711) | (a711 & c711) | (b_inv711 & c711);
  wire s712, sub712, and712, or712;
  wire b_inv712;
  assign b_inv712 = ~b712;
  assign s712  = a712 ^ b712 ^ c712;
  assign sub712 = a712 ^ b_inv712 ^ c712;
  assign and712 = a712 & b712;
  assign or712  = a712 | b712;
  assign c713 = (a712 & b712) | (a712 & c712) | (b712 & c712);
  wire c_sub713;
  assign c_sub713 = (a712 & b_inv712) | (a712 & c712) | (b_inv712 & c712);
  wire s713, sub713, and713, or713;
  wire b_inv713;
  assign b_inv713 = ~b713;
  assign s713  = a713 ^ b713 ^ c713;
  assign sub713 = a713 ^ b_inv713 ^ c713;
  assign and713 = a713 & b713;
  assign or713  = a713 | b713;
  assign c714 = (a713 & b713) | (a713 & c713) | (b713 & c713);
  wire c_sub714;
  assign c_sub714 = (a713 & b_inv713) | (a713 & c713) | (b_inv713 & c713);
  wire s714, sub714, and714, or714;
  wire b_inv714;
  assign b_inv714 = ~b714;
  assign s714  = a714 ^ b714 ^ c714;
  assign sub714 = a714 ^ b_inv714 ^ c714;
  assign and714 = a714 & b714;
  assign or714  = a714 | b714;
  assign c715 = (a714 & b714) | (a714 & c714) | (b714 & c714);
  wire c_sub715;
  assign c_sub715 = (a714 & b_inv714) | (a714 & c714) | (b_inv714 & c714);
  wire s715, sub715, and715, or715;
  wire b_inv715;
  assign b_inv715 = ~b715;
  assign s715  = a715 ^ b715 ^ c715;
  assign sub715 = a715 ^ b_inv715 ^ c715;
  assign and715 = a715 & b715;
  assign or715  = a715 | b715;
  assign c716 = (a715 & b715) | (a715 & c715) | (b715 & c715);
  wire c_sub716;
  assign c_sub716 = (a715 & b_inv715) | (a715 & c715) | (b_inv715 & c715);
  wire s716, sub716, and716, or716;
  wire b_inv716;
  assign b_inv716 = ~b716;
  assign s716  = a716 ^ b716 ^ c716;
  assign sub716 = a716 ^ b_inv716 ^ c716;
  assign and716 = a716 & b716;
  assign or716  = a716 | b716;
  assign c717 = (a716 & b716) | (a716 & c716) | (b716 & c716);
  wire c_sub717;
  assign c_sub717 = (a716 & b_inv716) | (a716 & c716) | (b_inv716 & c716);
  wire s717, sub717, and717, or717;
  wire b_inv717;
  assign b_inv717 = ~b717;
  assign s717  = a717 ^ b717 ^ c717;
  assign sub717 = a717 ^ b_inv717 ^ c717;
  assign and717 = a717 & b717;
  assign or717  = a717 | b717;
  assign c718 = (a717 & b717) | (a717 & c717) | (b717 & c717);
  wire c_sub718;
  assign c_sub718 = (a717 & b_inv717) | (a717 & c717) | (b_inv717 & c717);
  wire s718, sub718, and718, or718;
  wire b_inv718;
  assign b_inv718 = ~b718;
  assign s718  = a718 ^ b718 ^ c718;
  assign sub718 = a718 ^ b_inv718 ^ c718;
  assign and718 = a718 & b718;
  assign or718  = a718 | b718;
  assign c719 = (a718 & b718) | (a718 & c718) | (b718 & c718);
  wire c_sub719;
  assign c_sub719 = (a718 & b_inv718) | (a718 & c718) | (b_inv718 & c718);
  wire s719, sub719, and719, or719;
  wire b_inv719;
  assign b_inv719 = ~b719;
  assign s719  = a719 ^ b719 ^ c719;
  assign sub719 = a719 ^ b_inv719 ^ c719;
  assign and719 = a719 & b719;
  assign or719  = a719 | b719;
  assign c720 = (a719 & b719) | (a719 & c719) | (b719 & c719);
  wire c_sub720;
  assign c_sub720 = (a719 & b_inv719) | (a719 & c719) | (b_inv719 & c719);
  wire s720, sub720, and720, or720;
  wire b_inv720;
  assign b_inv720 = ~b720;
  assign s720  = a720 ^ b720 ^ c720;
  assign sub720 = a720 ^ b_inv720 ^ c720;
  assign and720 = a720 & b720;
  assign or720  = a720 | b720;
  assign c721 = (a720 & b720) | (a720 & c720) | (b720 & c720);
  wire c_sub721;
  assign c_sub721 = (a720 & b_inv720) | (a720 & c720) | (b_inv720 & c720);
  wire s721, sub721, and721, or721;
  wire b_inv721;
  assign b_inv721 = ~b721;
  assign s721  = a721 ^ b721 ^ c721;
  assign sub721 = a721 ^ b_inv721 ^ c721;
  assign and721 = a721 & b721;
  assign or721  = a721 | b721;
  assign c722 = (a721 & b721) | (a721 & c721) | (b721 & c721);
  wire c_sub722;
  assign c_sub722 = (a721 & b_inv721) | (a721 & c721) | (b_inv721 & c721);
  wire s722, sub722, and722, or722;
  wire b_inv722;
  assign b_inv722 = ~b722;
  assign s722  = a722 ^ b722 ^ c722;
  assign sub722 = a722 ^ b_inv722 ^ c722;
  assign and722 = a722 & b722;
  assign or722  = a722 | b722;
  assign c723 = (a722 & b722) | (a722 & c722) | (b722 & c722);
  wire c_sub723;
  assign c_sub723 = (a722 & b_inv722) | (a722 & c722) | (b_inv722 & c722);
  wire s723, sub723, and723, or723;
  wire b_inv723;
  assign b_inv723 = ~b723;
  assign s723  = a723 ^ b723 ^ c723;
  assign sub723 = a723 ^ b_inv723 ^ c723;
  assign and723 = a723 & b723;
  assign or723  = a723 | b723;
  assign c724 = (a723 & b723) | (a723 & c723) | (b723 & c723);
  wire c_sub724;
  assign c_sub724 = (a723 & b_inv723) | (a723 & c723) | (b_inv723 & c723);
  wire s724, sub724, and724, or724;
  wire b_inv724;
  assign b_inv724 = ~b724;
  assign s724  = a724 ^ b724 ^ c724;
  assign sub724 = a724 ^ b_inv724 ^ c724;
  assign and724 = a724 & b724;
  assign or724  = a724 | b724;
  assign c725 = (a724 & b724) | (a724 & c724) | (b724 & c724);
  wire c_sub725;
  assign c_sub725 = (a724 & b_inv724) | (a724 & c724) | (b_inv724 & c724);
  wire s725, sub725, and725, or725;
  wire b_inv725;
  assign b_inv725 = ~b725;
  assign s725  = a725 ^ b725 ^ c725;
  assign sub725 = a725 ^ b_inv725 ^ c725;
  assign and725 = a725 & b725;
  assign or725  = a725 | b725;
  assign c726 = (a725 & b725) | (a725 & c725) | (b725 & c725);
  wire c_sub726;
  assign c_sub726 = (a725 & b_inv725) | (a725 & c725) | (b_inv725 & c725);
  wire s726, sub726, and726, or726;
  wire b_inv726;
  assign b_inv726 = ~b726;
  assign s726  = a726 ^ b726 ^ c726;
  assign sub726 = a726 ^ b_inv726 ^ c726;
  assign and726 = a726 & b726;
  assign or726  = a726 | b726;
  assign c727 = (a726 & b726) | (a726 & c726) | (b726 & c726);
  wire c_sub727;
  assign c_sub727 = (a726 & b_inv726) | (a726 & c726) | (b_inv726 & c726);
  wire s727, sub727, and727, or727;
  wire b_inv727;
  assign b_inv727 = ~b727;
  assign s727  = a727 ^ b727 ^ c727;
  assign sub727 = a727 ^ b_inv727 ^ c727;
  assign and727 = a727 & b727;
  assign or727  = a727 | b727;
  assign c728 = (a727 & b727) | (a727 & c727) | (b727 & c727);
  wire c_sub728;
  assign c_sub728 = (a727 & b_inv727) | (a727 & c727) | (b_inv727 & c727);
  wire s728, sub728, and728, or728;
  wire b_inv728;
  assign b_inv728 = ~b728;
  assign s728  = a728 ^ b728 ^ c728;
  assign sub728 = a728 ^ b_inv728 ^ c728;
  assign and728 = a728 & b728;
  assign or728  = a728 | b728;
  assign c729 = (a728 & b728) | (a728 & c728) | (b728 & c728);
  wire c_sub729;
  assign c_sub729 = (a728 & b_inv728) | (a728 & c728) | (b_inv728 & c728);
  wire s729, sub729, and729, or729;
  wire b_inv729;
  assign b_inv729 = ~b729;
  assign s729  = a729 ^ b729 ^ c729;
  assign sub729 = a729 ^ b_inv729 ^ c729;
  assign and729 = a729 & b729;
  assign or729  = a729 | b729;
  assign c730 = (a729 & b729) | (a729 & c729) | (b729 & c729);
  wire c_sub730;
  assign c_sub730 = (a729 & b_inv729) | (a729 & c729) | (b_inv729 & c729);
  wire s730, sub730, and730, or730;
  wire b_inv730;
  assign b_inv730 = ~b730;
  assign s730  = a730 ^ b730 ^ c730;
  assign sub730 = a730 ^ b_inv730 ^ c730;
  assign and730 = a730 & b730;
  assign or730  = a730 | b730;
  assign c731 = (a730 & b730) | (a730 & c730) | (b730 & c730);
  wire c_sub731;
  assign c_sub731 = (a730 & b_inv730) | (a730 & c730) | (b_inv730 & c730);
  wire s731, sub731, and731, or731;
  wire b_inv731;
  assign b_inv731 = ~b731;
  assign s731  = a731 ^ b731 ^ c731;
  assign sub731 = a731 ^ b_inv731 ^ c731;
  assign and731 = a731 & b731;
  assign or731  = a731 | b731;
  assign c732 = (a731 & b731) | (a731 & c731) | (b731 & c731);
  wire c_sub732;
  assign c_sub732 = (a731 & b_inv731) | (a731 & c731) | (b_inv731 & c731);
  wire s732, sub732, and732, or732;
  wire b_inv732;
  assign b_inv732 = ~b732;
  assign s732  = a732 ^ b732 ^ c732;
  assign sub732 = a732 ^ b_inv732 ^ c732;
  assign and732 = a732 & b732;
  assign or732  = a732 | b732;
  assign c733 = (a732 & b732) | (a732 & c732) | (b732 & c732);
  wire c_sub733;
  assign c_sub733 = (a732 & b_inv732) | (a732 & c732) | (b_inv732 & c732);
  wire s733, sub733, and733, or733;
  wire b_inv733;
  assign b_inv733 = ~b733;
  assign s733  = a733 ^ b733 ^ c733;
  assign sub733 = a733 ^ b_inv733 ^ c733;
  assign and733 = a733 & b733;
  assign or733  = a733 | b733;
  assign c734 = (a733 & b733) | (a733 & c733) | (b733 & c733);
  wire c_sub734;
  assign c_sub734 = (a733 & b_inv733) | (a733 & c733) | (b_inv733 & c733);
  wire s734, sub734, and734, or734;
  wire b_inv734;
  assign b_inv734 = ~b734;
  assign s734  = a734 ^ b734 ^ c734;
  assign sub734 = a734 ^ b_inv734 ^ c734;
  assign and734 = a734 & b734;
  assign or734  = a734 | b734;
  assign c735 = (a734 & b734) | (a734 & c734) | (b734 & c734);
  wire c_sub735;
  assign c_sub735 = (a734 & b_inv734) | (a734 & c734) | (b_inv734 & c734);
  wire s735, sub735, and735, or735;
  wire b_inv735;
  assign b_inv735 = ~b735;
  assign s735  = a735 ^ b735 ^ c735;
  assign sub735 = a735 ^ b_inv735 ^ c735;
  assign and735 = a735 & b735;
  assign or735  = a735 | b735;
  assign c736 = (a735 & b735) | (a735 & c735) | (b735 & c735);
  wire c_sub736;
  assign c_sub736 = (a735 & b_inv735) | (a735 & c735) | (b_inv735 & c735);
  wire s736, sub736, and736, or736;
  wire b_inv736;
  assign b_inv736 = ~b736;
  assign s736  = a736 ^ b736 ^ c736;
  assign sub736 = a736 ^ b_inv736 ^ c736;
  assign and736 = a736 & b736;
  assign or736  = a736 | b736;
  assign c737 = (a736 & b736) | (a736 & c736) | (b736 & c736);
  wire c_sub737;
  assign c_sub737 = (a736 & b_inv736) | (a736 & c736) | (b_inv736 & c736);
  wire s737, sub737, and737, or737;
  wire b_inv737;
  assign b_inv737 = ~b737;
  assign s737  = a737 ^ b737 ^ c737;
  assign sub737 = a737 ^ b_inv737 ^ c737;
  assign and737 = a737 & b737;
  assign or737  = a737 | b737;
  assign c738 = (a737 & b737) | (a737 & c737) | (b737 & c737);
  wire c_sub738;
  assign c_sub738 = (a737 & b_inv737) | (a737 & c737) | (b_inv737 & c737);
  wire s738, sub738, and738, or738;
  wire b_inv738;
  assign b_inv738 = ~b738;
  assign s738  = a738 ^ b738 ^ c738;
  assign sub738 = a738 ^ b_inv738 ^ c738;
  assign and738 = a738 & b738;
  assign or738  = a738 | b738;
  assign c739 = (a738 & b738) | (a738 & c738) | (b738 & c738);
  wire c_sub739;
  assign c_sub739 = (a738 & b_inv738) | (a738 & c738) | (b_inv738 & c738);
  wire s739, sub739, and739, or739;
  wire b_inv739;
  assign b_inv739 = ~b739;
  assign s739  = a739 ^ b739 ^ c739;
  assign sub739 = a739 ^ b_inv739 ^ c739;
  assign and739 = a739 & b739;
  assign or739  = a739 | b739;
  assign c740 = (a739 & b739) | (a739 & c739) | (b739 & c739);
  wire c_sub740;
  assign c_sub740 = (a739 & b_inv739) | (a739 & c739) | (b_inv739 & c739);
  wire s740, sub740, and740, or740;
  wire b_inv740;
  assign b_inv740 = ~b740;
  assign s740  = a740 ^ b740 ^ c740;
  assign sub740 = a740 ^ b_inv740 ^ c740;
  assign and740 = a740 & b740;
  assign or740  = a740 | b740;
  assign c741 = (a740 & b740) | (a740 & c740) | (b740 & c740);
  wire c_sub741;
  assign c_sub741 = (a740 & b_inv740) | (a740 & c740) | (b_inv740 & c740);
  wire s741, sub741, and741, or741;
  wire b_inv741;
  assign b_inv741 = ~b741;
  assign s741  = a741 ^ b741 ^ c741;
  assign sub741 = a741 ^ b_inv741 ^ c741;
  assign and741 = a741 & b741;
  assign or741  = a741 | b741;
  assign c742 = (a741 & b741) | (a741 & c741) | (b741 & c741);
  wire c_sub742;
  assign c_sub742 = (a741 & b_inv741) | (a741 & c741) | (b_inv741 & c741);
  wire s742, sub742, and742, or742;
  wire b_inv742;
  assign b_inv742 = ~b742;
  assign s742  = a742 ^ b742 ^ c742;
  assign sub742 = a742 ^ b_inv742 ^ c742;
  assign and742 = a742 & b742;
  assign or742  = a742 | b742;
  assign c743 = (a742 & b742) | (a742 & c742) | (b742 & c742);
  wire c_sub743;
  assign c_sub743 = (a742 & b_inv742) | (a742 & c742) | (b_inv742 & c742);
  wire s743, sub743, and743, or743;
  wire b_inv743;
  assign b_inv743 = ~b743;
  assign s743  = a743 ^ b743 ^ c743;
  assign sub743 = a743 ^ b_inv743 ^ c743;
  assign and743 = a743 & b743;
  assign or743  = a743 | b743;
  assign c744 = (a743 & b743) | (a743 & c743) | (b743 & c743);
  wire c_sub744;
  assign c_sub744 = (a743 & b_inv743) | (a743 & c743) | (b_inv743 & c743);
  wire s744, sub744, and744, or744;
  wire b_inv744;
  assign b_inv744 = ~b744;
  assign s744  = a744 ^ b744 ^ c744;
  assign sub744 = a744 ^ b_inv744 ^ c744;
  assign and744 = a744 & b744;
  assign or744  = a744 | b744;
  assign c745 = (a744 & b744) | (a744 & c744) | (b744 & c744);
  wire c_sub745;
  assign c_sub745 = (a744 & b_inv744) | (a744 & c744) | (b_inv744 & c744);
  wire s745, sub745, and745, or745;
  wire b_inv745;
  assign b_inv745 = ~b745;
  assign s745  = a745 ^ b745 ^ c745;
  assign sub745 = a745 ^ b_inv745 ^ c745;
  assign and745 = a745 & b745;
  assign or745  = a745 | b745;
  assign c746 = (a745 & b745) | (a745 & c745) | (b745 & c745);
  wire c_sub746;
  assign c_sub746 = (a745 & b_inv745) | (a745 & c745) | (b_inv745 & c745);
  wire s746, sub746, and746, or746;
  wire b_inv746;
  assign b_inv746 = ~b746;
  assign s746  = a746 ^ b746 ^ c746;
  assign sub746 = a746 ^ b_inv746 ^ c746;
  assign and746 = a746 & b746;
  assign or746  = a746 | b746;
  assign c747 = (a746 & b746) | (a746 & c746) | (b746 & c746);
  wire c_sub747;
  assign c_sub747 = (a746 & b_inv746) | (a746 & c746) | (b_inv746 & c746);
  wire s747, sub747, and747, or747;
  wire b_inv747;
  assign b_inv747 = ~b747;
  assign s747  = a747 ^ b747 ^ c747;
  assign sub747 = a747 ^ b_inv747 ^ c747;
  assign and747 = a747 & b747;
  assign or747  = a747 | b747;
  assign c748 = (a747 & b747) | (a747 & c747) | (b747 & c747);
  wire c_sub748;
  assign c_sub748 = (a747 & b_inv747) | (a747 & c747) | (b_inv747 & c747);
  wire s748, sub748, and748, or748;
  wire b_inv748;
  assign b_inv748 = ~b748;
  assign s748  = a748 ^ b748 ^ c748;
  assign sub748 = a748 ^ b_inv748 ^ c748;
  assign and748 = a748 & b748;
  assign or748  = a748 | b748;
  assign c749 = (a748 & b748) | (a748 & c748) | (b748 & c748);
  wire c_sub749;
  assign c_sub749 = (a748 & b_inv748) | (a748 & c748) | (b_inv748 & c748);
  wire s749, sub749, and749, or749;
  wire b_inv749;
  assign b_inv749 = ~b749;
  assign s749  = a749 ^ b749 ^ c749;
  assign sub749 = a749 ^ b_inv749 ^ c749;
  assign and749 = a749 & b749;
  assign or749  = a749 | b749;
  assign c750 = (a749 & b749) | (a749 & c749) | (b749 & c749);
  wire c_sub750;
  assign c_sub750 = (a749 & b_inv749) | (a749 & c749) | (b_inv749 & c749);
  wire s750, sub750, and750, or750;
  wire b_inv750;
  assign b_inv750 = ~b750;
  assign s750  = a750 ^ b750 ^ c750;
  assign sub750 = a750 ^ b_inv750 ^ c750;
  assign and750 = a750 & b750;
  assign or750  = a750 | b750;
  assign c751 = (a750 & b750) | (a750 & c750) | (b750 & c750);
  wire c_sub751;
  assign c_sub751 = (a750 & b_inv750) | (a750 & c750) | (b_inv750 & c750);
  wire s751, sub751, and751, or751;
  wire b_inv751;
  assign b_inv751 = ~b751;
  assign s751  = a751 ^ b751 ^ c751;
  assign sub751 = a751 ^ b_inv751 ^ c751;
  assign and751 = a751 & b751;
  assign or751  = a751 | b751;
  assign c752 = (a751 & b751) | (a751 & c751) | (b751 & c751);
  wire c_sub752;
  assign c_sub752 = (a751 & b_inv751) | (a751 & c751) | (b_inv751 & c751);
  wire s752, sub752, and752, or752;
  wire b_inv752;
  assign b_inv752 = ~b752;
  assign s752  = a752 ^ b752 ^ c752;
  assign sub752 = a752 ^ b_inv752 ^ c752;
  assign and752 = a752 & b752;
  assign or752  = a752 | b752;
  assign c753 = (a752 & b752) | (a752 & c752) | (b752 & c752);
  wire c_sub753;
  assign c_sub753 = (a752 & b_inv752) | (a752 & c752) | (b_inv752 & c752);
  wire s753, sub753, and753, or753;
  wire b_inv753;
  assign b_inv753 = ~b753;
  assign s753  = a753 ^ b753 ^ c753;
  assign sub753 = a753 ^ b_inv753 ^ c753;
  assign and753 = a753 & b753;
  assign or753  = a753 | b753;
  assign c754 = (a753 & b753) | (a753 & c753) | (b753 & c753);
  wire c_sub754;
  assign c_sub754 = (a753 & b_inv753) | (a753 & c753) | (b_inv753 & c753);
  wire s754, sub754, and754, or754;
  wire b_inv754;
  assign b_inv754 = ~b754;
  assign s754  = a754 ^ b754 ^ c754;
  assign sub754 = a754 ^ b_inv754 ^ c754;
  assign and754 = a754 & b754;
  assign or754  = a754 | b754;
  assign c755 = (a754 & b754) | (a754 & c754) | (b754 & c754);
  wire c_sub755;
  assign c_sub755 = (a754 & b_inv754) | (a754 & c754) | (b_inv754 & c754);
  wire s755, sub755, and755, or755;
  wire b_inv755;
  assign b_inv755 = ~b755;
  assign s755  = a755 ^ b755 ^ c755;
  assign sub755 = a755 ^ b_inv755 ^ c755;
  assign and755 = a755 & b755;
  assign or755  = a755 | b755;
  assign c756 = (a755 & b755) | (a755 & c755) | (b755 & c755);
  wire c_sub756;
  assign c_sub756 = (a755 & b_inv755) | (a755 & c755) | (b_inv755 & c755);
  wire s756, sub756, and756, or756;
  wire b_inv756;
  assign b_inv756 = ~b756;
  assign s756  = a756 ^ b756 ^ c756;
  assign sub756 = a756 ^ b_inv756 ^ c756;
  assign and756 = a756 & b756;
  assign or756  = a756 | b756;
  assign c757 = (a756 & b756) | (a756 & c756) | (b756 & c756);
  wire c_sub757;
  assign c_sub757 = (a756 & b_inv756) | (a756 & c756) | (b_inv756 & c756);
  wire s757, sub757, and757, or757;
  wire b_inv757;
  assign b_inv757 = ~b757;
  assign s757  = a757 ^ b757 ^ c757;
  assign sub757 = a757 ^ b_inv757 ^ c757;
  assign and757 = a757 & b757;
  assign or757  = a757 | b757;
  assign c758 = (a757 & b757) | (a757 & c757) | (b757 & c757);
  wire c_sub758;
  assign c_sub758 = (a757 & b_inv757) | (a757 & c757) | (b_inv757 & c757);
  wire s758, sub758, and758, or758;
  wire b_inv758;
  assign b_inv758 = ~b758;
  assign s758  = a758 ^ b758 ^ c758;
  assign sub758 = a758 ^ b_inv758 ^ c758;
  assign and758 = a758 & b758;
  assign or758  = a758 | b758;
  assign c759 = (a758 & b758) | (a758 & c758) | (b758 & c758);
  wire c_sub759;
  assign c_sub759 = (a758 & b_inv758) | (a758 & c758) | (b_inv758 & c758);
  wire s759, sub759, and759, or759;
  wire b_inv759;
  assign b_inv759 = ~b759;
  assign s759  = a759 ^ b759 ^ c759;
  assign sub759 = a759 ^ b_inv759 ^ c759;
  assign and759 = a759 & b759;
  assign or759  = a759 | b759;
  assign c760 = (a759 & b759) | (a759 & c759) | (b759 & c759);
  wire c_sub760;
  assign c_sub760 = (a759 & b_inv759) | (a759 & c759) | (b_inv759 & c759);
  wire s760, sub760, and760, or760;
  wire b_inv760;
  assign b_inv760 = ~b760;
  assign s760  = a760 ^ b760 ^ c760;
  assign sub760 = a760 ^ b_inv760 ^ c760;
  assign and760 = a760 & b760;
  assign or760  = a760 | b760;
  assign c761 = (a760 & b760) | (a760 & c760) | (b760 & c760);
  wire c_sub761;
  assign c_sub761 = (a760 & b_inv760) | (a760 & c760) | (b_inv760 & c760);
  wire s761, sub761, and761, or761;
  wire b_inv761;
  assign b_inv761 = ~b761;
  assign s761  = a761 ^ b761 ^ c761;
  assign sub761 = a761 ^ b_inv761 ^ c761;
  assign and761 = a761 & b761;
  assign or761  = a761 | b761;
  assign c762 = (a761 & b761) | (a761 & c761) | (b761 & c761);
  wire c_sub762;
  assign c_sub762 = (a761 & b_inv761) | (a761 & c761) | (b_inv761 & c761);
  wire s762, sub762, and762, or762;
  wire b_inv762;
  assign b_inv762 = ~b762;
  assign s762  = a762 ^ b762 ^ c762;
  assign sub762 = a762 ^ b_inv762 ^ c762;
  assign and762 = a762 & b762;
  assign or762  = a762 | b762;
  assign c763 = (a762 & b762) | (a762 & c762) | (b762 & c762);
  wire c_sub763;
  assign c_sub763 = (a762 & b_inv762) | (a762 & c762) | (b_inv762 & c762);
  wire s763, sub763, and763, or763;
  wire b_inv763;
  assign b_inv763 = ~b763;
  assign s763  = a763 ^ b763 ^ c763;
  assign sub763 = a763 ^ b_inv763 ^ c763;
  assign and763 = a763 & b763;
  assign or763  = a763 | b763;
  assign c764 = (a763 & b763) | (a763 & c763) | (b763 & c763);
  wire c_sub764;
  assign c_sub764 = (a763 & b_inv763) | (a763 & c763) | (b_inv763 & c763);
  wire s764, sub764, and764, or764;
  wire b_inv764;
  assign b_inv764 = ~b764;
  assign s764  = a764 ^ b764 ^ c764;
  assign sub764 = a764 ^ b_inv764 ^ c764;
  assign and764 = a764 & b764;
  assign or764  = a764 | b764;
  assign c765 = (a764 & b764) | (a764 & c764) | (b764 & c764);
  wire c_sub765;
  assign c_sub765 = (a764 & b_inv764) | (a764 & c764) | (b_inv764 & c764);
  wire s765, sub765, and765, or765;
  wire b_inv765;
  assign b_inv765 = ~b765;
  assign s765  = a765 ^ b765 ^ c765;
  assign sub765 = a765 ^ b_inv765 ^ c765;
  assign and765 = a765 & b765;
  assign or765  = a765 | b765;
  assign c766 = (a765 & b765) | (a765 & c765) | (b765 & c765);
  wire c_sub766;
  assign c_sub766 = (a765 & b_inv765) | (a765 & c765) | (b_inv765 & c765);
  wire s766, sub766, and766, or766;
  wire b_inv766;
  assign b_inv766 = ~b766;
  assign s766  = a766 ^ b766 ^ c766;
  assign sub766 = a766 ^ b_inv766 ^ c766;
  assign and766 = a766 & b766;
  assign or766  = a766 | b766;
  assign c767 = (a766 & b766) | (a766 & c766) | (b766 & c766);
  wire c_sub767;
  assign c_sub767 = (a766 & b_inv766) | (a766 & c766) | (b_inv766 & c766);
  wire s767, sub767, and767, or767;
  wire b_inv767;
  assign b_inv767 = ~b767;
  assign s767  = a767 ^ b767 ^ c767;
  assign sub767 = a767 ^ b_inv767 ^ c767;
  assign and767 = a767 & b767;
  assign or767  = a767 | b767;
  assign c768 = (a767 & b767) | (a767 & c767) | (b767 & c767);
  wire c_sub768;
  assign c_sub768 = (a767 & b_inv767) | (a767 & c767) | (b_inv767 & c767);
  wire s768, sub768, and768, or768;
  wire b_inv768;
  assign b_inv768 = ~b768;
  assign s768  = a768 ^ b768 ^ c768;
  assign sub768 = a768 ^ b_inv768 ^ c768;
  assign and768 = a768 & b768;
  assign or768  = a768 | b768;
  assign c769 = (a768 & b768) | (a768 & c768) | (b768 & c768);
  wire c_sub769;
  assign c_sub769 = (a768 & b_inv768) | (a768 & c768) | (b_inv768 & c768);
  wire s769, sub769, and769, or769;
  wire b_inv769;
  assign b_inv769 = ~b769;
  assign s769  = a769 ^ b769 ^ c769;
  assign sub769 = a769 ^ b_inv769 ^ c769;
  assign and769 = a769 & b769;
  assign or769  = a769 | b769;
  assign c770 = (a769 & b769) | (a769 & c769) | (b769 & c769);
  wire c_sub770;
  assign c_sub770 = (a769 & b_inv769) | (a769 & c769) | (b_inv769 & c769);
  wire s770, sub770, and770, or770;
  wire b_inv770;
  assign b_inv770 = ~b770;
  assign s770  = a770 ^ b770 ^ c770;
  assign sub770 = a770 ^ b_inv770 ^ c770;
  assign and770 = a770 & b770;
  assign or770  = a770 | b770;
  assign c771 = (a770 & b770) | (a770 & c770) | (b770 & c770);
  wire c_sub771;
  assign c_sub771 = (a770 & b_inv770) | (a770 & c770) | (b_inv770 & c770);
  wire s771, sub771, and771, or771;
  wire b_inv771;
  assign b_inv771 = ~b771;
  assign s771  = a771 ^ b771 ^ c771;
  assign sub771 = a771 ^ b_inv771 ^ c771;
  assign and771 = a771 & b771;
  assign or771  = a771 | b771;
  assign c772 = (a771 & b771) | (a771 & c771) | (b771 & c771);
  wire c_sub772;
  assign c_sub772 = (a771 & b_inv771) | (a771 & c771) | (b_inv771 & c771);
  wire s772, sub772, and772, or772;
  wire b_inv772;
  assign b_inv772 = ~b772;
  assign s772  = a772 ^ b772 ^ c772;
  assign sub772 = a772 ^ b_inv772 ^ c772;
  assign and772 = a772 & b772;
  assign or772  = a772 | b772;
  assign c773 = (a772 & b772) | (a772 & c772) | (b772 & c772);
  wire c_sub773;
  assign c_sub773 = (a772 & b_inv772) | (a772 & c772) | (b_inv772 & c772);
  wire s773, sub773, and773, or773;
  wire b_inv773;
  assign b_inv773 = ~b773;
  assign s773  = a773 ^ b773 ^ c773;
  assign sub773 = a773 ^ b_inv773 ^ c773;
  assign and773 = a773 & b773;
  assign or773  = a773 | b773;
  assign c774 = (a773 & b773) | (a773 & c773) | (b773 & c773);
  wire c_sub774;
  assign c_sub774 = (a773 & b_inv773) | (a773 & c773) | (b_inv773 & c773);
  wire s774, sub774, and774, or774;
  wire b_inv774;
  assign b_inv774 = ~b774;
  assign s774  = a774 ^ b774 ^ c774;
  assign sub774 = a774 ^ b_inv774 ^ c774;
  assign and774 = a774 & b774;
  assign or774  = a774 | b774;
  assign c775 = (a774 & b774) | (a774 & c774) | (b774 & c774);
  wire c_sub775;
  assign c_sub775 = (a774 & b_inv774) | (a774 & c774) | (b_inv774 & c774);
  wire s775, sub775, and775, or775;
  wire b_inv775;
  assign b_inv775 = ~b775;
  assign s775  = a775 ^ b775 ^ c775;
  assign sub775 = a775 ^ b_inv775 ^ c775;
  assign and775 = a775 & b775;
  assign or775  = a775 | b775;
  assign c776 = (a775 & b775) | (a775 & c775) | (b775 & c775);
  wire c_sub776;
  assign c_sub776 = (a775 & b_inv775) | (a775 & c775) | (b_inv775 & c775);
  wire s776, sub776, and776, or776;
  wire b_inv776;
  assign b_inv776 = ~b776;
  assign s776  = a776 ^ b776 ^ c776;
  assign sub776 = a776 ^ b_inv776 ^ c776;
  assign and776 = a776 & b776;
  assign or776  = a776 | b776;
  assign c777 = (a776 & b776) | (a776 & c776) | (b776 & c776);
  wire c_sub777;
  assign c_sub777 = (a776 & b_inv776) | (a776 & c776) | (b_inv776 & c776);
  wire s777, sub777, and777, or777;
  wire b_inv777;
  assign b_inv777 = ~b777;
  assign s777  = a777 ^ b777 ^ c777;
  assign sub777 = a777 ^ b_inv777 ^ c777;
  assign and777 = a777 & b777;
  assign or777  = a777 | b777;
  assign c778 = (a777 & b777) | (a777 & c777) | (b777 & c777);
  wire c_sub778;
  assign c_sub778 = (a777 & b_inv777) | (a777 & c777) | (b_inv777 & c777);
  wire s778, sub778, and778, or778;
  wire b_inv778;
  assign b_inv778 = ~b778;
  assign s778  = a778 ^ b778 ^ c778;
  assign sub778 = a778 ^ b_inv778 ^ c778;
  assign and778 = a778 & b778;
  assign or778  = a778 | b778;
  assign c779 = (a778 & b778) | (a778 & c778) | (b778 & c778);
  wire c_sub779;
  assign c_sub779 = (a778 & b_inv778) | (a778 & c778) | (b_inv778 & c778);
  wire s779, sub779, and779, or779;
  wire b_inv779;
  assign b_inv779 = ~b779;
  assign s779  = a779 ^ b779 ^ c779;
  assign sub779 = a779 ^ b_inv779 ^ c779;
  assign and779 = a779 & b779;
  assign or779  = a779 | b779;
  assign c780 = (a779 & b779) | (a779 & c779) | (b779 & c779);
  wire c_sub780;
  assign c_sub780 = (a779 & b_inv779) | (a779 & c779) | (b_inv779 & c779);
  wire s780, sub780, and780, or780;
  wire b_inv780;
  assign b_inv780 = ~b780;
  assign s780  = a780 ^ b780 ^ c780;
  assign sub780 = a780 ^ b_inv780 ^ c780;
  assign and780 = a780 & b780;
  assign or780  = a780 | b780;
  assign c781 = (a780 & b780) | (a780 & c780) | (b780 & c780);
  wire c_sub781;
  assign c_sub781 = (a780 & b_inv780) | (a780 & c780) | (b_inv780 & c780);
  wire s781, sub781, and781, or781;
  wire b_inv781;
  assign b_inv781 = ~b781;
  assign s781  = a781 ^ b781 ^ c781;
  assign sub781 = a781 ^ b_inv781 ^ c781;
  assign and781 = a781 & b781;
  assign or781  = a781 | b781;
  assign c782 = (a781 & b781) | (a781 & c781) | (b781 & c781);
  wire c_sub782;
  assign c_sub782 = (a781 & b_inv781) | (a781 & c781) | (b_inv781 & c781);
  wire s782, sub782, and782, or782;
  wire b_inv782;
  assign b_inv782 = ~b782;
  assign s782  = a782 ^ b782 ^ c782;
  assign sub782 = a782 ^ b_inv782 ^ c782;
  assign and782 = a782 & b782;
  assign or782  = a782 | b782;
  assign c783 = (a782 & b782) | (a782 & c782) | (b782 & c782);
  wire c_sub783;
  assign c_sub783 = (a782 & b_inv782) | (a782 & c782) | (b_inv782 & c782);
  wire s783, sub783, and783, or783;
  wire b_inv783;
  assign b_inv783 = ~b783;
  assign s783  = a783 ^ b783 ^ c783;
  assign sub783 = a783 ^ b_inv783 ^ c783;
  assign and783 = a783 & b783;
  assign or783  = a783 | b783;
  assign c784 = (a783 & b783) | (a783 & c783) | (b783 & c783);
  wire c_sub784;
  assign c_sub784 = (a783 & b_inv783) | (a783 & c783) | (b_inv783 & c783);
  wire s784, sub784, and784, or784;
  wire b_inv784;
  assign b_inv784 = ~b784;
  assign s784  = a784 ^ b784 ^ c784;
  assign sub784 = a784 ^ b_inv784 ^ c784;
  assign and784 = a784 & b784;
  assign or784  = a784 | b784;
  assign c785 = (a784 & b784) | (a784 & c784) | (b784 & c784);
  wire c_sub785;
  assign c_sub785 = (a784 & b_inv784) | (a784 & c784) | (b_inv784 & c784);
  wire s785, sub785, and785, or785;
  wire b_inv785;
  assign b_inv785 = ~b785;
  assign s785  = a785 ^ b785 ^ c785;
  assign sub785 = a785 ^ b_inv785 ^ c785;
  assign and785 = a785 & b785;
  assign or785  = a785 | b785;
  assign c786 = (a785 & b785) | (a785 & c785) | (b785 & c785);
  wire c_sub786;
  assign c_sub786 = (a785 & b_inv785) | (a785 & c785) | (b_inv785 & c785);
  wire s786, sub786, and786, or786;
  wire b_inv786;
  assign b_inv786 = ~b786;
  assign s786  = a786 ^ b786 ^ c786;
  assign sub786 = a786 ^ b_inv786 ^ c786;
  assign and786 = a786 & b786;
  assign or786  = a786 | b786;
  assign c787 = (a786 & b786) | (a786 & c786) | (b786 & c786);
  wire c_sub787;
  assign c_sub787 = (a786 & b_inv786) | (a786 & c786) | (b_inv786 & c786);
  wire s787, sub787, and787, or787;
  wire b_inv787;
  assign b_inv787 = ~b787;
  assign s787  = a787 ^ b787 ^ c787;
  assign sub787 = a787 ^ b_inv787 ^ c787;
  assign and787 = a787 & b787;
  assign or787  = a787 | b787;
  assign c788 = (a787 & b787) | (a787 & c787) | (b787 & c787);
  wire c_sub788;
  assign c_sub788 = (a787 & b_inv787) | (a787 & c787) | (b_inv787 & c787);
  wire s788, sub788, and788, or788;
  wire b_inv788;
  assign b_inv788 = ~b788;
  assign s788  = a788 ^ b788 ^ c788;
  assign sub788 = a788 ^ b_inv788 ^ c788;
  assign and788 = a788 & b788;
  assign or788  = a788 | b788;
  assign c789 = (a788 & b788) | (a788 & c788) | (b788 & c788);
  wire c_sub789;
  assign c_sub789 = (a788 & b_inv788) | (a788 & c788) | (b_inv788 & c788);
  wire s789, sub789, and789, or789;
  wire b_inv789;
  assign b_inv789 = ~b789;
  assign s789  = a789 ^ b789 ^ c789;
  assign sub789 = a789 ^ b_inv789 ^ c789;
  assign and789 = a789 & b789;
  assign or789  = a789 | b789;
  assign c790 = (a789 & b789) | (a789 & c789) | (b789 & c789);
  wire c_sub790;
  assign c_sub790 = (a789 & b_inv789) | (a789 & c789) | (b_inv789 & c789);
  wire s790, sub790, and790, or790;
  wire b_inv790;
  assign b_inv790 = ~b790;
  assign s790  = a790 ^ b790 ^ c790;
  assign sub790 = a790 ^ b_inv790 ^ c790;
  assign and790 = a790 & b790;
  assign or790  = a790 | b790;
  assign c791 = (a790 & b790) | (a790 & c790) | (b790 & c790);
  wire c_sub791;
  assign c_sub791 = (a790 & b_inv790) | (a790 & c790) | (b_inv790 & c790);
  wire s791, sub791, and791, or791;
  wire b_inv791;
  assign b_inv791 = ~b791;
  assign s791  = a791 ^ b791 ^ c791;
  assign sub791 = a791 ^ b_inv791 ^ c791;
  assign and791 = a791 & b791;
  assign or791  = a791 | b791;
  assign c792 = (a791 & b791) | (a791 & c791) | (b791 & c791);
  wire c_sub792;
  assign c_sub792 = (a791 & b_inv791) | (a791 & c791) | (b_inv791 & c791);
  wire s792, sub792, and792, or792;
  wire b_inv792;
  assign b_inv792 = ~b792;
  assign s792  = a792 ^ b792 ^ c792;
  assign sub792 = a792 ^ b_inv792 ^ c792;
  assign and792 = a792 & b792;
  assign or792  = a792 | b792;
  assign c793 = (a792 & b792) | (a792 & c792) | (b792 & c792);
  wire c_sub793;
  assign c_sub793 = (a792 & b_inv792) | (a792 & c792) | (b_inv792 & c792);
  wire s793, sub793, and793, or793;
  wire b_inv793;
  assign b_inv793 = ~b793;
  assign s793  = a793 ^ b793 ^ c793;
  assign sub793 = a793 ^ b_inv793 ^ c793;
  assign and793 = a793 & b793;
  assign or793  = a793 | b793;
  assign c794 = (a793 & b793) | (a793 & c793) | (b793 & c793);
  wire c_sub794;
  assign c_sub794 = (a793 & b_inv793) | (a793 & c793) | (b_inv793 & c793);
  wire s794, sub794, and794, or794;
  wire b_inv794;
  assign b_inv794 = ~b794;
  assign s794  = a794 ^ b794 ^ c794;
  assign sub794 = a794 ^ b_inv794 ^ c794;
  assign and794 = a794 & b794;
  assign or794  = a794 | b794;
  assign c795 = (a794 & b794) | (a794 & c794) | (b794 & c794);
  wire c_sub795;
  assign c_sub795 = (a794 & b_inv794) | (a794 & c794) | (b_inv794 & c794);
  wire s795, sub795, and795, or795;
  wire b_inv795;
  assign b_inv795 = ~b795;
  assign s795  = a795 ^ b795 ^ c795;
  assign sub795 = a795 ^ b_inv795 ^ c795;
  assign and795 = a795 & b795;
  assign or795  = a795 | b795;
  assign c796 = (a795 & b795) | (a795 & c795) | (b795 & c795);
  wire c_sub796;
  assign c_sub796 = (a795 & b_inv795) | (a795 & c795) | (b_inv795 & c795);
  wire s796, sub796, and796, or796;
  wire b_inv796;
  assign b_inv796 = ~b796;
  assign s796  = a796 ^ b796 ^ c796;
  assign sub796 = a796 ^ b_inv796 ^ c796;
  assign and796 = a796 & b796;
  assign or796  = a796 | b796;
  assign c797 = (a796 & b796) | (a796 & c796) | (b796 & c796);
  wire c_sub797;
  assign c_sub797 = (a796 & b_inv796) | (a796 & c796) | (b_inv796 & c796);
  wire s797, sub797, and797, or797;
  wire b_inv797;
  assign b_inv797 = ~b797;
  assign s797  = a797 ^ b797 ^ c797;
  assign sub797 = a797 ^ b_inv797 ^ c797;
  assign and797 = a797 & b797;
  assign or797  = a797 | b797;
  assign c798 = (a797 & b797) | (a797 & c797) | (b797 & c797);
  wire c_sub798;
  assign c_sub798 = (a797 & b_inv797) | (a797 & c797) | (b_inv797 & c797);
  wire s798, sub798, and798, or798;
  wire b_inv798;
  assign b_inv798 = ~b798;
  assign s798  = a798 ^ b798 ^ c798;
  assign sub798 = a798 ^ b_inv798 ^ c798;
  assign and798 = a798 & b798;
  assign or798  = a798 | b798;
  assign c799 = (a798 & b798) | (a798 & c798) | (b798 & c798);
  wire c_sub799;
  assign c_sub799 = (a798 & b_inv798) | (a798 & c798) | (b_inv798 & c798);
  wire s799, sub799, and799, or799;
  wire b_inv799;
  assign b_inv799 = ~b799;
  assign s799  = a799 ^ b799 ^ c799;
  assign sub799 = a799 ^ b_inv799 ^ c799;
  assign and799 = a799 & b799;
  assign or799  = a799 | b799;
  assign c800 = (a799 & b799) | (a799 & c799) | (b799 & c799);
  wire c_sub800;
  assign c_sub800 = (a799 & b_inv799) | (a799 & c799) | (b_inv799 & c799);
  wire s800, sub800, and800, or800;
  wire b_inv800;
  assign b_inv800 = ~b800;
  assign s800  = a800 ^ b800 ^ c800;
  assign sub800 = a800 ^ b_inv800 ^ c800;
  assign and800 = a800 & b800;
  assign or800  = a800 | b800;
  assign c801 = (a800 & b800) | (a800 & c800) | (b800 & c800);
  wire c_sub801;
  assign c_sub801 = (a800 & b_inv800) | (a800 & c800) | (b_inv800 & c800);
  wire s801, sub801, and801, or801;
  wire b_inv801;
  assign b_inv801 = ~b801;
  assign s801  = a801 ^ b801 ^ c801;
  assign sub801 = a801 ^ b_inv801 ^ c801;
  assign and801 = a801 & b801;
  assign or801  = a801 | b801;
  assign c802 = (a801 & b801) | (a801 & c801) | (b801 & c801);
  wire c_sub802;
  assign c_sub802 = (a801 & b_inv801) | (a801 & c801) | (b_inv801 & c801);
  wire s802, sub802, and802, or802;
  wire b_inv802;
  assign b_inv802 = ~b802;
  assign s802  = a802 ^ b802 ^ c802;
  assign sub802 = a802 ^ b_inv802 ^ c802;
  assign and802 = a802 & b802;
  assign or802  = a802 | b802;
  assign c803 = (a802 & b802) | (a802 & c802) | (b802 & c802);
  wire c_sub803;
  assign c_sub803 = (a802 & b_inv802) | (a802 & c802) | (b_inv802 & c802);
  wire s803, sub803, and803, or803;
  wire b_inv803;
  assign b_inv803 = ~b803;
  assign s803  = a803 ^ b803 ^ c803;
  assign sub803 = a803 ^ b_inv803 ^ c803;
  assign and803 = a803 & b803;
  assign or803  = a803 | b803;
  assign c804 = (a803 & b803) | (a803 & c803) | (b803 & c803);
  wire c_sub804;
  assign c_sub804 = (a803 & b_inv803) | (a803 & c803) | (b_inv803 & c803);
  wire s804, sub804, and804, or804;
  wire b_inv804;
  assign b_inv804 = ~b804;
  assign s804  = a804 ^ b804 ^ c804;
  assign sub804 = a804 ^ b_inv804 ^ c804;
  assign and804 = a804 & b804;
  assign or804  = a804 | b804;
  assign c805 = (a804 & b804) | (a804 & c804) | (b804 & c804);
  wire c_sub805;
  assign c_sub805 = (a804 & b_inv804) | (a804 & c804) | (b_inv804 & c804);
  wire s805, sub805, and805, or805;
  wire b_inv805;
  assign b_inv805 = ~b805;
  assign s805  = a805 ^ b805 ^ c805;
  assign sub805 = a805 ^ b_inv805 ^ c805;
  assign and805 = a805 & b805;
  assign or805  = a805 | b805;
  assign c806 = (a805 & b805) | (a805 & c805) | (b805 & c805);
  wire c_sub806;
  assign c_sub806 = (a805 & b_inv805) | (a805 & c805) | (b_inv805 & c805);
  wire s806, sub806, and806, or806;
  wire b_inv806;
  assign b_inv806 = ~b806;
  assign s806  = a806 ^ b806 ^ c806;
  assign sub806 = a806 ^ b_inv806 ^ c806;
  assign and806 = a806 & b806;
  assign or806  = a806 | b806;
  assign c807 = (a806 & b806) | (a806 & c806) | (b806 & c806);
  wire c_sub807;
  assign c_sub807 = (a806 & b_inv806) | (a806 & c806) | (b_inv806 & c806);
  wire s807, sub807, and807, or807;
  wire b_inv807;
  assign b_inv807 = ~b807;
  assign s807  = a807 ^ b807 ^ c807;
  assign sub807 = a807 ^ b_inv807 ^ c807;
  assign and807 = a807 & b807;
  assign or807  = a807 | b807;
  assign c808 = (a807 & b807) | (a807 & c807) | (b807 & c807);
  wire c_sub808;
  assign c_sub808 = (a807 & b_inv807) | (a807 & c807) | (b_inv807 & c807);
  wire s808, sub808, and808, or808;
  wire b_inv808;
  assign b_inv808 = ~b808;
  assign s808  = a808 ^ b808 ^ c808;
  assign sub808 = a808 ^ b_inv808 ^ c808;
  assign and808 = a808 & b808;
  assign or808  = a808 | b808;
  assign c809 = (a808 & b808) | (a808 & c808) | (b808 & c808);
  wire c_sub809;
  assign c_sub809 = (a808 & b_inv808) | (a808 & c808) | (b_inv808 & c808);
  wire s809, sub809, and809, or809;
  wire b_inv809;
  assign b_inv809 = ~b809;
  assign s809  = a809 ^ b809 ^ c809;
  assign sub809 = a809 ^ b_inv809 ^ c809;
  assign and809 = a809 & b809;
  assign or809  = a809 | b809;
  assign c810 = (a809 & b809) | (a809 & c809) | (b809 & c809);
  wire c_sub810;
  assign c_sub810 = (a809 & b_inv809) | (a809 & c809) | (b_inv809 & c809);
  wire s810, sub810, and810, or810;
  wire b_inv810;
  assign b_inv810 = ~b810;
  assign s810  = a810 ^ b810 ^ c810;
  assign sub810 = a810 ^ b_inv810 ^ c810;
  assign and810 = a810 & b810;
  assign or810  = a810 | b810;
  assign c811 = (a810 & b810) | (a810 & c810) | (b810 & c810);
  wire c_sub811;
  assign c_sub811 = (a810 & b_inv810) | (a810 & c810) | (b_inv810 & c810);
  wire s811, sub811, and811, or811;
  wire b_inv811;
  assign b_inv811 = ~b811;
  assign s811  = a811 ^ b811 ^ c811;
  assign sub811 = a811 ^ b_inv811 ^ c811;
  assign and811 = a811 & b811;
  assign or811  = a811 | b811;
  assign c812 = (a811 & b811) | (a811 & c811) | (b811 & c811);
  wire c_sub812;
  assign c_sub812 = (a811 & b_inv811) | (a811 & c811) | (b_inv811 & c811);
  wire s812, sub812, and812, or812;
  wire b_inv812;
  assign b_inv812 = ~b812;
  assign s812  = a812 ^ b812 ^ c812;
  assign sub812 = a812 ^ b_inv812 ^ c812;
  assign and812 = a812 & b812;
  assign or812  = a812 | b812;
  assign c813 = (a812 & b812) | (a812 & c812) | (b812 & c812);
  wire c_sub813;
  assign c_sub813 = (a812 & b_inv812) | (a812 & c812) | (b_inv812 & c812);
  wire s813, sub813, and813, or813;
  wire b_inv813;
  assign b_inv813 = ~b813;
  assign s813  = a813 ^ b813 ^ c813;
  assign sub813 = a813 ^ b_inv813 ^ c813;
  assign and813 = a813 & b813;
  assign or813  = a813 | b813;
  assign c814 = (a813 & b813) | (a813 & c813) | (b813 & c813);
  wire c_sub814;
  assign c_sub814 = (a813 & b_inv813) | (a813 & c813) | (b_inv813 & c813);
  wire s814, sub814, and814, or814;
  wire b_inv814;
  assign b_inv814 = ~b814;
  assign s814  = a814 ^ b814 ^ c814;
  assign sub814 = a814 ^ b_inv814 ^ c814;
  assign and814 = a814 & b814;
  assign or814  = a814 | b814;
  assign c815 = (a814 & b814) | (a814 & c814) | (b814 & c814);
  wire c_sub815;
  assign c_sub815 = (a814 & b_inv814) | (a814 & c814) | (b_inv814 & c814);
  wire s815, sub815, and815, or815;
  wire b_inv815;
  assign b_inv815 = ~b815;
  assign s815  = a815 ^ b815 ^ c815;
  assign sub815 = a815 ^ b_inv815 ^ c815;
  assign and815 = a815 & b815;
  assign or815  = a815 | b815;
  assign c816 = (a815 & b815) | (a815 & c815) | (b815 & c815);
  wire c_sub816;
  assign c_sub816 = (a815 & b_inv815) | (a815 & c815) | (b_inv815 & c815);
  wire s816, sub816, and816, or816;
  wire b_inv816;
  assign b_inv816 = ~b816;
  assign s816  = a816 ^ b816 ^ c816;
  assign sub816 = a816 ^ b_inv816 ^ c816;
  assign and816 = a816 & b816;
  assign or816  = a816 | b816;
  assign c817 = (a816 & b816) | (a816 & c816) | (b816 & c816);
  wire c_sub817;
  assign c_sub817 = (a816 & b_inv816) | (a816 & c816) | (b_inv816 & c816);
  wire s817, sub817, and817, or817;
  wire b_inv817;
  assign b_inv817 = ~b817;
  assign s817  = a817 ^ b817 ^ c817;
  assign sub817 = a817 ^ b_inv817 ^ c817;
  assign and817 = a817 & b817;
  assign or817  = a817 | b817;
  assign c818 = (a817 & b817) | (a817 & c817) | (b817 & c817);
  wire c_sub818;
  assign c_sub818 = (a817 & b_inv817) | (a817 & c817) | (b_inv817 & c817);
  wire s818, sub818, and818, or818;
  wire b_inv818;
  assign b_inv818 = ~b818;
  assign s818  = a818 ^ b818 ^ c818;
  assign sub818 = a818 ^ b_inv818 ^ c818;
  assign and818 = a818 & b818;
  assign or818  = a818 | b818;
  assign c819 = (a818 & b818) | (a818 & c818) | (b818 & c818);
  wire c_sub819;
  assign c_sub819 = (a818 & b_inv818) | (a818 & c818) | (b_inv818 & c818);
  wire s819, sub819, and819, or819;
  wire b_inv819;
  assign b_inv819 = ~b819;
  assign s819  = a819 ^ b819 ^ c819;
  assign sub819 = a819 ^ b_inv819 ^ c819;
  assign and819 = a819 & b819;
  assign or819  = a819 | b819;
  assign c820 = (a819 & b819) | (a819 & c819) | (b819 & c819);
  wire c_sub820;
  assign c_sub820 = (a819 & b_inv819) | (a819 & c819) | (b_inv819 & c819);
  wire s820, sub820, and820, or820;
  wire b_inv820;
  assign b_inv820 = ~b820;
  assign s820  = a820 ^ b820 ^ c820;
  assign sub820 = a820 ^ b_inv820 ^ c820;
  assign and820 = a820 & b820;
  assign or820  = a820 | b820;
  assign c821 = (a820 & b820) | (a820 & c820) | (b820 & c820);
  wire c_sub821;
  assign c_sub821 = (a820 & b_inv820) | (a820 & c820) | (b_inv820 & c820);
  wire s821, sub821, and821, or821;
  wire b_inv821;
  assign b_inv821 = ~b821;
  assign s821  = a821 ^ b821 ^ c821;
  assign sub821 = a821 ^ b_inv821 ^ c821;
  assign and821 = a821 & b821;
  assign or821  = a821 | b821;
  assign c822 = (a821 & b821) | (a821 & c821) | (b821 & c821);
  wire c_sub822;
  assign c_sub822 = (a821 & b_inv821) | (a821 & c821) | (b_inv821 & c821);
  wire s822, sub822, and822, or822;
  wire b_inv822;
  assign b_inv822 = ~b822;
  assign s822  = a822 ^ b822 ^ c822;
  assign sub822 = a822 ^ b_inv822 ^ c822;
  assign and822 = a822 & b822;
  assign or822  = a822 | b822;
  assign c823 = (a822 & b822) | (a822 & c822) | (b822 & c822);
  wire c_sub823;
  assign c_sub823 = (a822 & b_inv822) | (a822 & c822) | (b_inv822 & c822);
  wire s823, sub823, and823, or823;
  wire b_inv823;
  assign b_inv823 = ~b823;
  assign s823  = a823 ^ b823 ^ c823;
  assign sub823 = a823 ^ b_inv823 ^ c823;
  assign and823 = a823 & b823;
  assign or823  = a823 | b823;
  assign c824 = (a823 & b823) | (a823 & c823) | (b823 & c823);
  wire c_sub824;
  assign c_sub824 = (a823 & b_inv823) | (a823 & c823) | (b_inv823 & c823);
  wire s824, sub824, and824, or824;
  wire b_inv824;
  assign b_inv824 = ~b824;
  assign s824  = a824 ^ b824 ^ c824;
  assign sub824 = a824 ^ b_inv824 ^ c824;
  assign and824 = a824 & b824;
  assign or824  = a824 | b824;
  assign c825 = (a824 & b824) | (a824 & c824) | (b824 & c824);
  wire c_sub825;
  assign c_sub825 = (a824 & b_inv824) | (a824 & c824) | (b_inv824 & c824);
  wire s825, sub825, and825, or825;
  wire b_inv825;
  assign b_inv825 = ~b825;
  assign s825  = a825 ^ b825 ^ c825;
  assign sub825 = a825 ^ b_inv825 ^ c825;
  assign and825 = a825 & b825;
  assign or825  = a825 | b825;
  assign c826 = (a825 & b825) | (a825 & c825) | (b825 & c825);
  wire c_sub826;
  assign c_sub826 = (a825 & b_inv825) | (a825 & c825) | (b_inv825 & c825);
  wire s826, sub826, and826, or826;
  wire b_inv826;
  assign b_inv826 = ~b826;
  assign s826  = a826 ^ b826 ^ c826;
  assign sub826 = a826 ^ b_inv826 ^ c826;
  assign and826 = a826 & b826;
  assign or826  = a826 | b826;
  assign c827 = (a826 & b826) | (a826 & c826) | (b826 & c826);
  wire c_sub827;
  assign c_sub827 = (a826 & b_inv826) | (a826 & c826) | (b_inv826 & c826);
  wire s827, sub827, and827, or827;
  wire b_inv827;
  assign b_inv827 = ~b827;
  assign s827  = a827 ^ b827 ^ c827;
  assign sub827 = a827 ^ b_inv827 ^ c827;
  assign and827 = a827 & b827;
  assign or827  = a827 | b827;
  assign c828 = (a827 & b827) | (a827 & c827) | (b827 & c827);
  wire c_sub828;
  assign c_sub828 = (a827 & b_inv827) | (a827 & c827) | (b_inv827 & c827);
  wire s828, sub828, and828, or828;
  wire b_inv828;
  assign b_inv828 = ~b828;
  assign s828  = a828 ^ b828 ^ c828;
  assign sub828 = a828 ^ b_inv828 ^ c828;
  assign and828 = a828 & b828;
  assign or828  = a828 | b828;
  assign c829 = (a828 & b828) | (a828 & c828) | (b828 & c828);
  wire c_sub829;
  assign c_sub829 = (a828 & b_inv828) | (a828 & c828) | (b_inv828 & c828);
  wire s829, sub829, and829, or829;
  wire b_inv829;
  assign b_inv829 = ~b829;
  assign s829  = a829 ^ b829 ^ c829;
  assign sub829 = a829 ^ b_inv829 ^ c829;
  assign and829 = a829 & b829;
  assign or829  = a829 | b829;
  assign c830 = (a829 & b829) | (a829 & c829) | (b829 & c829);
  wire c_sub830;
  assign c_sub830 = (a829 & b_inv829) | (a829 & c829) | (b_inv829 & c829);
  wire s830, sub830, and830, or830;
  wire b_inv830;
  assign b_inv830 = ~b830;
  assign s830  = a830 ^ b830 ^ c830;
  assign sub830 = a830 ^ b_inv830 ^ c830;
  assign and830 = a830 & b830;
  assign or830  = a830 | b830;
  assign c831 = (a830 & b830) | (a830 & c830) | (b830 & c830);
  wire c_sub831;
  assign c_sub831 = (a830 & b_inv830) | (a830 & c830) | (b_inv830 & c830);
  wire s831, sub831, and831, or831;
  wire b_inv831;
  assign b_inv831 = ~b831;
  assign s831  = a831 ^ b831 ^ c831;
  assign sub831 = a831 ^ b_inv831 ^ c831;
  assign and831 = a831 & b831;
  assign or831  = a831 | b831;
  assign c832 = (a831 & b831) | (a831 & c831) | (b831 & c831);
  wire c_sub832;
  assign c_sub832 = (a831 & b_inv831) | (a831 & c831) | (b_inv831 & c831);
  wire s832, sub832, and832, or832;
  wire b_inv832;
  assign b_inv832 = ~b832;
  assign s832  = a832 ^ b832 ^ c832;
  assign sub832 = a832 ^ b_inv832 ^ c832;
  assign and832 = a832 & b832;
  assign or832  = a832 | b832;
  assign c833 = (a832 & b832) | (a832 & c832) | (b832 & c832);
  wire c_sub833;
  assign c_sub833 = (a832 & b_inv832) | (a832 & c832) | (b_inv832 & c832);
  wire s833, sub833, and833, or833;
  wire b_inv833;
  assign b_inv833 = ~b833;
  assign s833  = a833 ^ b833 ^ c833;
  assign sub833 = a833 ^ b_inv833 ^ c833;
  assign and833 = a833 & b833;
  assign or833  = a833 | b833;
  assign c834 = (a833 & b833) | (a833 & c833) | (b833 & c833);
  wire c_sub834;
  assign c_sub834 = (a833 & b_inv833) | (a833 & c833) | (b_inv833 & c833);
  wire s834, sub834, and834, or834;
  wire b_inv834;
  assign b_inv834 = ~b834;
  assign s834  = a834 ^ b834 ^ c834;
  assign sub834 = a834 ^ b_inv834 ^ c834;
  assign and834 = a834 & b834;
  assign or834  = a834 | b834;
  assign c835 = (a834 & b834) | (a834 & c834) | (b834 & c834);
  wire c_sub835;
  assign c_sub835 = (a834 & b_inv834) | (a834 & c834) | (b_inv834 & c834);
  wire s835, sub835, and835, or835;
  wire b_inv835;
  assign b_inv835 = ~b835;
  assign s835  = a835 ^ b835 ^ c835;
  assign sub835 = a835 ^ b_inv835 ^ c835;
  assign and835 = a835 & b835;
  assign or835  = a835 | b835;
  assign c836 = (a835 & b835) | (a835 & c835) | (b835 & c835);
  wire c_sub836;
  assign c_sub836 = (a835 & b_inv835) | (a835 & c835) | (b_inv835 & c835);
  wire s836, sub836, and836, or836;
  wire b_inv836;
  assign b_inv836 = ~b836;
  assign s836  = a836 ^ b836 ^ c836;
  assign sub836 = a836 ^ b_inv836 ^ c836;
  assign and836 = a836 & b836;
  assign or836  = a836 | b836;
  assign c837 = (a836 & b836) | (a836 & c836) | (b836 & c836);
  wire c_sub837;
  assign c_sub837 = (a836 & b_inv836) | (a836 & c836) | (b_inv836 & c836);
  wire s837, sub837, and837, or837;
  wire b_inv837;
  assign b_inv837 = ~b837;
  assign s837  = a837 ^ b837 ^ c837;
  assign sub837 = a837 ^ b_inv837 ^ c837;
  assign and837 = a837 & b837;
  assign or837  = a837 | b837;
  assign c838 = (a837 & b837) | (a837 & c837) | (b837 & c837);
  wire c_sub838;
  assign c_sub838 = (a837 & b_inv837) | (a837 & c837) | (b_inv837 & c837);
  wire s838, sub838, and838, or838;
  wire b_inv838;
  assign b_inv838 = ~b838;
  assign s838  = a838 ^ b838 ^ c838;
  assign sub838 = a838 ^ b_inv838 ^ c838;
  assign and838 = a838 & b838;
  assign or838  = a838 | b838;
  assign c839 = (a838 & b838) | (a838 & c838) | (b838 & c838);
  wire c_sub839;
  assign c_sub839 = (a838 & b_inv838) | (a838 & c838) | (b_inv838 & c838);
  wire s839, sub839, and839, or839;
  wire b_inv839;
  assign b_inv839 = ~b839;
  assign s839  = a839 ^ b839 ^ c839;
  assign sub839 = a839 ^ b_inv839 ^ c839;
  assign and839 = a839 & b839;
  assign or839  = a839 | b839;
  assign c840 = (a839 & b839) | (a839 & c839) | (b839 & c839);
  wire c_sub840;
  assign c_sub840 = (a839 & b_inv839) | (a839 & c839) | (b_inv839 & c839);
  wire s840, sub840, and840, or840;
  wire b_inv840;
  assign b_inv840 = ~b840;
  assign s840  = a840 ^ b840 ^ c840;
  assign sub840 = a840 ^ b_inv840 ^ c840;
  assign and840 = a840 & b840;
  assign or840  = a840 | b840;
  assign c841 = (a840 & b840) | (a840 & c840) | (b840 & c840);
  wire c_sub841;
  assign c_sub841 = (a840 & b_inv840) | (a840 & c840) | (b_inv840 & c840);
  wire s841, sub841, and841, or841;
  wire b_inv841;
  assign b_inv841 = ~b841;
  assign s841  = a841 ^ b841 ^ c841;
  assign sub841 = a841 ^ b_inv841 ^ c841;
  assign and841 = a841 & b841;
  assign or841  = a841 | b841;
  assign c842 = (a841 & b841) | (a841 & c841) | (b841 & c841);
  wire c_sub842;
  assign c_sub842 = (a841 & b_inv841) | (a841 & c841) | (b_inv841 & c841);
  wire s842, sub842, and842, or842;
  wire b_inv842;
  assign b_inv842 = ~b842;
  assign s842  = a842 ^ b842 ^ c842;
  assign sub842 = a842 ^ b_inv842 ^ c842;
  assign and842 = a842 & b842;
  assign or842  = a842 | b842;
  assign c843 = (a842 & b842) | (a842 & c842) | (b842 & c842);
  wire c_sub843;
  assign c_sub843 = (a842 & b_inv842) | (a842 & c842) | (b_inv842 & c842);
  wire s843, sub843, and843, or843;
  wire b_inv843;
  assign b_inv843 = ~b843;
  assign s843  = a843 ^ b843 ^ c843;
  assign sub843 = a843 ^ b_inv843 ^ c843;
  assign and843 = a843 & b843;
  assign or843  = a843 | b843;
  assign c844 = (a843 & b843) | (a843 & c843) | (b843 & c843);
  wire c_sub844;
  assign c_sub844 = (a843 & b_inv843) | (a843 & c843) | (b_inv843 & c843);
  wire s844, sub844, and844, or844;
  wire b_inv844;
  assign b_inv844 = ~b844;
  assign s844  = a844 ^ b844 ^ c844;
  assign sub844 = a844 ^ b_inv844 ^ c844;
  assign and844 = a844 & b844;
  assign or844  = a844 | b844;
  assign c845 = (a844 & b844) | (a844 & c844) | (b844 & c844);
  wire c_sub845;
  assign c_sub845 = (a844 & b_inv844) | (a844 & c844) | (b_inv844 & c844);
  wire s845, sub845, and845, or845;
  wire b_inv845;
  assign b_inv845 = ~b845;
  assign s845  = a845 ^ b845 ^ c845;
  assign sub845 = a845 ^ b_inv845 ^ c845;
  assign and845 = a845 & b845;
  assign or845  = a845 | b845;
  assign c846 = (a845 & b845) | (a845 & c845) | (b845 & c845);
  wire c_sub846;
  assign c_sub846 = (a845 & b_inv845) | (a845 & c845) | (b_inv845 & c845);
  wire s846, sub846, and846, or846;
  wire b_inv846;
  assign b_inv846 = ~b846;
  assign s846  = a846 ^ b846 ^ c846;
  assign sub846 = a846 ^ b_inv846 ^ c846;
  assign and846 = a846 & b846;
  assign or846  = a846 | b846;
  assign c847 = (a846 & b846) | (a846 & c846) | (b846 & c846);
  wire c_sub847;
  assign c_sub847 = (a846 & b_inv846) | (a846 & c846) | (b_inv846 & c846);
  wire s847, sub847, and847, or847;
  wire b_inv847;
  assign b_inv847 = ~b847;
  assign s847  = a847 ^ b847 ^ c847;
  assign sub847 = a847 ^ b_inv847 ^ c847;
  assign and847 = a847 & b847;
  assign or847  = a847 | b847;
  assign c848 = (a847 & b847) | (a847 & c847) | (b847 & c847);
  wire c_sub848;
  assign c_sub848 = (a847 & b_inv847) | (a847 & c847) | (b_inv847 & c847);
  wire s848, sub848, and848, or848;
  wire b_inv848;
  assign b_inv848 = ~b848;
  assign s848  = a848 ^ b848 ^ c848;
  assign sub848 = a848 ^ b_inv848 ^ c848;
  assign and848 = a848 & b848;
  assign or848  = a848 | b848;
  assign c849 = (a848 & b848) | (a848 & c848) | (b848 & c848);
  wire c_sub849;
  assign c_sub849 = (a848 & b_inv848) | (a848 & c848) | (b_inv848 & c848);
  wire s849, sub849, and849, or849;
  wire b_inv849;
  assign b_inv849 = ~b849;
  assign s849  = a849 ^ b849 ^ c849;
  assign sub849 = a849 ^ b_inv849 ^ c849;
  assign and849 = a849 & b849;
  assign or849  = a849 | b849;
  assign c850 = (a849 & b849) | (a849 & c849) | (b849 & c849);
  wire c_sub850;
  assign c_sub850 = (a849 & b_inv849) | (a849 & c849) | (b_inv849 & c849);
  wire s850, sub850, and850, or850;
  wire b_inv850;
  assign b_inv850 = ~b850;
  assign s850  = a850 ^ b850 ^ c850;
  assign sub850 = a850 ^ b_inv850 ^ c850;
  assign and850 = a850 & b850;
  assign or850  = a850 | b850;
  assign c851 = (a850 & b850) | (a850 & c850) | (b850 & c850);
  wire c_sub851;
  assign c_sub851 = (a850 & b_inv850) | (a850 & c850) | (b_inv850 & c850);
  wire s851, sub851, and851, or851;
  wire b_inv851;
  assign b_inv851 = ~b851;
  assign s851  = a851 ^ b851 ^ c851;
  assign sub851 = a851 ^ b_inv851 ^ c851;
  assign and851 = a851 & b851;
  assign or851  = a851 | b851;
  assign c852 = (a851 & b851) | (a851 & c851) | (b851 & c851);
  wire c_sub852;
  assign c_sub852 = (a851 & b_inv851) | (a851 & c851) | (b_inv851 & c851);
  wire s852, sub852, and852, or852;
  wire b_inv852;
  assign b_inv852 = ~b852;
  assign s852  = a852 ^ b852 ^ c852;
  assign sub852 = a852 ^ b_inv852 ^ c852;
  assign and852 = a852 & b852;
  assign or852  = a852 | b852;
  assign c853 = (a852 & b852) | (a852 & c852) | (b852 & c852);
  wire c_sub853;
  assign c_sub853 = (a852 & b_inv852) | (a852 & c852) | (b_inv852 & c852);
  wire s853, sub853, and853, or853;
  wire b_inv853;
  assign b_inv853 = ~b853;
  assign s853  = a853 ^ b853 ^ c853;
  assign sub853 = a853 ^ b_inv853 ^ c853;
  assign and853 = a853 & b853;
  assign or853  = a853 | b853;
  assign c854 = (a853 & b853) | (a853 & c853) | (b853 & c853);
  wire c_sub854;
  assign c_sub854 = (a853 & b_inv853) | (a853 & c853) | (b_inv853 & c853);
  wire s854, sub854, and854, or854;
  wire b_inv854;
  assign b_inv854 = ~b854;
  assign s854  = a854 ^ b854 ^ c854;
  assign sub854 = a854 ^ b_inv854 ^ c854;
  assign and854 = a854 & b854;
  assign or854  = a854 | b854;
  assign c855 = (a854 & b854) | (a854 & c854) | (b854 & c854);
  wire c_sub855;
  assign c_sub855 = (a854 & b_inv854) | (a854 & c854) | (b_inv854 & c854);
  wire s855, sub855, and855, or855;
  wire b_inv855;
  assign b_inv855 = ~b855;
  assign s855  = a855 ^ b855 ^ c855;
  assign sub855 = a855 ^ b_inv855 ^ c855;
  assign and855 = a855 & b855;
  assign or855  = a855 | b855;
  assign c856 = (a855 & b855) | (a855 & c855) | (b855 & c855);
  wire c_sub856;
  assign c_sub856 = (a855 & b_inv855) | (a855 & c855) | (b_inv855 & c855);
  wire s856, sub856, and856, or856;
  wire b_inv856;
  assign b_inv856 = ~b856;
  assign s856  = a856 ^ b856 ^ c856;
  assign sub856 = a856 ^ b_inv856 ^ c856;
  assign and856 = a856 & b856;
  assign or856  = a856 | b856;
  assign c857 = (a856 & b856) | (a856 & c856) | (b856 & c856);
  wire c_sub857;
  assign c_sub857 = (a856 & b_inv856) | (a856 & c856) | (b_inv856 & c856);
  wire s857, sub857, and857, or857;
  wire b_inv857;
  assign b_inv857 = ~b857;
  assign s857  = a857 ^ b857 ^ c857;
  assign sub857 = a857 ^ b_inv857 ^ c857;
  assign and857 = a857 & b857;
  assign or857  = a857 | b857;
  assign c858 = (a857 & b857) | (a857 & c857) | (b857 & c857);
  wire c_sub858;
  assign c_sub858 = (a857 & b_inv857) | (a857 & c857) | (b_inv857 & c857);
  wire s858, sub858, and858, or858;
  wire b_inv858;
  assign b_inv858 = ~b858;
  assign s858  = a858 ^ b858 ^ c858;
  assign sub858 = a858 ^ b_inv858 ^ c858;
  assign and858 = a858 & b858;
  assign or858  = a858 | b858;
  assign c859 = (a858 & b858) | (a858 & c858) | (b858 & c858);
  wire c_sub859;
  assign c_sub859 = (a858 & b_inv858) | (a858 & c858) | (b_inv858 & c858);
  wire s859, sub859, and859, or859;
  wire b_inv859;
  assign b_inv859 = ~b859;
  assign s859  = a859 ^ b859 ^ c859;
  assign sub859 = a859 ^ b_inv859 ^ c859;
  assign and859 = a859 & b859;
  assign or859  = a859 | b859;
  assign c860 = (a859 & b859) | (a859 & c859) | (b859 & c859);
  wire c_sub860;
  assign c_sub860 = (a859 & b_inv859) | (a859 & c859) | (b_inv859 & c859);
  wire s860, sub860, and860, or860;
  wire b_inv860;
  assign b_inv860 = ~b860;
  assign s860  = a860 ^ b860 ^ c860;
  assign sub860 = a860 ^ b_inv860 ^ c860;
  assign and860 = a860 & b860;
  assign or860  = a860 | b860;
  assign c861 = (a860 & b860) | (a860 & c860) | (b860 & c860);
  wire c_sub861;
  assign c_sub861 = (a860 & b_inv860) | (a860 & c860) | (b_inv860 & c860);
  wire s861, sub861, and861, or861;
  wire b_inv861;
  assign b_inv861 = ~b861;
  assign s861  = a861 ^ b861 ^ c861;
  assign sub861 = a861 ^ b_inv861 ^ c861;
  assign and861 = a861 & b861;
  assign or861  = a861 | b861;
  assign c862 = (a861 & b861) | (a861 & c861) | (b861 & c861);
  wire c_sub862;
  assign c_sub862 = (a861 & b_inv861) | (a861 & c861) | (b_inv861 & c861);
  wire s862, sub862, and862, or862;
  wire b_inv862;
  assign b_inv862 = ~b862;
  assign s862  = a862 ^ b862 ^ c862;
  assign sub862 = a862 ^ b_inv862 ^ c862;
  assign and862 = a862 & b862;
  assign or862  = a862 | b862;
  assign c863 = (a862 & b862) | (a862 & c862) | (b862 & c862);
  wire c_sub863;
  assign c_sub863 = (a862 & b_inv862) | (a862 & c862) | (b_inv862 & c862);
  wire s863, sub863, and863, or863;
  wire b_inv863;
  assign b_inv863 = ~b863;
  assign s863  = a863 ^ b863 ^ c863;
  assign sub863 = a863 ^ b_inv863 ^ c863;
  assign and863 = a863 & b863;
  assign or863  = a863 | b863;
  assign c864 = (a863 & b863) | (a863 & c863) | (b863 & c863);
  wire c_sub864;
  assign c_sub864 = (a863 & b_inv863) | (a863 & c863) | (b_inv863 & c863);
  wire s864, sub864, and864, or864;
  wire b_inv864;
  assign b_inv864 = ~b864;
  assign s864  = a864 ^ b864 ^ c864;
  assign sub864 = a864 ^ b_inv864 ^ c864;
  assign and864 = a864 & b864;
  assign or864  = a864 | b864;
  assign c865 = (a864 & b864) | (a864 & c864) | (b864 & c864);
  wire c_sub865;
  assign c_sub865 = (a864 & b_inv864) | (a864 & c864) | (b_inv864 & c864);
  wire s865, sub865, and865, or865;
  wire b_inv865;
  assign b_inv865 = ~b865;
  assign s865  = a865 ^ b865 ^ c865;
  assign sub865 = a865 ^ b_inv865 ^ c865;
  assign and865 = a865 & b865;
  assign or865  = a865 | b865;
  assign c866 = (a865 & b865) | (a865 & c865) | (b865 & c865);
  wire c_sub866;
  assign c_sub866 = (a865 & b_inv865) | (a865 & c865) | (b_inv865 & c865);
  wire s866, sub866, and866, or866;
  wire b_inv866;
  assign b_inv866 = ~b866;
  assign s866  = a866 ^ b866 ^ c866;
  assign sub866 = a866 ^ b_inv866 ^ c866;
  assign and866 = a866 & b866;
  assign or866  = a866 | b866;
  assign c867 = (a866 & b866) | (a866 & c866) | (b866 & c866);
  wire c_sub867;
  assign c_sub867 = (a866 & b_inv866) | (a866 & c866) | (b_inv866 & c866);
  wire s867, sub867, and867, or867;
  wire b_inv867;
  assign b_inv867 = ~b867;
  assign s867  = a867 ^ b867 ^ c867;
  assign sub867 = a867 ^ b_inv867 ^ c867;
  assign and867 = a867 & b867;
  assign or867  = a867 | b867;
  assign c868 = (a867 & b867) | (a867 & c867) | (b867 & c867);
  wire c_sub868;
  assign c_sub868 = (a867 & b_inv867) | (a867 & c867) | (b_inv867 & c867);
  wire s868, sub868, and868, or868;
  wire b_inv868;
  assign b_inv868 = ~b868;
  assign s868  = a868 ^ b868 ^ c868;
  assign sub868 = a868 ^ b_inv868 ^ c868;
  assign and868 = a868 & b868;
  assign or868  = a868 | b868;
  assign c869 = (a868 & b868) | (a868 & c868) | (b868 & c868);
  wire c_sub869;
  assign c_sub869 = (a868 & b_inv868) | (a868 & c868) | (b_inv868 & c868);
  wire s869, sub869, and869, or869;
  wire b_inv869;
  assign b_inv869 = ~b869;
  assign s869  = a869 ^ b869 ^ c869;
  assign sub869 = a869 ^ b_inv869 ^ c869;
  assign and869 = a869 & b869;
  assign or869  = a869 | b869;
  assign c870 = (a869 & b869) | (a869 & c869) | (b869 & c869);
  wire c_sub870;
  assign c_sub870 = (a869 & b_inv869) | (a869 & c869) | (b_inv869 & c869);
  wire s870, sub870, and870, or870;
  wire b_inv870;
  assign b_inv870 = ~b870;
  assign s870  = a870 ^ b870 ^ c870;
  assign sub870 = a870 ^ b_inv870 ^ c870;
  assign and870 = a870 & b870;
  assign or870  = a870 | b870;
  assign c871 = (a870 & b870) | (a870 & c870) | (b870 & c870);
  wire c_sub871;
  assign c_sub871 = (a870 & b_inv870) | (a870 & c870) | (b_inv870 & c870);
  wire s871, sub871, and871, or871;
  wire b_inv871;
  assign b_inv871 = ~b871;
  assign s871  = a871 ^ b871 ^ c871;
  assign sub871 = a871 ^ b_inv871 ^ c871;
  assign and871 = a871 & b871;
  assign or871  = a871 | b871;
  assign c872 = (a871 & b871) | (a871 & c871) | (b871 & c871);
  wire c_sub872;
  assign c_sub872 = (a871 & b_inv871) | (a871 & c871) | (b_inv871 & c871);
  wire s872, sub872, and872, or872;
  wire b_inv872;
  assign b_inv872 = ~b872;
  assign s872  = a872 ^ b872 ^ c872;
  assign sub872 = a872 ^ b_inv872 ^ c872;
  assign and872 = a872 & b872;
  assign or872  = a872 | b872;
  assign c873 = (a872 & b872) | (a872 & c872) | (b872 & c872);
  wire c_sub873;
  assign c_sub873 = (a872 & b_inv872) | (a872 & c872) | (b_inv872 & c872);
  wire s873, sub873, and873, or873;
  wire b_inv873;
  assign b_inv873 = ~b873;
  assign s873  = a873 ^ b873 ^ c873;
  assign sub873 = a873 ^ b_inv873 ^ c873;
  assign and873 = a873 & b873;
  assign or873  = a873 | b873;
  assign c874 = (a873 & b873) | (a873 & c873) | (b873 & c873);
  wire c_sub874;
  assign c_sub874 = (a873 & b_inv873) | (a873 & c873) | (b_inv873 & c873);
  wire s874, sub874, and874, or874;
  wire b_inv874;
  assign b_inv874 = ~b874;
  assign s874  = a874 ^ b874 ^ c874;
  assign sub874 = a874 ^ b_inv874 ^ c874;
  assign and874 = a874 & b874;
  assign or874  = a874 | b874;
  assign c875 = (a874 & b874) | (a874 & c874) | (b874 & c874);
  wire c_sub875;
  assign c_sub875 = (a874 & b_inv874) | (a874 & c874) | (b_inv874 & c874);
  wire s875, sub875, and875, or875;
  wire b_inv875;
  assign b_inv875 = ~b875;
  assign s875  = a875 ^ b875 ^ c875;
  assign sub875 = a875 ^ b_inv875 ^ c875;
  assign and875 = a875 & b875;
  assign or875  = a875 | b875;
  assign c876 = (a875 & b875) | (a875 & c875) | (b875 & c875);
  wire c_sub876;
  assign c_sub876 = (a875 & b_inv875) | (a875 & c875) | (b_inv875 & c875);
  wire s876, sub876, and876, or876;
  wire b_inv876;
  assign b_inv876 = ~b876;
  assign s876  = a876 ^ b876 ^ c876;
  assign sub876 = a876 ^ b_inv876 ^ c876;
  assign and876 = a876 & b876;
  assign or876  = a876 | b876;
  assign c877 = (a876 & b876) | (a876 & c876) | (b876 & c876);
  wire c_sub877;
  assign c_sub877 = (a876 & b_inv876) | (a876 & c876) | (b_inv876 & c876);
  wire s877, sub877, and877, or877;
  wire b_inv877;
  assign b_inv877 = ~b877;
  assign s877  = a877 ^ b877 ^ c877;
  assign sub877 = a877 ^ b_inv877 ^ c877;
  assign and877 = a877 & b877;
  assign or877  = a877 | b877;
  assign c878 = (a877 & b877) | (a877 & c877) | (b877 & c877);
  wire c_sub878;
  assign c_sub878 = (a877 & b_inv877) | (a877 & c877) | (b_inv877 & c877);
  wire s878, sub878, and878, or878;
  wire b_inv878;
  assign b_inv878 = ~b878;
  assign s878  = a878 ^ b878 ^ c878;
  assign sub878 = a878 ^ b_inv878 ^ c878;
  assign and878 = a878 & b878;
  assign or878  = a878 | b878;
  assign c879 = (a878 & b878) | (a878 & c878) | (b878 & c878);
  wire c_sub879;
  assign c_sub879 = (a878 & b_inv878) | (a878 & c878) | (b_inv878 & c878);
  wire s879, sub879, and879, or879;
  wire b_inv879;
  assign b_inv879 = ~b879;
  assign s879  = a879 ^ b879 ^ c879;
  assign sub879 = a879 ^ b_inv879 ^ c879;
  assign and879 = a879 & b879;
  assign or879  = a879 | b879;
  assign c880 = (a879 & b879) | (a879 & c879) | (b879 & c879);
  wire c_sub880;
  assign c_sub880 = (a879 & b_inv879) | (a879 & c879) | (b_inv879 & c879);
  wire s880, sub880, and880, or880;
  wire b_inv880;
  assign b_inv880 = ~b880;
  assign s880  = a880 ^ b880 ^ c880;
  assign sub880 = a880 ^ b_inv880 ^ c880;
  assign and880 = a880 & b880;
  assign or880  = a880 | b880;
  assign c881 = (a880 & b880) | (a880 & c880) | (b880 & c880);
  wire c_sub881;
  assign c_sub881 = (a880 & b_inv880) | (a880 & c880) | (b_inv880 & c880);
  wire s881, sub881, and881, or881;
  wire b_inv881;
  assign b_inv881 = ~b881;
  assign s881  = a881 ^ b881 ^ c881;
  assign sub881 = a881 ^ b_inv881 ^ c881;
  assign and881 = a881 & b881;
  assign or881  = a881 | b881;
  assign c882 = (a881 & b881) | (a881 & c881) | (b881 & c881);
  wire c_sub882;
  assign c_sub882 = (a881 & b_inv881) | (a881 & c881) | (b_inv881 & c881);
  wire s882, sub882, and882, or882;
  wire b_inv882;
  assign b_inv882 = ~b882;
  assign s882  = a882 ^ b882 ^ c882;
  assign sub882 = a882 ^ b_inv882 ^ c882;
  assign and882 = a882 & b882;
  assign or882  = a882 | b882;
  assign c883 = (a882 & b882) | (a882 & c882) | (b882 & c882);
  wire c_sub883;
  assign c_sub883 = (a882 & b_inv882) | (a882 & c882) | (b_inv882 & c882);
  wire s883, sub883, and883, or883;
  wire b_inv883;
  assign b_inv883 = ~b883;
  assign s883  = a883 ^ b883 ^ c883;
  assign sub883 = a883 ^ b_inv883 ^ c883;
  assign and883 = a883 & b883;
  assign or883  = a883 | b883;
  assign c884 = (a883 & b883) | (a883 & c883) | (b883 & c883);
  wire c_sub884;
  assign c_sub884 = (a883 & b_inv883) | (a883 & c883) | (b_inv883 & c883);
  wire s884, sub884, and884, or884;
  wire b_inv884;
  assign b_inv884 = ~b884;
  assign s884  = a884 ^ b884 ^ c884;
  assign sub884 = a884 ^ b_inv884 ^ c884;
  assign and884 = a884 & b884;
  assign or884  = a884 | b884;
  assign c885 = (a884 & b884) | (a884 & c884) | (b884 & c884);
  wire c_sub885;
  assign c_sub885 = (a884 & b_inv884) | (a884 & c884) | (b_inv884 & c884);
  wire s885, sub885, and885, or885;
  wire b_inv885;
  assign b_inv885 = ~b885;
  assign s885  = a885 ^ b885 ^ c885;
  assign sub885 = a885 ^ b_inv885 ^ c885;
  assign and885 = a885 & b885;
  assign or885  = a885 | b885;
  assign c886 = (a885 & b885) | (a885 & c885) | (b885 & c885);
  wire c_sub886;
  assign c_sub886 = (a885 & b_inv885) | (a885 & c885) | (b_inv885 & c885);
  wire s886, sub886, and886, or886;
  wire b_inv886;
  assign b_inv886 = ~b886;
  assign s886  = a886 ^ b886 ^ c886;
  assign sub886 = a886 ^ b_inv886 ^ c886;
  assign and886 = a886 & b886;
  assign or886  = a886 | b886;
  assign c887 = (a886 & b886) | (a886 & c886) | (b886 & c886);
  wire c_sub887;
  assign c_sub887 = (a886 & b_inv886) | (a886 & c886) | (b_inv886 & c886);
  wire s887, sub887, and887, or887;
  wire b_inv887;
  assign b_inv887 = ~b887;
  assign s887  = a887 ^ b887 ^ c887;
  assign sub887 = a887 ^ b_inv887 ^ c887;
  assign and887 = a887 & b887;
  assign or887  = a887 | b887;
  assign c888 = (a887 & b887) | (a887 & c887) | (b887 & c887);
  wire c_sub888;
  assign c_sub888 = (a887 & b_inv887) | (a887 & c887) | (b_inv887 & c887);
  wire s888, sub888, and888, or888;
  wire b_inv888;
  assign b_inv888 = ~b888;
  assign s888  = a888 ^ b888 ^ c888;
  assign sub888 = a888 ^ b_inv888 ^ c888;
  assign and888 = a888 & b888;
  assign or888  = a888 | b888;
  assign c889 = (a888 & b888) | (a888 & c888) | (b888 & c888);
  wire c_sub889;
  assign c_sub889 = (a888 & b_inv888) | (a888 & c888) | (b_inv888 & c888);
  wire s889, sub889, and889, or889;
  wire b_inv889;
  assign b_inv889 = ~b889;
  assign s889  = a889 ^ b889 ^ c889;
  assign sub889 = a889 ^ b_inv889 ^ c889;
  assign and889 = a889 & b889;
  assign or889  = a889 | b889;
  assign c890 = (a889 & b889) | (a889 & c889) | (b889 & c889);
  wire c_sub890;
  assign c_sub890 = (a889 & b_inv889) | (a889 & c889) | (b_inv889 & c889);
  wire s890, sub890, and890, or890;
  wire b_inv890;
  assign b_inv890 = ~b890;
  assign s890  = a890 ^ b890 ^ c890;
  assign sub890 = a890 ^ b_inv890 ^ c890;
  assign and890 = a890 & b890;
  assign or890  = a890 | b890;
  assign c891 = (a890 & b890) | (a890 & c890) | (b890 & c890);
  wire c_sub891;
  assign c_sub891 = (a890 & b_inv890) | (a890 & c890) | (b_inv890 & c890);
  wire s891, sub891, and891, or891;
  wire b_inv891;
  assign b_inv891 = ~b891;
  assign s891  = a891 ^ b891 ^ c891;
  assign sub891 = a891 ^ b_inv891 ^ c891;
  assign and891 = a891 & b891;
  assign or891  = a891 | b891;
  assign c892 = (a891 & b891) | (a891 & c891) | (b891 & c891);
  wire c_sub892;
  assign c_sub892 = (a891 & b_inv891) | (a891 & c891) | (b_inv891 & c891);
  wire s892, sub892, and892, or892;
  wire b_inv892;
  assign b_inv892 = ~b892;
  assign s892  = a892 ^ b892 ^ c892;
  assign sub892 = a892 ^ b_inv892 ^ c892;
  assign and892 = a892 & b892;
  assign or892  = a892 | b892;
  assign c893 = (a892 & b892) | (a892 & c892) | (b892 & c892);
  wire c_sub893;
  assign c_sub893 = (a892 & b_inv892) | (a892 & c892) | (b_inv892 & c892);
  wire s893, sub893, and893, or893;
  wire b_inv893;
  assign b_inv893 = ~b893;
  assign s893  = a893 ^ b893 ^ c893;
  assign sub893 = a893 ^ b_inv893 ^ c893;
  assign and893 = a893 & b893;
  assign or893  = a893 | b893;
  assign c894 = (a893 & b893) | (a893 & c893) | (b893 & c893);
  wire c_sub894;
  assign c_sub894 = (a893 & b_inv893) | (a893 & c893) | (b_inv893 & c893);
  wire s894, sub894, and894, or894;
  wire b_inv894;
  assign b_inv894 = ~b894;
  assign s894  = a894 ^ b894 ^ c894;
  assign sub894 = a894 ^ b_inv894 ^ c894;
  assign and894 = a894 & b894;
  assign or894  = a894 | b894;
  assign c895 = (a894 & b894) | (a894 & c894) | (b894 & c894);
  wire c_sub895;
  assign c_sub895 = (a894 & b_inv894) | (a894 & c894) | (b_inv894 & c894);
  wire s895, sub895, and895, or895;
  wire b_inv895;
  assign b_inv895 = ~b895;
  assign s895  = a895 ^ b895 ^ c895;
  assign sub895 = a895 ^ b_inv895 ^ c895;
  assign and895 = a895 & b895;
  assign or895  = a895 | b895;
  assign c896 = (a895 & b895) | (a895 & c895) | (b895 & c895);
  wire c_sub896;
  assign c_sub896 = (a895 & b_inv895) | (a895 & c895) | (b_inv895 & c895);
  wire s896, sub896, and896, or896;
  wire b_inv896;
  assign b_inv896 = ~b896;
  assign s896  = a896 ^ b896 ^ c896;
  assign sub896 = a896 ^ b_inv896 ^ c896;
  assign and896 = a896 & b896;
  assign or896  = a896 | b896;
  assign c897 = (a896 & b896) | (a896 & c896) | (b896 & c896);
  wire c_sub897;
  assign c_sub897 = (a896 & b_inv896) | (a896 & c896) | (b_inv896 & c896);
  wire s897, sub897, and897, or897;
  wire b_inv897;
  assign b_inv897 = ~b897;
  assign s897  = a897 ^ b897 ^ c897;
  assign sub897 = a897 ^ b_inv897 ^ c897;
  assign and897 = a897 & b897;
  assign or897  = a897 | b897;
  assign c898 = (a897 & b897) | (a897 & c897) | (b897 & c897);
  wire c_sub898;
  assign c_sub898 = (a897 & b_inv897) | (a897 & c897) | (b_inv897 & c897);
  wire s898, sub898, and898, or898;
  wire b_inv898;
  assign b_inv898 = ~b898;
  assign s898  = a898 ^ b898 ^ c898;
  assign sub898 = a898 ^ b_inv898 ^ c898;
  assign and898 = a898 & b898;
  assign or898  = a898 | b898;
  assign c899 = (a898 & b898) | (a898 & c898) | (b898 & c898);
  wire c_sub899;
  assign c_sub899 = (a898 & b_inv898) | (a898 & c898) | (b_inv898 & c898);
  wire s899, sub899, and899, or899;
  wire b_inv899;
  assign b_inv899 = ~b899;
  assign s899  = a899 ^ b899 ^ c899;
  assign sub899 = a899 ^ b_inv899 ^ c899;
  assign and899 = a899 & b899;
  assign or899  = a899 | b899;
  assign c900 = (a899 & b899) | (a899 & c899) | (b899 & c899);
  wire c_sub900;
  assign c_sub900 = (a899 & b_inv899) | (a899 & c899) | (b_inv899 & c899);
  wire s900, sub900, and900, or900;
  wire b_inv900;
  assign b_inv900 = ~b900;
  assign s900  = a900 ^ b900 ^ c900;
  assign sub900 = a900 ^ b_inv900 ^ c900;
  assign and900 = a900 & b900;
  assign or900  = a900 | b900;
  assign c901 = (a900 & b900) | (a900 & c900) | (b900 & c900);
  wire c_sub901;
  assign c_sub901 = (a900 & b_inv900) | (a900 & c900) | (b_inv900 & c900);
  wire s901, sub901, and901, or901;
  wire b_inv901;
  assign b_inv901 = ~b901;
  assign s901  = a901 ^ b901 ^ c901;
  assign sub901 = a901 ^ b_inv901 ^ c901;
  assign and901 = a901 & b901;
  assign or901  = a901 | b901;
  assign c902 = (a901 & b901) | (a901 & c901) | (b901 & c901);
  wire c_sub902;
  assign c_sub902 = (a901 & b_inv901) | (a901 & c901) | (b_inv901 & c901);
  wire s902, sub902, and902, or902;
  wire b_inv902;
  assign b_inv902 = ~b902;
  assign s902  = a902 ^ b902 ^ c902;
  assign sub902 = a902 ^ b_inv902 ^ c902;
  assign and902 = a902 & b902;
  assign or902  = a902 | b902;
  assign c903 = (a902 & b902) | (a902 & c902) | (b902 & c902);
  wire c_sub903;
  assign c_sub903 = (a902 & b_inv902) | (a902 & c902) | (b_inv902 & c902);
  wire s903, sub903, and903, or903;
  wire b_inv903;
  assign b_inv903 = ~b903;
  assign s903  = a903 ^ b903 ^ c903;
  assign sub903 = a903 ^ b_inv903 ^ c903;
  assign and903 = a903 & b903;
  assign or903  = a903 | b903;
  assign c904 = (a903 & b903) | (a903 & c903) | (b903 & c903);
  wire c_sub904;
  assign c_sub904 = (a903 & b_inv903) | (a903 & c903) | (b_inv903 & c903);
  wire s904, sub904, and904, or904;
  wire b_inv904;
  assign b_inv904 = ~b904;
  assign s904  = a904 ^ b904 ^ c904;
  assign sub904 = a904 ^ b_inv904 ^ c904;
  assign and904 = a904 & b904;
  assign or904  = a904 | b904;
  assign c905 = (a904 & b904) | (a904 & c904) | (b904 & c904);
  wire c_sub905;
  assign c_sub905 = (a904 & b_inv904) | (a904 & c904) | (b_inv904 & c904);
  wire s905, sub905, and905, or905;
  wire b_inv905;
  assign b_inv905 = ~b905;
  assign s905  = a905 ^ b905 ^ c905;
  assign sub905 = a905 ^ b_inv905 ^ c905;
  assign and905 = a905 & b905;
  assign or905  = a905 | b905;
  assign c906 = (a905 & b905) | (a905 & c905) | (b905 & c905);
  wire c_sub906;
  assign c_sub906 = (a905 & b_inv905) | (a905 & c905) | (b_inv905 & c905);
  wire s906, sub906, and906, or906;
  wire b_inv906;
  assign b_inv906 = ~b906;
  assign s906  = a906 ^ b906 ^ c906;
  assign sub906 = a906 ^ b_inv906 ^ c906;
  assign and906 = a906 & b906;
  assign or906  = a906 | b906;
  assign c907 = (a906 & b906) | (a906 & c906) | (b906 & c906);
  wire c_sub907;
  assign c_sub907 = (a906 & b_inv906) | (a906 & c906) | (b_inv906 & c906);
  wire s907, sub907, and907, or907;
  wire b_inv907;
  assign b_inv907 = ~b907;
  assign s907  = a907 ^ b907 ^ c907;
  assign sub907 = a907 ^ b_inv907 ^ c907;
  assign and907 = a907 & b907;
  assign or907  = a907 | b907;
  assign c908 = (a907 & b907) | (a907 & c907) | (b907 & c907);
  wire c_sub908;
  assign c_sub908 = (a907 & b_inv907) | (a907 & c907) | (b_inv907 & c907);
  wire s908, sub908, and908, or908;
  wire b_inv908;
  assign b_inv908 = ~b908;
  assign s908  = a908 ^ b908 ^ c908;
  assign sub908 = a908 ^ b_inv908 ^ c908;
  assign and908 = a908 & b908;
  assign or908  = a908 | b908;
  assign c909 = (a908 & b908) | (a908 & c908) | (b908 & c908);
  wire c_sub909;
  assign c_sub909 = (a908 & b_inv908) | (a908 & c908) | (b_inv908 & c908);
  wire s909, sub909, and909, or909;
  wire b_inv909;
  assign b_inv909 = ~b909;
  assign s909  = a909 ^ b909 ^ c909;
  assign sub909 = a909 ^ b_inv909 ^ c909;
  assign and909 = a909 & b909;
  assign or909  = a909 | b909;
  assign c910 = (a909 & b909) | (a909 & c909) | (b909 & c909);
  wire c_sub910;
  assign c_sub910 = (a909 & b_inv909) | (a909 & c909) | (b_inv909 & c909);
  wire s910, sub910, and910, or910;
  wire b_inv910;
  assign b_inv910 = ~b910;
  assign s910  = a910 ^ b910 ^ c910;
  assign sub910 = a910 ^ b_inv910 ^ c910;
  assign and910 = a910 & b910;
  assign or910  = a910 | b910;
  assign c911 = (a910 & b910) | (a910 & c910) | (b910 & c910);
  wire c_sub911;
  assign c_sub911 = (a910 & b_inv910) | (a910 & c910) | (b_inv910 & c910);
  wire s911, sub911, and911, or911;
  wire b_inv911;
  assign b_inv911 = ~b911;
  assign s911  = a911 ^ b911 ^ c911;
  assign sub911 = a911 ^ b_inv911 ^ c911;
  assign and911 = a911 & b911;
  assign or911  = a911 | b911;
  assign c912 = (a911 & b911) | (a911 & c911) | (b911 & c911);
  wire c_sub912;
  assign c_sub912 = (a911 & b_inv911) | (a911 & c911) | (b_inv911 & c911);
  wire s912, sub912, and912, or912;
  wire b_inv912;
  assign b_inv912 = ~b912;
  assign s912  = a912 ^ b912 ^ c912;
  assign sub912 = a912 ^ b_inv912 ^ c912;
  assign and912 = a912 & b912;
  assign or912  = a912 | b912;
  assign c913 = (a912 & b912) | (a912 & c912) | (b912 & c912);
  wire c_sub913;
  assign c_sub913 = (a912 & b_inv912) | (a912 & c912) | (b_inv912 & c912);
  wire s913, sub913, and913, or913;
  wire b_inv913;
  assign b_inv913 = ~b913;
  assign s913  = a913 ^ b913 ^ c913;
  assign sub913 = a913 ^ b_inv913 ^ c913;
  assign and913 = a913 & b913;
  assign or913  = a913 | b913;
  assign c914 = (a913 & b913) | (a913 & c913) | (b913 & c913);
  wire c_sub914;
  assign c_sub914 = (a913 & b_inv913) | (a913 & c913) | (b_inv913 & c913);
  wire s914, sub914, and914, or914;
  wire b_inv914;
  assign b_inv914 = ~b914;
  assign s914  = a914 ^ b914 ^ c914;
  assign sub914 = a914 ^ b_inv914 ^ c914;
  assign and914 = a914 & b914;
  assign or914  = a914 | b914;
  assign c915 = (a914 & b914) | (a914 & c914) | (b914 & c914);
  wire c_sub915;
  assign c_sub915 = (a914 & b_inv914) | (a914 & c914) | (b_inv914 & c914);
  wire s915, sub915, and915, or915;
  wire b_inv915;
  assign b_inv915 = ~b915;
  assign s915  = a915 ^ b915 ^ c915;
  assign sub915 = a915 ^ b_inv915 ^ c915;
  assign and915 = a915 & b915;
  assign or915  = a915 | b915;
  assign c916 = (a915 & b915) | (a915 & c915) | (b915 & c915);
  wire c_sub916;
  assign c_sub916 = (a915 & b_inv915) | (a915 & c915) | (b_inv915 & c915);
  wire s916, sub916, and916, or916;
  wire b_inv916;
  assign b_inv916 = ~b916;
  assign s916  = a916 ^ b916 ^ c916;
  assign sub916 = a916 ^ b_inv916 ^ c916;
  assign and916 = a916 & b916;
  assign or916  = a916 | b916;
  assign c917 = (a916 & b916) | (a916 & c916) | (b916 & c916);
  wire c_sub917;
  assign c_sub917 = (a916 & b_inv916) | (a916 & c916) | (b_inv916 & c916);
  wire s917, sub917, and917, or917;
  wire b_inv917;
  assign b_inv917 = ~b917;
  assign s917  = a917 ^ b917 ^ c917;
  assign sub917 = a917 ^ b_inv917 ^ c917;
  assign and917 = a917 & b917;
  assign or917  = a917 | b917;
  assign c918 = (a917 & b917) | (a917 & c917) | (b917 & c917);
  wire c_sub918;
  assign c_sub918 = (a917 & b_inv917) | (a917 & c917) | (b_inv917 & c917);
  wire s918, sub918, and918, or918;
  wire b_inv918;
  assign b_inv918 = ~b918;
  assign s918  = a918 ^ b918 ^ c918;
  assign sub918 = a918 ^ b_inv918 ^ c918;
  assign and918 = a918 & b918;
  assign or918  = a918 | b918;
  assign c919 = (a918 & b918) | (a918 & c918) | (b918 & c918);
  wire c_sub919;
  assign c_sub919 = (a918 & b_inv918) | (a918 & c918) | (b_inv918 & c918);
  wire s919, sub919, and919, or919;
  wire b_inv919;
  assign b_inv919 = ~b919;
  assign s919  = a919 ^ b919 ^ c919;
  assign sub919 = a919 ^ b_inv919 ^ c919;
  assign and919 = a919 & b919;
  assign or919  = a919 | b919;
  assign c920 = (a919 & b919) | (a919 & c919) | (b919 & c919);
  wire c_sub920;
  assign c_sub920 = (a919 & b_inv919) | (a919 & c919) | (b_inv919 & c919);
  wire s920, sub920, and920, or920;
  wire b_inv920;
  assign b_inv920 = ~b920;
  assign s920  = a920 ^ b920 ^ c920;
  assign sub920 = a920 ^ b_inv920 ^ c920;
  assign and920 = a920 & b920;
  assign or920  = a920 | b920;
  assign c921 = (a920 & b920) | (a920 & c920) | (b920 & c920);
  wire c_sub921;
  assign c_sub921 = (a920 & b_inv920) | (a920 & c920) | (b_inv920 & c920);
  wire s921, sub921, and921, or921;
  wire b_inv921;
  assign b_inv921 = ~b921;
  assign s921  = a921 ^ b921 ^ c921;
  assign sub921 = a921 ^ b_inv921 ^ c921;
  assign and921 = a921 & b921;
  assign or921  = a921 | b921;
  assign c922 = (a921 & b921) | (a921 & c921) | (b921 & c921);
  wire c_sub922;
  assign c_sub922 = (a921 & b_inv921) | (a921 & c921) | (b_inv921 & c921);
  wire s922, sub922, and922, or922;
  wire b_inv922;
  assign b_inv922 = ~b922;
  assign s922  = a922 ^ b922 ^ c922;
  assign sub922 = a922 ^ b_inv922 ^ c922;
  assign and922 = a922 & b922;
  assign or922  = a922 | b922;
  assign c923 = (a922 & b922) | (a922 & c922) | (b922 & c922);
  wire c_sub923;
  assign c_sub923 = (a922 & b_inv922) | (a922 & c922) | (b_inv922 & c922);
  wire s923, sub923, and923, or923;
  wire b_inv923;
  assign b_inv923 = ~b923;
  assign s923  = a923 ^ b923 ^ c923;
  assign sub923 = a923 ^ b_inv923 ^ c923;
  assign and923 = a923 & b923;
  assign or923  = a923 | b923;
  assign c924 = (a923 & b923) | (a923 & c923) | (b923 & c923);
  wire c_sub924;
  assign c_sub924 = (a923 & b_inv923) | (a923 & c923) | (b_inv923 & c923);
  wire s924, sub924, and924, or924;
  wire b_inv924;
  assign b_inv924 = ~b924;
  assign s924  = a924 ^ b924 ^ c924;
  assign sub924 = a924 ^ b_inv924 ^ c924;
  assign and924 = a924 & b924;
  assign or924  = a924 | b924;
  assign c925 = (a924 & b924) | (a924 & c924) | (b924 & c924);
  wire c_sub925;
  assign c_sub925 = (a924 & b_inv924) | (a924 & c924) | (b_inv924 & c924);
  wire s925, sub925, and925, or925;
  wire b_inv925;
  assign b_inv925 = ~b925;
  assign s925  = a925 ^ b925 ^ c925;
  assign sub925 = a925 ^ b_inv925 ^ c925;
  assign and925 = a925 & b925;
  assign or925  = a925 | b925;
  assign c926 = (a925 & b925) | (a925 & c925) | (b925 & c925);
  wire c_sub926;
  assign c_sub926 = (a925 & b_inv925) | (a925 & c925) | (b_inv925 & c925);
  wire s926, sub926, and926, or926;
  wire b_inv926;
  assign b_inv926 = ~b926;
  assign s926  = a926 ^ b926 ^ c926;
  assign sub926 = a926 ^ b_inv926 ^ c926;
  assign and926 = a926 & b926;
  assign or926  = a926 | b926;
  assign c927 = (a926 & b926) | (a926 & c926) | (b926 & c926);
  wire c_sub927;
  assign c_sub927 = (a926 & b_inv926) | (a926 & c926) | (b_inv926 & c926);
  wire s927, sub927, and927, or927;
  wire b_inv927;
  assign b_inv927 = ~b927;
  assign s927  = a927 ^ b927 ^ c927;
  assign sub927 = a927 ^ b_inv927 ^ c927;
  assign and927 = a927 & b927;
  assign or927  = a927 | b927;
  assign c928 = (a927 & b927) | (a927 & c927) | (b927 & c927);
  wire c_sub928;
  assign c_sub928 = (a927 & b_inv927) | (a927 & c927) | (b_inv927 & c927);
  wire s928, sub928, and928, or928;
  wire b_inv928;
  assign b_inv928 = ~b928;
  assign s928  = a928 ^ b928 ^ c928;
  assign sub928 = a928 ^ b_inv928 ^ c928;
  assign and928 = a928 & b928;
  assign or928  = a928 | b928;
  assign c929 = (a928 & b928) | (a928 & c928) | (b928 & c928);
  wire c_sub929;
  assign c_sub929 = (a928 & b_inv928) | (a928 & c928) | (b_inv928 & c928);
  wire s929, sub929, and929, or929;
  wire b_inv929;
  assign b_inv929 = ~b929;
  assign s929  = a929 ^ b929 ^ c929;
  assign sub929 = a929 ^ b_inv929 ^ c929;
  assign and929 = a929 & b929;
  assign or929  = a929 | b929;
  assign c930 = (a929 & b929) | (a929 & c929) | (b929 & c929);
  wire c_sub930;
  assign c_sub930 = (a929 & b_inv929) | (a929 & c929) | (b_inv929 & c929);
  wire s930, sub930, and930, or930;
  wire b_inv930;
  assign b_inv930 = ~b930;
  assign s930  = a930 ^ b930 ^ c930;
  assign sub930 = a930 ^ b_inv930 ^ c930;
  assign and930 = a930 & b930;
  assign or930  = a930 | b930;
  assign c931 = (a930 & b930) | (a930 & c930) | (b930 & c930);
  wire c_sub931;
  assign c_sub931 = (a930 & b_inv930) | (a930 & c930) | (b_inv930 & c930);
  wire s931, sub931, and931, or931;
  wire b_inv931;
  assign b_inv931 = ~b931;
  assign s931  = a931 ^ b931 ^ c931;
  assign sub931 = a931 ^ b_inv931 ^ c931;
  assign and931 = a931 & b931;
  assign or931  = a931 | b931;
  assign c932 = (a931 & b931) | (a931 & c931) | (b931 & c931);
  wire c_sub932;
  assign c_sub932 = (a931 & b_inv931) | (a931 & c931) | (b_inv931 & c931);
  wire s932, sub932, and932, or932;
  wire b_inv932;
  assign b_inv932 = ~b932;
  assign s932  = a932 ^ b932 ^ c932;
  assign sub932 = a932 ^ b_inv932 ^ c932;
  assign and932 = a932 & b932;
  assign or932  = a932 | b932;
  assign c933 = (a932 & b932) | (a932 & c932) | (b932 & c932);
  wire c_sub933;
  assign c_sub933 = (a932 & b_inv932) | (a932 & c932) | (b_inv932 & c932);
  wire s933, sub933, and933, or933;
  wire b_inv933;
  assign b_inv933 = ~b933;
  assign s933  = a933 ^ b933 ^ c933;
  assign sub933 = a933 ^ b_inv933 ^ c933;
  assign and933 = a933 & b933;
  assign or933  = a933 | b933;
  assign c934 = (a933 & b933) | (a933 & c933) | (b933 & c933);
  wire c_sub934;
  assign c_sub934 = (a933 & b_inv933) | (a933 & c933) | (b_inv933 & c933);
  wire s934, sub934, and934, or934;
  wire b_inv934;
  assign b_inv934 = ~b934;
  assign s934  = a934 ^ b934 ^ c934;
  assign sub934 = a934 ^ b_inv934 ^ c934;
  assign and934 = a934 & b934;
  assign or934  = a934 | b934;
  assign c935 = (a934 & b934) | (a934 & c934) | (b934 & c934);
  wire c_sub935;
  assign c_sub935 = (a934 & b_inv934) | (a934 & c934) | (b_inv934 & c934);
  wire s935, sub935, and935, or935;
  wire b_inv935;
  assign b_inv935 = ~b935;
  assign s935  = a935 ^ b935 ^ c935;
  assign sub935 = a935 ^ b_inv935 ^ c935;
  assign and935 = a935 & b935;
  assign or935  = a935 | b935;
  assign c936 = (a935 & b935) | (a935 & c935) | (b935 & c935);
  wire c_sub936;
  assign c_sub936 = (a935 & b_inv935) | (a935 & c935) | (b_inv935 & c935);
  wire s936, sub936, and936, or936;
  wire b_inv936;
  assign b_inv936 = ~b936;
  assign s936  = a936 ^ b936 ^ c936;
  assign sub936 = a936 ^ b_inv936 ^ c936;
  assign and936 = a936 & b936;
  assign or936  = a936 | b936;
  assign c937 = (a936 & b936) | (a936 & c936) | (b936 & c936);
  wire c_sub937;
  assign c_sub937 = (a936 & b_inv936) | (a936 & c936) | (b_inv936 & c936);
  wire s937, sub937, and937, or937;
  wire b_inv937;
  assign b_inv937 = ~b937;
  assign s937  = a937 ^ b937 ^ c937;
  assign sub937 = a937 ^ b_inv937 ^ c937;
  assign and937 = a937 & b937;
  assign or937  = a937 | b937;
  assign c938 = (a937 & b937) | (a937 & c937) | (b937 & c937);
  wire c_sub938;
  assign c_sub938 = (a937 & b_inv937) | (a937 & c937) | (b_inv937 & c937);
  wire s938, sub938, and938, or938;
  wire b_inv938;
  assign b_inv938 = ~b938;
  assign s938  = a938 ^ b938 ^ c938;
  assign sub938 = a938 ^ b_inv938 ^ c938;
  assign and938 = a938 & b938;
  assign or938  = a938 | b938;
  assign c939 = (a938 & b938) | (a938 & c938) | (b938 & c938);
  wire c_sub939;
  assign c_sub939 = (a938 & b_inv938) | (a938 & c938) | (b_inv938 & c938);
  wire s939, sub939, and939, or939;
  wire b_inv939;
  assign b_inv939 = ~b939;
  assign s939  = a939 ^ b939 ^ c939;
  assign sub939 = a939 ^ b_inv939 ^ c939;
  assign and939 = a939 & b939;
  assign or939  = a939 | b939;
  assign c940 = (a939 & b939) | (a939 & c939) | (b939 & c939);
  wire c_sub940;
  assign c_sub940 = (a939 & b_inv939) | (a939 & c939) | (b_inv939 & c939);
  wire s940, sub940, and940, or940;
  wire b_inv940;
  assign b_inv940 = ~b940;
  assign s940  = a940 ^ b940 ^ c940;
  assign sub940 = a940 ^ b_inv940 ^ c940;
  assign and940 = a940 & b940;
  assign or940  = a940 | b940;
  assign c941 = (a940 & b940) | (a940 & c940) | (b940 & c940);
  wire c_sub941;
  assign c_sub941 = (a940 & b_inv940) | (a940 & c940) | (b_inv940 & c940);
  wire s941, sub941, and941, or941;
  wire b_inv941;
  assign b_inv941 = ~b941;
  assign s941  = a941 ^ b941 ^ c941;
  assign sub941 = a941 ^ b_inv941 ^ c941;
  assign and941 = a941 & b941;
  assign or941  = a941 | b941;
  assign c942 = (a941 & b941) | (a941 & c941) | (b941 & c941);
  wire c_sub942;
  assign c_sub942 = (a941 & b_inv941) | (a941 & c941) | (b_inv941 & c941);
  wire s942, sub942, and942, or942;
  wire b_inv942;
  assign b_inv942 = ~b942;
  assign s942  = a942 ^ b942 ^ c942;
  assign sub942 = a942 ^ b_inv942 ^ c942;
  assign and942 = a942 & b942;
  assign or942  = a942 | b942;
  assign c943 = (a942 & b942) | (a942 & c942) | (b942 & c942);
  wire c_sub943;
  assign c_sub943 = (a942 & b_inv942) | (a942 & c942) | (b_inv942 & c942);
  wire s943, sub943, and943, or943;
  wire b_inv943;
  assign b_inv943 = ~b943;
  assign s943  = a943 ^ b943 ^ c943;
  assign sub943 = a943 ^ b_inv943 ^ c943;
  assign and943 = a943 & b943;
  assign or943  = a943 | b943;
  assign c944 = (a943 & b943) | (a943 & c943) | (b943 & c943);
  wire c_sub944;
  assign c_sub944 = (a943 & b_inv943) | (a943 & c943) | (b_inv943 & c943);
  wire s944, sub944, and944, or944;
  wire b_inv944;
  assign b_inv944 = ~b944;
  assign s944  = a944 ^ b944 ^ c944;
  assign sub944 = a944 ^ b_inv944 ^ c944;
  assign and944 = a944 & b944;
  assign or944  = a944 | b944;
  assign c945 = (a944 & b944) | (a944 & c944) | (b944 & c944);
  wire c_sub945;
  assign c_sub945 = (a944 & b_inv944) | (a944 & c944) | (b_inv944 & c944);
  wire s945, sub945, and945, or945;
  wire b_inv945;
  assign b_inv945 = ~b945;
  assign s945  = a945 ^ b945 ^ c945;
  assign sub945 = a945 ^ b_inv945 ^ c945;
  assign and945 = a945 & b945;
  assign or945  = a945 | b945;
  assign c946 = (a945 & b945) | (a945 & c945) | (b945 & c945);
  wire c_sub946;
  assign c_sub946 = (a945 & b_inv945) | (a945 & c945) | (b_inv945 & c945);
  wire s946, sub946, and946, or946;
  wire b_inv946;
  assign b_inv946 = ~b946;
  assign s946  = a946 ^ b946 ^ c946;
  assign sub946 = a946 ^ b_inv946 ^ c946;
  assign and946 = a946 & b946;
  assign or946  = a946 | b946;
  assign c947 = (a946 & b946) | (a946 & c946) | (b946 & c946);
  wire c_sub947;
  assign c_sub947 = (a946 & b_inv946) | (a946 & c946) | (b_inv946 & c946);
  wire s947, sub947, and947, or947;
  wire b_inv947;
  assign b_inv947 = ~b947;
  assign s947  = a947 ^ b947 ^ c947;
  assign sub947 = a947 ^ b_inv947 ^ c947;
  assign and947 = a947 & b947;
  assign or947  = a947 | b947;
  assign c948 = (a947 & b947) | (a947 & c947) | (b947 & c947);
  wire c_sub948;
  assign c_sub948 = (a947 & b_inv947) | (a947 & c947) | (b_inv947 & c947);
  wire s948, sub948, and948, or948;
  wire b_inv948;
  assign b_inv948 = ~b948;
  assign s948  = a948 ^ b948 ^ c948;
  assign sub948 = a948 ^ b_inv948 ^ c948;
  assign and948 = a948 & b948;
  assign or948  = a948 | b948;
  assign c949 = (a948 & b948) | (a948 & c948) | (b948 & c948);
  wire c_sub949;
  assign c_sub949 = (a948 & b_inv948) | (a948 & c948) | (b_inv948 & c948);
  wire s949, sub949, and949, or949;
  wire b_inv949;
  assign b_inv949 = ~b949;
  assign s949  = a949 ^ b949 ^ c949;
  assign sub949 = a949 ^ b_inv949 ^ c949;
  assign and949 = a949 & b949;
  assign or949  = a949 | b949;
  assign c950 = (a949 & b949) | (a949 & c949) | (b949 & c949);
  wire c_sub950;
  assign c_sub950 = (a949 & b_inv949) | (a949 & c949) | (b_inv949 & c949);
  wire s950, sub950, and950, or950;
  wire b_inv950;
  assign b_inv950 = ~b950;
  assign s950  = a950 ^ b950 ^ c950;
  assign sub950 = a950 ^ b_inv950 ^ c950;
  assign and950 = a950 & b950;
  assign or950  = a950 | b950;
  assign c951 = (a950 & b950) | (a950 & c950) | (b950 & c950);
  wire c_sub951;
  assign c_sub951 = (a950 & b_inv950) | (a950 & c950) | (b_inv950 & c950);
  wire s951, sub951, and951, or951;
  wire b_inv951;
  assign b_inv951 = ~b951;
  assign s951  = a951 ^ b951 ^ c951;
  assign sub951 = a951 ^ b_inv951 ^ c951;
  assign and951 = a951 & b951;
  assign or951  = a951 | b951;
  assign c952 = (a951 & b951) | (a951 & c951) | (b951 & c951);
  wire c_sub952;
  assign c_sub952 = (a951 & b_inv951) | (a951 & c951) | (b_inv951 & c951);
  wire s952, sub952, and952, or952;
  wire b_inv952;
  assign b_inv952 = ~b952;
  assign s952  = a952 ^ b952 ^ c952;
  assign sub952 = a952 ^ b_inv952 ^ c952;
  assign and952 = a952 & b952;
  assign or952  = a952 | b952;
  assign c953 = (a952 & b952) | (a952 & c952) | (b952 & c952);
  wire c_sub953;
  assign c_sub953 = (a952 & b_inv952) | (a952 & c952) | (b_inv952 & c952);
  wire s953, sub953, and953, or953;
  wire b_inv953;
  assign b_inv953 = ~b953;
  assign s953  = a953 ^ b953 ^ c953;
  assign sub953 = a953 ^ b_inv953 ^ c953;
  assign and953 = a953 & b953;
  assign or953  = a953 | b953;
  assign c954 = (a953 & b953) | (a953 & c953) | (b953 & c953);
  wire c_sub954;
  assign c_sub954 = (a953 & b_inv953) | (a953 & c953) | (b_inv953 & c953);
  wire s954, sub954, and954, or954;
  wire b_inv954;
  assign b_inv954 = ~b954;
  assign s954  = a954 ^ b954 ^ c954;
  assign sub954 = a954 ^ b_inv954 ^ c954;
  assign and954 = a954 & b954;
  assign or954  = a954 | b954;
  assign c955 = (a954 & b954) | (a954 & c954) | (b954 & c954);
  wire c_sub955;
  assign c_sub955 = (a954 & b_inv954) | (a954 & c954) | (b_inv954 & c954);
  wire s955, sub955, and955, or955;
  wire b_inv955;
  assign b_inv955 = ~b955;
  assign s955  = a955 ^ b955 ^ c955;
  assign sub955 = a955 ^ b_inv955 ^ c955;
  assign and955 = a955 & b955;
  assign or955  = a955 | b955;
  assign c956 = (a955 & b955) | (a955 & c955) | (b955 & c955);
  wire c_sub956;
  assign c_sub956 = (a955 & b_inv955) | (a955 & c955) | (b_inv955 & c955);
  wire s956, sub956, and956, or956;
  wire b_inv956;
  assign b_inv956 = ~b956;
  assign s956  = a956 ^ b956 ^ c956;
  assign sub956 = a956 ^ b_inv956 ^ c956;
  assign and956 = a956 & b956;
  assign or956  = a956 | b956;
  assign c957 = (a956 & b956) | (a956 & c956) | (b956 & c956);
  wire c_sub957;
  assign c_sub957 = (a956 & b_inv956) | (a956 & c956) | (b_inv956 & c956);
  wire s957, sub957, and957, or957;
  wire b_inv957;
  assign b_inv957 = ~b957;
  assign s957  = a957 ^ b957 ^ c957;
  assign sub957 = a957 ^ b_inv957 ^ c957;
  assign and957 = a957 & b957;
  assign or957  = a957 | b957;
  assign c958 = (a957 & b957) | (a957 & c957) | (b957 & c957);
  wire c_sub958;
  assign c_sub958 = (a957 & b_inv957) | (a957 & c957) | (b_inv957 & c957);
  wire s958, sub958, and958, or958;
  wire b_inv958;
  assign b_inv958 = ~b958;
  assign s958  = a958 ^ b958 ^ c958;
  assign sub958 = a958 ^ b_inv958 ^ c958;
  assign and958 = a958 & b958;
  assign or958  = a958 | b958;
  assign c959 = (a958 & b958) | (a958 & c958) | (b958 & c958);
  wire c_sub959;
  assign c_sub959 = (a958 & b_inv958) | (a958 & c958) | (b_inv958 & c958);
  wire s959, sub959, and959, or959;
  wire b_inv959;
  assign b_inv959 = ~b959;
  assign s959  = a959 ^ b959 ^ c959;
  assign sub959 = a959 ^ b_inv959 ^ c959;
  assign and959 = a959 & b959;
  assign or959  = a959 | b959;
  assign c960 = (a959 & b959) | (a959 & c959) | (b959 & c959);
  wire c_sub960;
  assign c_sub960 = (a959 & b_inv959) | (a959 & c959) | (b_inv959 & c959);
  wire s960, sub960, and960, or960;
  wire b_inv960;
  assign b_inv960 = ~b960;
  assign s960  = a960 ^ b960 ^ c960;
  assign sub960 = a960 ^ b_inv960 ^ c960;
  assign and960 = a960 & b960;
  assign or960  = a960 | b960;
  assign c961 = (a960 & b960) | (a960 & c960) | (b960 & c960);
  wire c_sub961;
  assign c_sub961 = (a960 & b_inv960) | (a960 & c960) | (b_inv960 & c960);
  wire s961, sub961, and961, or961;
  wire b_inv961;
  assign b_inv961 = ~b961;
  assign s961  = a961 ^ b961 ^ c961;
  assign sub961 = a961 ^ b_inv961 ^ c961;
  assign and961 = a961 & b961;
  assign or961  = a961 | b961;
  assign c962 = (a961 & b961) | (a961 & c961) | (b961 & c961);
  wire c_sub962;
  assign c_sub962 = (a961 & b_inv961) | (a961 & c961) | (b_inv961 & c961);
  wire s962, sub962, and962, or962;
  wire b_inv962;
  assign b_inv962 = ~b962;
  assign s962  = a962 ^ b962 ^ c962;
  assign sub962 = a962 ^ b_inv962 ^ c962;
  assign and962 = a962 & b962;
  assign or962  = a962 | b962;
  assign c963 = (a962 & b962) | (a962 & c962) | (b962 & c962);
  wire c_sub963;
  assign c_sub963 = (a962 & b_inv962) | (a962 & c962) | (b_inv962 & c962);
  wire s963, sub963, and963, or963;
  wire b_inv963;
  assign b_inv963 = ~b963;
  assign s963  = a963 ^ b963 ^ c963;
  assign sub963 = a963 ^ b_inv963 ^ c963;
  assign and963 = a963 & b963;
  assign or963  = a963 | b963;
  assign c964 = (a963 & b963) | (a963 & c963) | (b963 & c963);
  wire c_sub964;
  assign c_sub964 = (a963 & b_inv963) | (a963 & c963) | (b_inv963 & c963);
  wire s964, sub964, and964, or964;
  wire b_inv964;
  assign b_inv964 = ~b964;
  assign s964  = a964 ^ b964 ^ c964;
  assign sub964 = a964 ^ b_inv964 ^ c964;
  assign and964 = a964 & b964;
  assign or964  = a964 | b964;
  assign c965 = (a964 & b964) | (a964 & c964) | (b964 & c964);
  wire c_sub965;
  assign c_sub965 = (a964 & b_inv964) | (a964 & c964) | (b_inv964 & c964);
  wire s965, sub965, and965, or965;
  wire b_inv965;
  assign b_inv965 = ~b965;
  assign s965  = a965 ^ b965 ^ c965;
  assign sub965 = a965 ^ b_inv965 ^ c965;
  assign and965 = a965 & b965;
  assign or965  = a965 | b965;
  assign c966 = (a965 & b965) | (a965 & c965) | (b965 & c965);
  wire c_sub966;
  assign c_sub966 = (a965 & b_inv965) | (a965 & c965) | (b_inv965 & c965);
  wire s966, sub966, and966, or966;
  wire b_inv966;
  assign b_inv966 = ~b966;
  assign s966  = a966 ^ b966 ^ c966;
  assign sub966 = a966 ^ b_inv966 ^ c966;
  assign and966 = a966 & b966;
  assign or966  = a966 | b966;
  assign c967 = (a966 & b966) | (a966 & c966) | (b966 & c966);
  wire c_sub967;
  assign c_sub967 = (a966 & b_inv966) | (a966 & c966) | (b_inv966 & c966);
  wire s967, sub967, and967, or967;
  wire b_inv967;
  assign b_inv967 = ~b967;
  assign s967  = a967 ^ b967 ^ c967;
  assign sub967 = a967 ^ b_inv967 ^ c967;
  assign and967 = a967 & b967;
  assign or967  = a967 | b967;
  assign c968 = (a967 & b967) | (a967 & c967) | (b967 & c967);
  wire c_sub968;
  assign c_sub968 = (a967 & b_inv967) | (a967 & c967) | (b_inv967 & c967);
  wire s968, sub968, and968, or968;
  wire b_inv968;
  assign b_inv968 = ~b968;
  assign s968  = a968 ^ b968 ^ c968;
  assign sub968 = a968 ^ b_inv968 ^ c968;
  assign and968 = a968 & b968;
  assign or968  = a968 | b968;
  assign c969 = (a968 & b968) | (a968 & c968) | (b968 & c968);
  wire c_sub969;
  assign c_sub969 = (a968 & b_inv968) | (a968 & c968) | (b_inv968 & c968);
  wire s969, sub969, and969, or969;
  wire b_inv969;
  assign b_inv969 = ~b969;
  assign s969  = a969 ^ b969 ^ c969;
  assign sub969 = a969 ^ b_inv969 ^ c969;
  assign and969 = a969 & b969;
  assign or969  = a969 | b969;
  assign c970 = (a969 & b969) | (a969 & c969) | (b969 & c969);
  wire c_sub970;
  assign c_sub970 = (a969 & b_inv969) | (a969 & c969) | (b_inv969 & c969);
  wire s970, sub970, and970, or970;
  wire b_inv970;
  assign b_inv970 = ~b970;
  assign s970  = a970 ^ b970 ^ c970;
  assign sub970 = a970 ^ b_inv970 ^ c970;
  assign and970 = a970 & b970;
  assign or970  = a970 | b970;
  assign c971 = (a970 & b970) | (a970 & c970) | (b970 & c970);
  wire c_sub971;
  assign c_sub971 = (a970 & b_inv970) | (a970 & c970) | (b_inv970 & c970);
  wire s971, sub971, and971, or971;
  wire b_inv971;
  assign b_inv971 = ~b971;
  assign s971  = a971 ^ b971 ^ c971;
  assign sub971 = a971 ^ b_inv971 ^ c971;
  assign and971 = a971 & b971;
  assign or971  = a971 | b971;
  assign c972 = (a971 & b971) | (a971 & c971) | (b971 & c971);
  wire c_sub972;
  assign c_sub972 = (a971 & b_inv971) | (a971 & c971) | (b_inv971 & c971);
  wire s972, sub972, and972, or972;
  wire b_inv972;
  assign b_inv972 = ~b972;
  assign s972  = a972 ^ b972 ^ c972;
  assign sub972 = a972 ^ b_inv972 ^ c972;
  assign and972 = a972 & b972;
  assign or972  = a972 | b972;
  assign c973 = (a972 & b972) | (a972 & c972) | (b972 & c972);
  wire c_sub973;
  assign c_sub973 = (a972 & b_inv972) | (a972 & c972) | (b_inv972 & c972);
  wire s973, sub973, and973, or973;
  wire b_inv973;
  assign b_inv973 = ~b973;
  assign s973  = a973 ^ b973 ^ c973;
  assign sub973 = a973 ^ b_inv973 ^ c973;
  assign and973 = a973 & b973;
  assign or973  = a973 | b973;
  assign c974 = (a973 & b973) | (a973 & c973) | (b973 & c973);
  wire c_sub974;
  assign c_sub974 = (a973 & b_inv973) | (a973 & c973) | (b_inv973 & c973);
  wire s974, sub974, and974, or974;
  wire b_inv974;
  assign b_inv974 = ~b974;
  assign s974  = a974 ^ b974 ^ c974;
  assign sub974 = a974 ^ b_inv974 ^ c974;
  assign and974 = a974 & b974;
  assign or974  = a974 | b974;
  assign c975 = (a974 & b974) | (a974 & c974) | (b974 & c974);
  wire c_sub975;
  assign c_sub975 = (a974 & b_inv974) | (a974 & c974) | (b_inv974 & c974);
  wire s975, sub975, and975, or975;
  wire b_inv975;
  assign b_inv975 = ~b975;
  assign s975  = a975 ^ b975 ^ c975;
  assign sub975 = a975 ^ b_inv975 ^ c975;
  assign and975 = a975 & b975;
  assign or975  = a975 | b975;
  assign c976 = (a975 & b975) | (a975 & c975) | (b975 & c975);
  wire c_sub976;
  assign c_sub976 = (a975 & b_inv975) | (a975 & c975) | (b_inv975 & c975);
  wire s976, sub976, and976, or976;
  wire b_inv976;
  assign b_inv976 = ~b976;
  assign s976  = a976 ^ b976 ^ c976;
  assign sub976 = a976 ^ b_inv976 ^ c976;
  assign and976 = a976 & b976;
  assign or976  = a976 | b976;
  assign c977 = (a976 & b976) | (a976 & c976) | (b976 & c976);
  wire c_sub977;
  assign c_sub977 = (a976 & b_inv976) | (a976 & c976) | (b_inv976 & c976);
  wire s977, sub977, and977, or977;
  wire b_inv977;
  assign b_inv977 = ~b977;
  assign s977  = a977 ^ b977 ^ c977;
  assign sub977 = a977 ^ b_inv977 ^ c977;
  assign and977 = a977 & b977;
  assign or977  = a977 | b977;
  assign c978 = (a977 & b977) | (a977 & c977) | (b977 & c977);
  wire c_sub978;
  assign c_sub978 = (a977 & b_inv977) | (a977 & c977) | (b_inv977 & c977);
  wire s978, sub978, and978, or978;
  wire b_inv978;
  assign b_inv978 = ~b978;
  assign s978  = a978 ^ b978 ^ c978;
  assign sub978 = a978 ^ b_inv978 ^ c978;
  assign and978 = a978 & b978;
  assign or978  = a978 | b978;
  assign c979 = (a978 & b978) | (a978 & c978) | (b978 & c978);
  wire c_sub979;
  assign c_sub979 = (a978 & b_inv978) | (a978 & c978) | (b_inv978 & c978);
  wire s979, sub979, and979, or979;
  wire b_inv979;
  assign b_inv979 = ~b979;
  assign s979  = a979 ^ b979 ^ c979;
  assign sub979 = a979 ^ b_inv979 ^ c979;
  assign and979 = a979 & b979;
  assign or979  = a979 | b979;
  assign c980 = (a979 & b979) | (a979 & c979) | (b979 & c979);
  wire c_sub980;
  assign c_sub980 = (a979 & b_inv979) | (a979 & c979) | (b_inv979 & c979);
  wire s980, sub980, and980, or980;
  wire b_inv980;
  assign b_inv980 = ~b980;
  assign s980  = a980 ^ b980 ^ c980;
  assign sub980 = a980 ^ b_inv980 ^ c980;
  assign and980 = a980 & b980;
  assign or980  = a980 | b980;
  assign c981 = (a980 & b980) | (a980 & c980) | (b980 & c980);
  wire c_sub981;
  assign c_sub981 = (a980 & b_inv980) | (a980 & c980) | (b_inv980 & c980);
  wire s981, sub981, and981, or981;
  wire b_inv981;
  assign b_inv981 = ~b981;
  assign s981  = a981 ^ b981 ^ c981;
  assign sub981 = a981 ^ b_inv981 ^ c981;
  assign and981 = a981 & b981;
  assign or981  = a981 | b981;
  assign c982 = (a981 & b981) | (a981 & c981) | (b981 & c981);
  wire c_sub982;
  assign c_sub982 = (a981 & b_inv981) | (a981 & c981) | (b_inv981 & c981);
  wire s982, sub982, and982, or982;
  wire b_inv982;
  assign b_inv982 = ~b982;
  assign s982  = a982 ^ b982 ^ c982;
  assign sub982 = a982 ^ b_inv982 ^ c982;
  assign and982 = a982 & b982;
  assign or982  = a982 | b982;
  assign c983 = (a982 & b982) | (a982 & c982) | (b982 & c982);
  wire c_sub983;
  assign c_sub983 = (a982 & b_inv982) | (a982 & c982) | (b_inv982 & c982);
  wire s983, sub983, and983, or983;
  wire b_inv983;
  assign b_inv983 = ~b983;
  assign s983  = a983 ^ b983 ^ c983;
  assign sub983 = a983 ^ b_inv983 ^ c983;
  assign and983 = a983 & b983;
  assign or983  = a983 | b983;
  assign c984 = (a983 & b983) | (a983 & c983) | (b983 & c983);
  wire c_sub984;
  assign c_sub984 = (a983 & b_inv983) | (a983 & c983) | (b_inv983 & c983);
  wire s984, sub984, and984, or984;
  wire b_inv984;
  assign b_inv984 = ~b984;
  assign s984  = a984 ^ b984 ^ c984;
  assign sub984 = a984 ^ b_inv984 ^ c984;
  assign and984 = a984 & b984;
  assign or984  = a984 | b984;
  assign c985 = (a984 & b984) | (a984 & c984) | (b984 & c984);
  wire c_sub985;
  assign c_sub985 = (a984 & b_inv984) | (a984 & c984) | (b_inv984 & c984);
  wire s985, sub985, and985, or985;
  wire b_inv985;
  assign b_inv985 = ~b985;
  assign s985  = a985 ^ b985 ^ c985;
  assign sub985 = a985 ^ b_inv985 ^ c985;
  assign and985 = a985 & b985;
  assign or985  = a985 | b985;
  assign c986 = (a985 & b985) | (a985 & c985) | (b985 & c985);
  wire c_sub986;
  assign c_sub986 = (a985 & b_inv985) | (a985 & c985) | (b_inv985 & c985);
  wire s986, sub986, and986, or986;
  wire b_inv986;
  assign b_inv986 = ~b986;
  assign s986  = a986 ^ b986 ^ c986;
  assign sub986 = a986 ^ b_inv986 ^ c986;
  assign and986 = a986 & b986;
  assign or986  = a986 | b986;
  assign c987 = (a986 & b986) | (a986 & c986) | (b986 & c986);
  wire c_sub987;
  assign c_sub987 = (a986 & b_inv986) | (a986 & c986) | (b_inv986 & c986);
  wire s987, sub987, and987, or987;
  wire b_inv987;
  assign b_inv987 = ~b987;
  assign s987  = a987 ^ b987 ^ c987;
  assign sub987 = a987 ^ b_inv987 ^ c987;
  assign and987 = a987 & b987;
  assign or987  = a987 | b987;
  assign c988 = (a987 & b987) | (a987 & c987) | (b987 & c987);
  wire c_sub988;
  assign c_sub988 = (a987 & b_inv987) | (a987 & c987) | (b_inv987 & c987);
  wire s988, sub988, and988, or988;
  wire b_inv988;
  assign b_inv988 = ~b988;
  assign s988  = a988 ^ b988 ^ c988;
  assign sub988 = a988 ^ b_inv988 ^ c988;
  assign and988 = a988 & b988;
  assign or988  = a988 | b988;
  assign c989 = (a988 & b988) | (a988 & c988) | (b988 & c988);
  wire c_sub989;
  assign c_sub989 = (a988 & b_inv988) | (a988 & c988) | (b_inv988 & c988);
  wire s989, sub989, and989, or989;
  wire b_inv989;
  assign b_inv989 = ~b989;
  assign s989  = a989 ^ b989 ^ c989;
  assign sub989 = a989 ^ b_inv989 ^ c989;
  assign and989 = a989 & b989;
  assign or989  = a989 | b989;
  assign c990 = (a989 & b989) | (a989 & c989) | (b989 & c989);
  wire c_sub990;
  assign c_sub990 = (a989 & b_inv989) | (a989 & c989) | (b_inv989 & c989);
  wire s990, sub990, and990, or990;
  wire b_inv990;
  assign b_inv990 = ~b990;
  assign s990  = a990 ^ b990 ^ c990;
  assign sub990 = a990 ^ b_inv990 ^ c990;
  assign and990 = a990 & b990;
  assign or990  = a990 | b990;
  assign c991 = (a990 & b990) | (a990 & c990) | (b990 & c990);
  wire c_sub991;
  assign c_sub991 = (a990 & b_inv990) | (a990 & c990) | (b_inv990 & c990);
  wire s991, sub991, and991, or991;
  wire b_inv991;
  assign b_inv991 = ~b991;
  assign s991  = a991 ^ b991 ^ c991;
  assign sub991 = a991 ^ b_inv991 ^ c991;
  assign and991 = a991 & b991;
  assign or991  = a991 | b991;
  assign c992 = (a991 & b991) | (a991 & c991) | (b991 & c991);
  wire c_sub992;
  assign c_sub992 = (a991 & b_inv991) | (a991 & c991) | (b_inv991 & c991);
  wire s992, sub992, and992, or992;
  wire b_inv992;
  assign b_inv992 = ~b992;
  assign s992  = a992 ^ b992 ^ c992;
  assign sub992 = a992 ^ b_inv992 ^ c992;
  assign and992 = a992 & b992;
  assign or992  = a992 | b992;
  assign c993 = (a992 & b992) | (a992 & c992) | (b992 & c992);
  wire c_sub993;
  assign c_sub993 = (a992 & b_inv992) | (a992 & c992) | (b_inv992 & c992);
  wire s993, sub993, and993, or993;
  wire b_inv993;
  assign b_inv993 = ~b993;
  assign s993  = a993 ^ b993 ^ c993;
  assign sub993 = a993 ^ b_inv993 ^ c993;
  assign and993 = a993 & b993;
  assign or993  = a993 | b993;
  assign c994 = (a993 & b993) | (a993 & c993) | (b993 & c993);
  wire c_sub994;
  assign c_sub994 = (a993 & b_inv993) | (a993 & c993) | (b_inv993 & c993);
  wire s994, sub994, and994, or994;
  wire b_inv994;
  assign b_inv994 = ~b994;
  assign s994  = a994 ^ b994 ^ c994;
  assign sub994 = a994 ^ b_inv994 ^ c994;
  assign and994 = a994 & b994;
  assign or994  = a994 | b994;
  assign c995 = (a994 & b994) | (a994 & c994) | (b994 & c994);
  wire c_sub995;
  assign c_sub995 = (a994 & b_inv994) | (a994 & c994) | (b_inv994 & c994);
  wire s995, sub995, and995, or995;
  wire b_inv995;
  assign b_inv995 = ~b995;
  assign s995  = a995 ^ b995 ^ c995;
  assign sub995 = a995 ^ b_inv995 ^ c995;
  assign and995 = a995 & b995;
  assign or995  = a995 | b995;
  assign c996 = (a995 & b995) | (a995 & c995) | (b995 & c995);
  wire c_sub996;
  assign c_sub996 = (a995 & b_inv995) | (a995 & c995) | (b_inv995 & c995);
  wire s996, sub996, and996, or996;
  wire b_inv996;
  assign b_inv996 = ~b996;
  assign s996  = a996 ^ b996 ^ c996;
  assign sub996 = a996 ^ b_inv996 ^ c996;
  assign and996 = a996 & b996;
  assign or996  = a996 | b996;
  assign c997 = (a996 & b996) | (a996 & c996) | (b996 & c996);
  wire c_sub997;
  assign c_sub997 = (a996 & b_inv996) | (a996 & c996) | (b_inv996 & c996);
  wire s997, sub997, and997, or997;
  wire b_inv997;
  assign b_inv997 = ~b997;
  assign s997  = a997 ^ b997 ^ c997;
  assign sub997 = a997 ^ b_inv997 ^ c997;
  assign and997 = a997 & b997;
  assign or997  = a997 | b997;
  assign c998 = (a997 & b997) | (a997 & c997) | (b997 & c997);
  wire c_sub998;
  assign c_sub998 = (a997 & b_inv997) | (a997 & c997) | (b_inv997 & c997);
  wire s998, sub998, and998, or998;
  wire b_inv998;
  assign b_inv998 = ~b998;
  assign s998  = a998 ^ b998 ^ c998;
  assign sub998 = a998 ^ b_inv998 ^ c998;
  assign and998 = a998 & b998;
  assign or998  = a998 | b998;
  assign c999 = (a998 & b998) | (a998 & c998) | (b998 & c998);
  wire c_sub999;
  assign c_sub999 = (a998 & b_inv998) | (a998 & c998) | (b_inv998 & c998);
  wire s999, sub999, and999, or999;
  wire b_inv999;
  assign b_inv999 = ~b999;
  assign s999  = a999 ^ b999 ^ c999;
  assign sub999 = a999 ^ b_inv999 ^ c999;
  assign and999 = a999 & b999;
  assign or999  = a999 | b999;
  assign c1000 = (a999 & b999) | (a999 & c999) | (b999 & c999);
  wire c_sub1000;
  assign c_sub1000 = (a999 & b_inv999) | (a999 & c999) | (b_inv999 & c999);
  wire s1000, sub1000, and1000, or1000;
  wire b_inv1000;
  assign b_inv1000 = ~b1000;
  assign s1000  = a1000 ^ b1000 ^ c1000;
  assign sub1000 = a1000 ^ b_inv1000 ^ c1000;
  assign and1000 = a1000 & b1000;
  assign or1000  = a1000 | b1000;
  assign c1001 = (a1000 & b1000) | (a1000 & c1000) | (b1000 & c1000);
  wire c_sub1001;
  assign c_sub1001 = (a1000 & b_inv1000) | (a1000 & c1000) | (b_inv1000 & c1000);
  wire s1001, sub1001, and1001, or1001;
  wire b_inv1001;
  assign b_inv1001 = ~b1001;
  assign s1001  = a1001 ^ b1001 ^ c1001;
  assign sub1001 = a1001 ^ b_inv1001 ^ c1001;
  assign and1001 = a1001 & b1001;
  assign or1001  = a1001 | b1001;
  assign c1002 = (a1001 & b1001) | (a1001 & c1001) | (b1001 & c1001);
  wire c_sub1002;
  assign c_sub1002 = (a1001 & b_inv1001) | (a1001 & c1001) | (b_inv1001 & c1001);
  wire s1002, sub1002, and1002, or1002;
  wire b_inv1002;
  assign b_inv1002 = ~b1002;
  assign s1002  = a1002 ^ b1002 ^ c1002;
  assign sub1002 = a1002 ^ b_inv1002 ^ c1002;
  assign and1002 = a1002 & b1002;
  assign or1002  = a1002 | b1002;
  assign c1003 = (a1002 & b1002) | (a1002 & c1002) | (b1002 & c1002);
  wire c_sub1003;
  assign c_sub1003 = (a1002 & b_inv1002) | (a1002 & c1002) | (b_inv1002 & c1002);
  wire s1003, sub1003, and1003, or1003;
  wire b_inv1003;
  assign b_inv1003 = ~b1003;
  assign s1003  = a1003 ^ b1003 ^ c1003;
  assign sub1003 = a1003 ^ b_inv1003 ^ c1003;
  assign and1003 = a1003 & b1003;
  assign or1003  = a1003 | b1003;
  assign c1004 = (a1003 & b1003) | (a1003 & c1003) | (b1003 & c1003);
  wire c_sub1004;
  assign c_sub1004 = (a1003 & b_inv1003) | (a1003 & c1003) | (b_inv1003 & c1003);
  wire s1004, sub1004, and1004, or1004;
  wire b_inv1004;
  assign b_inv1004 = ~b1004;
  assign s1004  = a1004 ^ b1004 ^ c1004;
  assign sub1004 = a1004 ^ b_inv1004 ^ c1004;
  assign and1004 = a1004 & b1004;
  assign or1004  = a1004 | b1004;
  assign c1005 = (a1004 & b1004) | (a1004 & c1004) | (b1004 & c1004);
  wire c_sub1005;
  assign c_sub1005 = (a1004 & b_inv1004) | (a1004 & c1004) | (b_inv1004 & c1004);
  wire s1005, sub1005, and1005, or1005;
  wire b_inv1005;
  assign b_inv1005 = ~b1005;
  assign s1005  = a1005 ^ b1005 ^ c1005;
  assign sub1005 = a1005 ^ b_inv1005 ^ c1005;
  assign and1005 = a1005 & b1005;
  assign or1005  = a1005 | b1005;
  assign c1006 = (a1005 & b1005) | (a1005 & c1005) | (b1005 & c1005);
  wire c_sub1006;
  assign c_sub1006 = (a1005 & b_inv1005) | (a1005 & c1005) | (b_inv1005 & c1005);
  wire s1006, sub1006, and1006, or1006;
  wire b_inv1006;
  assign b_inv1006 = ~b1006;
  assign s1006  = a1006 ^ b1006 ^ c1006;
  assign sub1006 = a1006 ^ b_inv1006 ^ c1006;
  assign and1006 = a1006 & b1006;
  assign or1006  = a1006 | b1006;
  assign c1007 = (a1006 & b1006) | (a1006 & c1006) | (b1006 & c1006);
  wire c_sub1007;
  assign c_sub1007 = (a1006 & b_inv1006) | (a1006 & c1006) | (b_inv1006 & c1006);
  wire s1007, sub1007, and1007, or1007;
  wire b_inv1007;
  assign b_inv1007 = ~b1007;
  assign s1007  = a1007 ^ b1007 ^ c1007;
  assign sub1007 = a1007 ^ b_inv1007 ^ c1007;
  assign and1007 = a1007 & b1007;
  assign or1007  = a1007 | b1007;
  assign c1008 = (a1007 & b1007) | (a1007 & c1007) | (b1007 & c1007);
  wire c_sub1008;
  assign c_sub1008 = (a1007 & b_inv1007) | (a1007 & c1007) | (b_inv1007 & c1007);
  wire s1008, sub1008, and1008, or1008;
  wire b_inv1008;
  assign b_inv1008 = ~b1008;
  assign s1008  = a1008 ^ b1008 ^ c1008;
  assign sub1008 = a1008 ^ b_inv1008 ^ c1008;
  assign and1008 = a1008 & b1008;
  assign or1008  = a1008 | b1008;
  assign c1009 = (a1008 & b1008) | (a1008 & c1008) | (b1008 & c1008);
  wire c_sub1009;
  assign c_sub1009 = (a1008 & b_inv1008) | (a1008 & c1008) | (b_inv1008 & c1008);
  wire s1009, sub1009, and1009, or1009;
  wire b_inv1009;
  assign b_inv1009 = ~b1009;
  assign s1009  = a1009 ^ b1009 ^ c1009;
  assign sub1009 = a1009 ^ b_inv1009 ^ c1009;
  assign and1009 = a1009 & b1009;
  assign or1009  = a1009 | b1009;
  assign c1010 = (a1009 & b1009) | (a1009 & c1009) | (b1009 & c1009);
  wire c_sub1010;
  assign c_sub1010 = (a1009 & b_inv1009) | (a1009 & c1009) | (b_inv1009 & c1009);
  wire s1010, sub1010, and1010, or1010;
  wire b_inv1010;
  assign b_inv1010 = ~b1010;
  assign s1010  = a1010 ^ b1010 ^ c1010;
  assign sub1010 = a1010 ^ b_inv1010 ^ c1010;
  assign and1010 = a1010 & b1010;
  assign or1010  = a1010 | b1010;
  assign c1011 = (a1010 & b1010) | (a1010 & c1010) | (b1010 & c1010);
  wire c_sub1011;
  assign c_sub1011 = (a1010 & b_inv1010) | (a1010 & c1010) | (b_inv1010 & c1010);
  wire s1011, sub1011, and1011, or1011;
  wire b_inv1011;
  assign b_inv1011 = ~b1011;
  assign s1011  = a1011 ^ b1011 ^ c1011;
  assign sub1011 = a1011 ^ b_inv1011 ^ c1011;
  assign and1011 = a1011 & b1011;
  assign or1011  = a1011 | b1011;
  assign c1012 = (a1011 & b1011) | (a1011 & c1011) | (b1011 & c1011);
  wire c_sub1012;
  assign c_sub1012 = (a1011 & b_inv1011) | (a1011 & c1011) | (b_inv1011 & c1011);
  wire s1012, sub1012, and1012, or1012;
  wire b_inv1012;
  assign b_inv1012 = ~b1012;
  assign s1012  = a1012 ^ b1012 ^ c1012;
  assign sub1012 = a1012 ^ b_inv1012 ^ c1012;
  assign and1012 = a1012 & b1012;
  assign or1012  = a1012 | b1012;
  assign c1013 = (a1012 & b1012) | (a1012 & c1012) | (b1012 & c1012);
  wire c_sub1013;
  assign c_sub1013 = (a1012 & b_inv1012) | (a1012 & c1012) | (b_inv1012 & c1012);
  wire s1013, sub1013, and1013, or1013;
  wire b_inv1013;
  assign b_inv1013 = ~b1013;
  assign s1013  = a1013 ^ b1013 ^ c1013;
  assign sub1013 = a1013 ^ b_inv1013 ^ c1013;
  assign and1013 = a1013 & b1013;
  assign or1013  = a1013 | b1013;
  assign c1014 = (a1013 & b1013) | (a1013 & c1013) | (b1013 & c1013);
  wire c_sub1014;
  assign c_sub1014 = (a1013 & b_inv1013) | (a1013 & c1013) | (b_inv1013 & c1013);
  wire s1014, sub1014, and1014, or1014;
  wire b_inv1014;
  assign b_inv1014 = ~b1014;
  assign s1014  = a1014 ^ b1014 ^ c1014;
  assign sub1014 = a1014 ^ b_inv1014 ^ c1014;
  assign and1014 = a1014 & b1014;
  assign or1014  = a1014 | b1014;
  assign c1015 = (a1014 & b1014) | (a1014 & c1014) | (b1014 & c1014);
  wire c_sub1015;
  assign c_sub1015 = (a1014 & b_inv1014) | (a1014 & c1014) | (b_inv1014 & c1014);
  wire s1015, sub1015, and1015, or1015;
  wire b_inv1015;
  assign b_inv1015 = ~b1015;
  assign s1015  = a1015 ^ b1015 ^ c1015;
  assign sub1015 = a1015 ^ b_inv1015 ^ c1015;
  assign and1015 = a1015 & b1015;
  assign or1015  = a1015 | b1015;
  assign c1016 = (a1015 & b1015) | (a1015 & c1015) | (b1015 & c1015);
  wire c_sub1016;
  assign c_sub1016 = (a1015 & b_inv1015) | (a1015 & c1015) | (b_inv1015 & c1015);
  wire s1016, sub1016, and1016, or1016;
  wire b_inv1016;
  assign b_inv1016 = ~b1016;
  assign s1016  = a1016 ^ b1016 ^ c1016;
  assign sub1016 = a1016 ^ b_inv1016 ^ c1016;
  assign and1016 = a1016 & b1016;
  assign or1016  = a1016 | b1016;
  assign c1017 = (a1016 & b1016) | (a1016 & c1016) | (b1016 & c1016);
  wire c_sub1017;
  assign c_sub1017 = (a1016 & b_inv1016) | (a1016 & c1016) | (b_inv1016 & c1016);
  wire s1017, sub1017, and1017, or1017;
  wire b_inv1017;
  assign b_inv1017 = ~b1017;
  assign s1017  = a1017 ^ b1017 ^ c1017;
  assign sub1017 = a1017 ^ b_inv1017 ^ c1017;
  assign and1017 = a1017 & b1017;
  assign or1017  = a1017 | b1017;
  assign c1018 = (a1017 & b1017) | (a1017 & c1017) | (b1017 & c1017);
  wire c_sub1018;
  assign c_sub1018 = (a1017 & b_inv1017) | (a1017 & c1017) | (b_inv1017 & c1017);
  wire s1018, sub1018, and1018, or1018;
  wire b_inv1018;
  assign b_inv1018 = ~b1018;
  assign s1018  = a1018 ^ b1018 ^ c1018;
  assign sub1018 = a1018 ^ b_inv1018 ^ c1018;
  assign and1018 = a1018 & b1018;
  assign or1018  = a1018 | b1018;
  assign c1019 = (a1018 & b1018) | (a1018 & c1018) | (b1018 & c1018);
  wire c_sub1019;
  assign c_sub1019 = (a1018 & b_inv1018) | (a1018 & c1018) | (b_inv1018 & c1018);
  wire s1019, sub1019, and1019, or1019;
  wire b_inv1019;
  assign b_inv1019 = ~b1019;
  assign s1019  = a1019 ^ b1019 ^ c1019;
  assign sub1019 = a1019 ^ b_inv1019 ^ c1019;
  assign and1019 = a1019 & b1019;
  assign or1019  = a1019 | b1019;
  assign c1020 = (a1019 & b1019) | (a1019 & c1019) | (b1019 & c1019);
  wire c_sub1020;
  assign c_sub1020 = (a1019 & b_inv1019) | (a1019 & c1019) | (b_inv1019 & c1019);
  wire s1020, sub1020, and1020, or1020;
  wire b_inv1020;
  assign b_inv1020 = ~b1020;
  assign s1020  = a1020 ^ b1020 ^ c1020;
  assign sub1020 = a1020 ^ b_inv1020 ^ c1020;
  assign and1020 = a1020 & b1020;
  assign or1020  = a1020 | b1020;
  assign c1021 = (a1020 & b1020) | (a1020 & c1020) | (b1020 & c1020);
  wire c_sub1021;
  assign c_sub1021 = (a1020 & b_inv1020) | (a1020 & c1020) | (b_inv1020 & c1020);
  wire s1021, sub1021, and1021, or1021;
  wire b_inv1021;
  assign b_inv1021 = ~b1021;
  assign s1021  = a1021 ^ b1021 ^ c1021;
  assign sub1021 = a1021 ^ b_inv1021 ^ c1021;
  assign and1021 = a1021 & b1021;
  assign or1021  = a1021 | b1021;
  assign c1022 = (a1021 & b1021) | (a1021 & c1021) | (b1021 & c1021);
  wire c_sub1022;
  assign c_sub1022 = (a1021 & b_inv1021) | (a1021 & c1021) | (b_inv1021 & c1021);
  wire s1022, sub1022, and1022, or1022;
  wire b_inv1022;
  assign b_inv1022 = ~b1022;
  assign s1022  = a1022 ^ b1022 ^ c1022;
  assign sub1022 = a1022 ^ b_inv1022 ^ c1022;
  assign and1022 = a1022 & b1022;
  assign or1022  = a1022 | b1022;
  assign c1023 = (a1022 & b1022) | (a1022 & c1022) | (b1022 & c1022);
  wire c_sub1023;
  assign c_sub1023 = (a1022 & b_inv1022) | (a1022 & c1022) | (b_inv1022 & c1022);
  wire s1023, sub1023, and1023, or1023;
  wire b_inv1023;
  assign b_inv1023 = ~b1023;
  assign s1023  = a1023 ^ b1023 ^ c1023;
  assign sub1023 = a1023 ^ b_inv1023 ^ c1023;
  assign and1023 = a1023 & b1023;
  assign or1023  = a1023 | b1023;
  assign c1024 = (a1023 & b1023) | (a1023 & c1023) | (b1023 & c1023);
  wire c_sub1024;
  assign c_sub1024 = (a1023 & b_inv1023) | (a1023 & c1023) | (b_inv1023 & c1023);
  wire s1024, sub1024, and1024, or1024;
  wire b_inv1024;
  assign b_inv1024 = ~b1024;
  assign s1024  = a1024 ^ b1024 ^ c1024;
  assign sub1024 = a1024 ^ b_inv1024 ^ c1024;
  assign and1024 = a1024 & b1024;
  assign or1024  = a1024 | b1024;
  assign c1025 = (a1024 & b1024) | (a1024 & c1024) | (b1024 & c1024);
  wire c_sub1025;
  assign c_sub1025 = (a1024 & b_inv1024) | (a1024 & c1024) | (b_inv1024 & c1024);
  wire s1025, sub1025, and1025, or1025;
  wire b_inv1025;
  assign b_inv1025 = ~b1025;
  assign s1025  = a1025 ^ b1025 ^ c1025;
  assign sub1025 = a1025 ^ b_inv1025 ^ c1025;
  assign and1025 = a1025 & b1025;
  assign or1025  = a1025 | b1025;
  assign c1026 = (a1025 & b1025) | (a1025 & c1025) | (b1025 & c1025);
  wire c_sub1026;
  assign c_sub1026 = (a1025 & b_inv1025) | (a1025 & c1025) | (b_inv1025 & c1025);
  wire s1026, sub1026, and1026, or1026;
  wire b_inv1026;
  assign b_inv1026 = ~b1026;
  assign s1026  = a1026 ^ b1026 ^ c1026;
  assign sub1026 = a1026 ^ b_inv1026 ^ c1026;
  assign and1026 = a1026 & b1026;
  assign or1026  = a1026 | b1026;
  assign c1027 = (a1026 & b1026) | (a1026 & c1026) | (b1026 & c1026);
  wire c_sub1027;
  assign c_sub1027 = (a1026 & b_inv1026) | (a1026 & c1026) | (b_inv1026 & c1026);
  wire s1027, sub1027, and1027, or1027;
  wire b_inv1027;
  assign b_inv1027 = ~b1027;
  assign s1027  = a1027 ^ b1027 ^ c1027;
  assign sub1027 = a1027 ^ b_inv1027 ^ c1027;
  assign and1027 = a1027 & b1027;
  assign or1027  = a1027 | b1027;
  assign c1028 = (a1027 & b1027) | (a1027 & c1027) | (b1027 & c1027);
  wire c_sub1028;
  assign c_sub1028 = (a1027 & b_inv1027) | (a1027 & c1027) | (b_inv1027 & c1027);
  wire s1028, sub1028, and1028, or1028;
  wire b_inv1028;
  assign b_inv1028 = ~b1028;
  assign s1028  = a1028 ^ b1028 ^ c1028;
  assign sub1028 = a1028 ^ b_inv1028 ^ c1028;
  assign and1028 = a1028 & b1028;
  assign or1028  = a1028 | b1028;
  assign c1029 = (a1028 & b1028) | (a1028 & c1028) | (b1028 & c1028);
  wire c_sub1029;
  assign c_sub1029 = (a1028 & b_inv1028) | (a1028 & c1028) | (b_inv1028 & c1028);
  wire s1029, sub1029, and1029, or1029;
  wire b_inv1029;
  assign b_inv1029 = ~b1029;
  assign s1029  = a1029 ^ b1029 ^ c1029;
  assign sub1029 = a1029 ^ b_inv1029 ^ c1029;
  assign and1029 = a1029 & b1029;
  assign or1029  = a1029 | b1029;
  assign c1030 = (a1029 & b1029) | (a1029 & c1029) | (b1029 & c1029);
  wire c_sub1030;
  assign c_sub1030 = (a1029 & b_inv1029) | (a1029 & c1029) | (b_inv1029 & c1029);
  wire s1030, sub1030, and1030, or1030;
  wire b_inv1030;
  assign b_inv1030 = ~b1030;
  assign s1030  = a1030 ^ b1030 ^ c1030;
  assign sub1030 = a1030 ^ b_inv1030 ^ c1030;
  assign and1030 = a1030 & b1030;
  assign or1030  = a1030 | b1030;
  assign c1031 = (a1030 & b1030) | (a1030 & c1030) | (b1030 & c1030);
  wire c_sub1031;
  assign c_sub1031 = (a1030 & b_inv1030) | (a1030 & c1030) | (b_inv1030 & c1030);
  wire s1031, sub1031, and1031, or1031;
  wire b_inv1031;
  assign b_inv1031 = ~b1031;
  assign s1031  = a1031 ^ b1031 ^ c1031;
  assign sub1031 = a1031 ^ b_inv1031 ^ c1031;
  assign and1031 = a1031 & b1031;
  assign or1031  = a1031 | b1031;
  assign c1032 = (a1031 & b1031) | (a1031 & c1031) | (b1031 & c1031);
  wire c_sub1032;
  assign c_sub1032 = (a1031 & b_inv1031) | (a1031 & c1031) | (b_inv1031 & c1031);
  wire s1032, sub1032, and1032, or1032;
  wire b_inv1032;
  assign b_inv1032 = ~b1032;
  assign s1032  = a1032 ^ b1032 ^ c1032;
  assign sub1032 = a1032 ^ b_inv1032 ^ c1032;
  assign and1032 = a1032 & b1032;
  assign or1032  = a1032 | b1032;
  assign c1033 = (a1032 & b1032) | (a1032 & c1032) | (b1032 & c1032);
  wire c_sub1033;
  assign c_sub1033 = (a1032 & b_inv1032) | (a1032 & c1032) | (b_inv1032 & c1032);
  wire s1033, sub1033, and1033, or1033;
  wire b_inv1033;
  assign b_inv1033 = ~b1033;
  assign s1033  = a1033 ^ b1033 ^ c1033;
  assign sub1033 = a1033 ^ b_inv1033 ^ c1033;
  assign and1033 = a1033 & b1033;
  assign or1033  = a1033 | b1033;
  assign c1034 = (a1033 & b1033) | (a1033 & c1033) | (b1033 & c1033);
  wire c_sub1034;
  assign c_sub1034 = (a1033 & b_inv1033) | (a1033 & c1033) | (b_inv1033 & c1033);
  wire s1034, sub1034, and1034, or1034;
  wire b_inv1034;
  assign b_inv1034 = ~b1034;
  assign s1034  = a1034 ^ b1034 ^ c1034;
  assign sub1034 = a1034 ^ b_inv1034 ^ c1034;
  assign and1034 = a1034 & b1034;
  assign or1034  = a1034 | b1034;
  assign c1035 = (a1034 & b1034) | (a1034 & c1034) | (b1034 & c1034);
  wire c_sub1035;
  assign c_sub1035 = (a1034 & b_inv1034) | (a1034 & c1034) | (b_inv1034 & c1034);
  wire s1035, sub1035, and1035, or1035;
  wire b_inv1035;
  assign b_inv1035 = ~b1035;
  assign s1035  = a1035 ^ b1035 ^ c1035;
  assign sub1035 = a1035 ^ b_inv1035 ^ c1035;
  assign and1035 = a1035 & b1035;
  assign or1035  = a1035 | b1035;
  assign c1036 = (a1035 & b1035) | (a1035 & c1035) | (b1035 & c1035);
  wire c_sub1036;
  assign c_sub1036 = (a1035 & b_inv1035) | (a1035 & c1035) | (b_inv1035 & c1035);
  wire s1036, sub1036, and1036, or1036;
  wire b_inv1036;
  assign b_inv1036 = ~b1036;
  assign s1036  = a1036 ^ b1036 ^ c1036;
  assign sub1036 = a1036 ^ b_inv1036 ^ c1036;
  assign and1036 = a1036 & b1036;
  assign or1036  = a1036 | b1036;
  assign c1037 = (a1036 & b1036) | (a1036 & c1036) | (b1036 & c1036);
  wire c_sub1037;
  assign c_sub1037 = (a1036 & b_inv1036) | (a1036 & c1036) | (b_inv1036 & c1036);
  wire s1037, sub1037, and1037, or1037;
  wire b_inv1037;
  assign b_inv1037 = ~b1037;
  assign s1037  = a1037 ^ b1037 ^ c1037;
  assign sub1037 = a1037 ^ b_inv1037 ^ c1037;
  assign and1037 = a1037 & b1037;
  assign or1037  = a1037 | b1037;
  assign c1038 = (a1037 & b1037) | (a1037 & c1037) | (b1037 & c1037);
  wire c_sub1038;
  assign c_sub1038 = (a1037 & b_inv1037) | (a1037 & c1037) | (b_inv1037 & c1037);
  wire s1038, sub1038, and1038, or1038;
  wire b_inv1038;
  assign b_inv1038 = ~b1038;
  assign s1038  = a1038 ^ b1038 ^ c1038;
  assign sub1038 = a1038 ^ b_inv1038 ^ c1038;
  assign and1038 = a1038 & b1038;
  assign or1038  = a1038 | b1038;
  assign c1039 = (a1038 & b1038) | (a1038 & c1038) | (b1038 & c1038);
  wire c_sub1039;
  assign c_sub1039 = (a1038 & b_inv1038) | (a1038 & c1038) | (b_inv1038 & c1038);
  wire s1039, sub1039, and1039, or1039;
  wire b_inv1039;
  assign b_inv1039 = ~b1039;
  assign s1039  = a1039 ^ b1039 ^ c1039;
  assign sub1039 = a1039 ^ b_inv1039 ^ c1039;
  assign and1039 = a1039 & b1039;
  assign or1039  = a1039 | b1039;
  assign c1040 = (a1039 & b1039) | (a1039 & c1039) | (b1039 & c1039);
  wire c_sub1040;
  assign c_sub1040 = (a1039 & b_inv1039) | (a1039 & c1039) | (b_inv1039 & c1039);
  wire s1040, sub1040, and1040, or1040;
  wire b_inv1040;
  assign b_inv1040 = ~b1040;
  assign s1040  = a1040 ^ b1040 ^ c1040;
  assign sub1040 = a1040 ^ b_inv1040 ^ c1040;
  assign and1040 = a1040 & b1040;
  assign or1040  = a1040 | b1040;
  assign c1041 = (a1040 & b1040) | (a1040 & c1040) | (b1040 & c1040);
  wire c_sub1041;
  assign c_sub1041 = (a1040 & b_inv1040) | (a1040 & c1040) | (b_inv1040 & c1040);
  wire s1041, sub1041, and1041, or1041;
  wire b_inv1041;
  assign b_inv1041 = ~b1041;
  assign s1041  = a1041 ^ b1041 ^ c1041;
  assign sub1041 = a1041 ^ b_inv1041 ^ c1041;
  assign and1041 = a1041 & b1041;
  assign or1041  = a1041 | b1041;
  assign c1042 = (a1041 & b1041) | (a1041 & c1041) | (b1041 & c1041);
  wire c_sub1042;
  assign c_sub1042 = (a1041 & b_inv1041) | (a1041 & c1041) | (b_inv1041 & c1041);
  wire s1042, sub1042, and1042, or1042;
  wire b_inv1042;
  assign b_inv1042 = ~b1042;
  assign s1042  = a1042 ^ b1042 ^ c1042;
  assign sub1042 = a1042 ^ b_inv1042 ^ c1042;
  assign and1042 = a1042 & b1042;
  assign or1042  = a1042 | b1042;
  assign c1043 = (a1042 & b1042) | (a1042 & c1042) | (b1042 & c1042);
  wire c_sub1043;
  assign c_sub1043 = (a1042 & b_inv1042) | (a1042 & c1042) | (b_inv1042 & c1042);
  wire s1043, sub1043, and1043, or1043;
  wire b_inv1043;
  assign b_inv1043 = ~b1043;
  assign s1043  = a1043 ^ b1043 ^ c1043;
  assign sub1043 = a1043 ^ b_inv1043 ^ c1043;
  assign and1043 = a1043 & b1043;
  assign or1043  = a1043 | b1043;
  assign c1044 = (a1043 & b1043) | (a1043 & c1043) | (b1043 & c1043);
  wire c_sub1044;
  assign c_sub1044 = (a1043 & b_inv1043) | (a1043 & c1043) | (b_inv1043 & c1043);
  wire s1044, sub1044, and1044, or1044;
  wire b_inv1044;
  assign b_inv1044 = ~b1044;
  assign s1044  = a1044 ^ b1044 ^ c1044;
  assign sub1044 = a1044 ^ b_inv1044 ^ c1044;
  assign and1044 = a1044 & b1044;
  assign or1044  = a1044 | b1044;
  assign c1045 = (a1044 & b1044) | (a1044 & c1044) | (b1044 & c1044);
  wire c_sub1045;
  assign c_sub1045 = (a1044 & b_inv1044) | (a1044 & c1044) | (b_inv1044 & c1044);
  wire s1045, sub1045, and1045, or1045;
  wire b_inv1045;
  assign b_inv1045 = ~b1045;
  assign s1045  = a1045 ^ b1045 ^ c1045;
  assign sub1045 = a1045 ^ b_inv1045 ^ c1045;
  assign and1045 = a1045 & b1045;
  assign or1045  = a1045 | b1045;
  assign c1046 = (a1045 & b1045) | (a1045 & c1045) | (b1045 & c1045);
  wire c_sub1046;
  assign c_sub1046 = (a1045 & b_inv1045) | (a1045 & c1045) | (b_inv1045 & c1045);
  wire s1046, sub1046, and1046, or1046;
  wire b_inv1046;
  assign b_inv1046 = ~b1046;
  assign s1046  = a1046 ^ b1046 ^ c1046;
  assign sub1046 = a1046 ^ b_inv1046 ^ c1046;
  assign and1046 = a1046 & b1046;
  assign or1046  = a1046 | b1046;
  assign c1047 = (a1046 & b1046) | (a1046 & c1046) | (b1046 & c1046);
  wire c_sub1047;
  assign c_sub1047 = (a1046 & b_inv1046) | (a1046 & c1046) | (b_inv1046 & c1046);
  wire s1047, sub1047, and1047, or1047;
  wire b_inv1047;
  assign b_inv1047 = ~b1047;
  assign s1047  = a1047 ^ b1047 ^ c1047;
  assign sub1047 = a1047 ^ b_inv1047 ^ c1047;
  assign and1047 = a1047 & b1047;
  assign or1047  = a1047 | b1047;
  assign c1048 = (a1047 & b1047) | (a1047 & c1047) | (b1047 & c1047);
  wire c_sub1048;
  assign c_sub1048 = (a1047 & b_inv1047) | (a1047 & c1047) | (b_inv1047 & c1047);
  wire s1048, sub1048, and1048, or1048;
  wire b_inv1048;
  assign b_inv1048 = ~b1048;
  assign s1048  = a1048 ^ b1048 ^ c1048;
  assign sub1048 = a1048 ^ b_inv1048 ^ c1048;
  assign and1048 = a1048 & b1048;
  assign or1048  = a1048 | b1048;
  assign c1049 = (a1048 & b1048) | (a1048 & c1048) | (b1048 & c1048);
  wire c_sub1049;
  assign c_sub1049 = (a1048 & b_inv1048) | (a1048 & c1048) | (b_inv1048 & c1048);
  wire s1049, sub1049, and1049, or1049;
  wire b_inv1049;
  assign b_inv1049 = ~b1049;
  assign s1049  = a1049 ^ b1049 ^ c1049;
  assign sub1049 = a1049 ^ b_inv1049 ^ c1049;
  assign and1049 = a1049 & b1049;
  assign or1049  = a1049 | b1049;
  assign c1050 = (a1049 & b1049) | (a1049 & c1049) | (b1049 & c1049);
  wire c_sub1050;
  assign c_sub1050 = (a1049 & b_inv1049) | (a1049 & c1049) | (b_inv1049 & c1049);
  wire s1050, sub1050, and1050, or1050;
  wire b_inv1050;
  assign b_inv1050 = ~b1050;
  assign s1050  = a1050 ^ b1050 ^ c1050;
  assign sub1050 = a1050 ^ b_inv1050 ^ c1050;
  assign and1050 = a1050 & b1050;
  assign or1050  = a1050 | b1050;
  assign c1051 = (a1050 & b1050) | (a1050 & c1050) | (b1050 & c1050);
  wire c_sub1051;
  assign c_sub1051 = (a1050 & b_inv1050) | (a1050 & c1050) | (b_inv1050 & c1050);
  wire s1051, sub1051, and1051, or1051;
  wire b_inv1051;
  assign b_inv1051 = ~b1051;
  assign s1051  = a1051 ^ b1051 ^ c1051;
  assign sub1051 = a1051 ^ b_inv1051 ^ c1051;
  assign and1051 = a1051 & b1051;
  assign or1051  = a1051 | b1051;
  assign c1052 = (a1051 & b1051) | (a1051 & c1051) | (b1051 & c1051);
  wire c_sub1052;
  assign c_sub1052 = (a1051 & b_inv1051) | (a1051 & c1051) | (b_inv1051 & c1051);
  wire s1052, sub1052, and1052, or1052;
  wire b_inv1052;
  assign b_inv1052 = ~b1052;
  assign s1052  = a1052 ^ b1052 ^ c1052;
  assign sub1052 = a1052 ^ b_inv1052 ^ c1052;
  assign and1052 = a1052 & b1052;
  assign or1052  = a1052 | b1052;
  assign c1053 = (a1052 & b1052) | (a1052 & c1052) | (b1052 & c1052);
  wire c_sub1053;
  assign c_sub1053 = (a1052 & b_inv1052) | (a1052 & c1052) | (b_inv1052 & c1052);
  wire s1053, sub1053, and1053, or1053;
  wire b_inv1053;
  assign b_inv1053 = ~b1053;
  assign s1053  = a1053 ^ b1053 ^ c1053;
  assign sub1053 = a1053 ^ b_inv1053 ^ c1053;
  assign and1053 = a1053 & b1053;
  assign or1053  = a1053 | b1053;
  assign c1054 = (a1053 & b1053) | (a1053 & c1053) | (b1053 & c1053);
  wire c_sub1054;
  assign c_sub1054 = (a1053 & b_inv1053) | (a1053 & c1053) | (b_inv1053 & c1053);
  wire s1054, sub1054, and1054, or1054;
  wire b_inv1054;
  assign b_inv1054 = ~b1054;
  assign s1054  = a1054 ^ b1054 ^ c1054;
  assign sub1054 = a1054 ^ b_inv1054 ^ c1054;
  assign and1054 = a1054 & b1054;
  assign or1054  = a1054 | b1054;
  assign c1055 = (a1054 & b1054) | (a1054 & c1054) | (b1054 & c1054);
  wire c_sub1055;
  assign c_sub1055 = (a1054 & b_inv1054) | (a1054 & c1054) | (b_inv1054 & c1054);
  wire s1055, sub1055, and1055, or1055;
  wire b_inv1055;
  assign b_inv1055 = ~b1055;
  assign s1055  = a1055 ^ b1055 ^ c1055;
  assign sub1055 = a1055 ^ b_inv1055 ^ c1055;
  assign and1055 = a1055 & b1055;
  assign or1055  = a1055 | b1055;
  assign c1056 = (a1055 & b1055) | (a1055 & c1055) | (b1055 & c1055);
  wire c_sub1056;
  assign c_sub1056 = (a1055 & b_inv1055) | (a1055 & c1055) | (b_inv1055 & c1055);
  wire s1056, sub1056, and1056, or1056;
  wire b_inv1056;
  assign b_inv1056 = ~b1056;
  assign s1056  = a1056 ^ b1056 ^ c1056;
  assign sub1056 = a1056 ^ b_inv1056 ^ c1056;
  assign and1056 = a1056 & b1056;
  assign or1056  = a1056 | b1056;
  assign c1057 = (a1056 & b1056) | (a1056 & c1056) | (b1056 & c1056);
  wire c_sub1057;
  assign c_sub1057 = (a1056 & b_inv1056) | (a1056 & c1056) | (b_inv1056 & c1056);
  wire s1057, sub1057, and1057, or1057;
  wire b_inv1057;
  assign b_inv1057 = ~b1057;
  assign s1057  = a1057 ^ b1057 ^ c1057;
  assign sub1057 = a1057 ^ b_inv1057 ^ c1057;
  assign and1057 = a1057 & b1057;
  assign or1057  = a1057 | b1057;
  assign c1058 = (a1057 & b1057) | (a1057 & c1057) | (b1057 & c1057);
  wire c_sub1058;
  assign c_sub1058 = (a1057 & b_inv1057) | (a1057 & c1057) | (b_inv1057 & c1057);
  wire s1058, sub1058, and1058, or1058;
  wire b_inv1058;
  assign b_inv1058 = ~b1058;
  assign s1058  = a1058 ^ b1058 ^ c1058;
  assign sub1058 = a1058 ^ b_inv1058 ^ c1058;
  assign and1058 = a1058 & b1058;
  assign or1058  = a1058 | b1058;
  assign c1059 = (a1058 & b1058) | (a1058 & c1058) | (b1058 & c1058);
  wire c_sub1059;
  assign c_sub1059 = (a1058 & b_inv1058) | (a1058 & c1058) | (b_inv1058 & c1058);
  wire s1059, sub1059, and1059, or1059;
  wire b_inv1059;
  assign b_inv1059 = ~b1059;
  assign s1059  = a1059 ^ b1059 ^ c1059;
  assign sub1059 = a1059 ^ b_inv1059 ^ c1059;
  assign and1059 = a1059 & b1059;
  assign or1059  = a1059 | b1059;
  assign c1060 = (a1059 & b1059) | (a1059 & c1059) | (b1059 & c1059);
  wire c_sub1060;
  assign c_sub1060 = (a1059 & b_inv1059) | (a1059 & c1059) | (b_inv1059 & c1059);
  wire s1060, sub1060, and1060, or1060;
  wire b_inv1060;
  assign b_inv1060 = ~b1060;
  assign s1060  = a1060 ^ b1060 ^ c1060;
  assign sub1060 = a1060 ^ b_inv1060 ^ c1060;
  assign and1060 = a1060 & b1060;
  assign or1060  = a1060 | b1060;
  assign c1061 = (a1060 & b1060) | (a1060 & c1060) | (b1060 & c1060);
  wire c_sub1061;
  assign c_sub1061 = (a1060 & b_inv1060) | (a1060 & c1060) | (b_inv1060 & c1060);
  wire s1061, sub1061, and1061, or1061;
  wire b_inv1061;
  assign b_inv1061 = ~b1061;
  assign s1061  = a1061 ^ b1061 ^ c1061;
  assign sub1061 = a1061 ^ b_inv1061 ^ c1061;
  assign and1061 = a1061 & b1061;
  assign or1061  = a1061 | b1061;
  assign c1062 = (a1061 & b1061) | (a1061 & c1061) | (b1061 & c1061);
  wire c_sub1062;
  assign c_sub1062 = (a1061 & b_inv1061) | (a1061 & c1061) | (b_inv1061 & c1061);
  wire s1062, sub1062, and1062, or1062;
  wire b_inv1062;
  assign b_inv1062 = ~b1062;
  assign s1062  = a1062 ^ b1062 ^ c1062;
  assign sub1062 = a1062 ^ b_inv1062 ^ c1062;
  assign and1062 = a1062 & b1062;
  assign or1062  = a1062 | b1062;
  assign c1063 = (a1062 & b1062) | (a1062 & c1062) | (b1062 & c1062);
  wire c_sub1063;
  assign c_sub1063 = (a1062 & b_inv1062) | (a1062 & c1062) | (b_inv1062 & c1062);
  wire s1063, sub1063, and1063, or1063;
  wire b_inv1063;
  assign b_inv1063 = ~b1063;
  assign s1063  = a1063 ^ b1063 ^ c1063;
  assign sub1063 = a1063 ^ b_inv1063 ^ c1063;
  assign and1063 = a1063 & b1063;
  assign or1063  = a1063 | b1063;
  assign c1064 = (a1063 & b1063) | (a1063 & c1063) | (b1063 & c1063);
  wire c_sub1064;
  assign c_sub1064 = (a1063 & b_inv1063) | (a1063 & c1063) | (b_inv1063 & c1063);
  wire s1064, sub1064, and1064, or1064;
  wire b_inv1064;
  assign b_inv1064 = ~b1064;
  assign s1064  = a1064 ^ b1064 ^ c1064;
  assign sub1064 = a1064 ^ b_inv1064 ^ c1064;
  assign and1064 = a1064 & b1064;
  assign or1064  = a1064 | b1064;
  assign c1065 = (a1064 & b1064) | (a1064 & c1064) | (b1064 & c1064);
  wire c_sub1065;
  assign c_sub1065 = (a1064 & b_inv1064) | (a1064 & c1064) | (b_inv1064 & c1064);
  wire s1065, sub1065, and1065, or1065;
  wire b_inv1065;
  assign b_inv1065 = ~b1065;
  assign s1065  = a1065 ^ b1065 ^ c1065;
  assign sub1065 = a1065 ^ b_inv1065 ^ c1065;
  assign and1065 = a1065 & b1065;
  assign or1065  = a1065 | b1065;
  assign c1066 = (a1065 & b1065) | (a1065 & c1065) | (b1065 & c1065);
  wire c_sub1066;
  assign c_sub1066 = (a1065 & b_inv1065) | (a1065 & c1065) | (b_inv1065 & c1065);
  wire s1066, sub1066, and1066, or1066;
  wire b_inv1066;
  assign b_inv1066 = ~b1066;
  assign s1066  = a1066 ^ b1066 ^ c1066;
  assign sub1066 = a1066 ^ b_inv1066 ^ c1066;
  assign and1066 = a1066 & b1066;
  assign or1066  = a1066 | b1066;
  assign c1067 = (a1066 & b1066) | (a1066 & c1066) | (b1066 & c1066);
  wire c_sub1067;
  assign c_sub1067 = (a1066 & b_inv1066) | (a1066 & c1066) | (b_inv1066 & c1066);
  wire s1067, sub1067, and1067, or1067;
  wire b_inv1067;
  assign b_inv1067 = ~b1067;
  assign s1067  = a1067 ^ b1067 ^ c1067;
  assign sub1067 = a1067 ^ b_inv1067 ^ c1067;
  assign and1067 = a1067 & b1067;
  assign or1067  = a1067 | b1067;
  assign c1068 = (a1067 & b1067) | (a1067 & c1067) | (b1067 & c1067);
  wire c_sub1068;
  assign c_sub1068 = (a1067 & b_inv1067) | (a1067 & c1067) | (b_inv1067 & c1067);
  wire s1068, sub1068, and1068, or1068;
  wire b_inv1068;
  assign b_inv1068 = ~b1068;
  assign s1068  = a1068 ^ b1068 ^ c1068;
  assign sub1068 = a1068 ^ b_inv1068 ^ c1068;
  assign and1068 = a1068 & b1068;
  assign or1068  = a1068 | b1068;
  assign c1069 = (a1068 & b1068) | (a1068 & c1068) | (b1068 & c1068);
  wire c_sub1069;
  assign c_sub1069 = (a1068 & b_inv1068) | (a1068 & c1068) | (b_inv1068 & c1068);
  wire s1069, sub1069, and1069, or1069;
  wire b_inv1069;
  assign b_inv1069 = ~b1069;
  assign s1069  = a1069 ^ b1069 ^ c1069;
  assign sub1069 = a1069 ^ b_inv1069 ^ c1069;
  assign and1069 = a1069 & b1069;
  assign or1069  = a1069 | b1069;
  assign c1070 = (a1069 & b1069) | (a1069 & c1069) | (b1069 & c1069);
  wire c_sub1070;
  assign c_sub1070 = (a1069 & b_inv1069) | (a1069 & c1069) | (b_inv1069 & c1069);
  wire s1070, sub1070, and1070, or1070;
  wire b_inv1070;
  assign b_inv1070 = ~b1070;
  assign s1070  = a1070 ^ b1070 ^ c1070;
  assign sub1070 = a1070 ^ b_inv1070 ^ c1070;
  assign and1070 = a1070 & b1070;
  assign or1070  = a1070 | b1070;
  assign c1071 = (a1070 & b1070) | (a1070 & c1070) | (b1070 & c1070);
  wire c_sub1071;
  assign c_sub1071 = (a1070 & b_inv1070) | (a1070 & c1070) | (b_inv1070 & c1070);
  wire s1071, sub1071, and1071, or1071;
  wire b_inv1071;
  assign b_inv1071 = ~b1071;
  assign s1071  = a1071 ^ b1071 ^ c1071;
  assign sub1071 = a1071 ^ b_inv1071 ^ c1071;
  assign and1071 = a1071 & b1071;
  assign or1071  = a1071 | b1071;
  assign c1072 = (a1071 & b1071) | (a1071 & c1071) | (b1071 & c1071);
  wire c_sub1072;
  assign c_sub1072 = (a1071 & b_inv1071) | (a1071 & c1071) | (b_inv1071 & c1071);
  wire s1072, sub1072, and1072, or1072;
  wire b_inv1072;
  assign b_inv1072 = ~b1072;
  assign s1072  = a1072 ^ b1072 ^ c1072;
  assign sub1072 = a1072 ^ b_inv1072 ^ c1072;
  assign and1072 = a1072 & b1072;
  assign or1072  = a1072 | b1072;
  assign c1073 = (a1072 & b1072) | (a1072 & c1072) | (b1072 & c1072);
  wire c_sub1073;
  assign c_sub1073 = (a1072 & b_inv1072) | (a1072 & c1072) | (b_inv1072 & c1072);
  wire s1073, sub1073, and1073, or1073;
  wire b_inv1073;
  assign b_inv1073 = ~b1073;
  assign s1073  = a1073 ^ b1073 ^ c1073;
  assign sub1073 = a1073 ^ b_inv1073 ^ c1073;
  assign and1073 = a1073 & b1073;
  assign or1073  = a1073 | b1073;
  assign c1074 = (a1073 & b1073) | (a1073 & c1073) | (b1073 & c1073);
  wire c_sub1074;
  assign c_sub1074 = (a1073 & b_inv1073) | (a1073 & c1073) | (b_inv1073 & c1073);
  wire s1074, sub1074, and1074, or1074;
  wire b_inv1074;
  assign b_inv1074 = ~b1074;
  assign s1074  = a1074 ^ b1074 ^ c1074;
  assign sub1074 = a1074 ^ b_inv1074 ^ c1074;
  assign and1074 = a1074 & b1074;
  assign or1074  = a1074 | b1074;
  assign c1075 = (a1074 & b1074) | (a1074 & c1074) | (b1074 & c1074);
  wire c_sub1075;
  assign c_sub1075 = (a1074 & b_inv1074) | (a1074 & c1074) | (b_inv1074 & c1074);
  wire s1075, sub1075, and1075, or1075;
  wire b_inv1075;
  assign b_inv1075 = ~b1075;
  assign s1075  = a1075 ^ b1075 ^ c1075;
  assign sub1075 = a1075 ^ b_inv1075 ^ c1075;
  assign and1075 = a1075 & b1075;
  assign or1075  = a1075 | b1075;
  assign c1076 = (a1075 & b1075) | (a1075 & c1075) | (b1075 & c1075);
  wire c_sub1076;
  assign c_sub1076 = (a1075 & b_inv1075) | (a1075 & c1075) | (b_inv1075 & c1075);
  wire s1076, sub1076, and1076, or1076;
  wire b_inv1076;
  assign b_inv1076 = ~b1076;
  assign s1076  = a1076 ^ b1076 ^ c1076;
  assign sub1076 = a1076 ^ b_inv1076 ^ c1076;
  assign and1076 = a1076 & b1076;
  assign or1076  = a1076 | b1076;
  assign c1077 = (a1076 & b1076) | (a1076 & c1076) | (b1076 & c1076);
  wire c_sub1077;
  assign c_sub1077 = (a1076 & b_inv1076) | (a1076 & c1076) | (b_inv1076 & c1076);
  wire s1077, sub1077, and1077, or1077;
  wire b_inv1077;
  assign b_inv1077 = ~b1077;
  assign s1077  = a1077 ^ b1077 ^ c1077;
  assign sub1077 = a1077 ^ b_inv1077 ^ c1077;
  assign and1077 = a1077 & b1077;
  assign or1077  = a1077 | b1077;
  assign c1078 = (a1077 & b1077) | (a1077 & c1077) | (b1077 & c1077);
  wire c_sub1078;
  assign c_sub1078 = (a1077 & b_inv1077) | (a1077 & c1077) | (b_inv1077 & c1077);
  wire s1078, sub1078, and1078, or1078;
  wire b_inv1078;
  assign b_inv1078 = ~b1078;
  assign s1078  = a1078 ^ b1078 ^ c1078;
  assign sub1078 = a1078 ^ b_inv1078 ^ c1078;
  assign and1078 = a1078 & b1078;
  assign or1078  = a1078 | b1078;
  assign c1079 = (a1078 & b1078) | (a1078 & c1078) | (b1078 & c1078);
  wire c_sub1079;
  assign c_sub1079 = (a1078 & b_inv1078) | (a1078 & c1078) | (b_inv1078 & c1078);
  wire s1079, sub1079, and1079, or1079;
  wire b_inv1079;
  assign b_inv1079 = ~b1079;
  assign s1079  = a1079 ^ b1079 ^ c1079;
  assign sub1079 = a1079 ^ b_inv1079 ^ c1079;
  assign and1079 = a1079 & b1079;
  assign or1079  = a1079 | b1079;
  assign c1080 = (a1079 & b1079) | (a1079 & c1079) | (b1079 & c1079);
  wire c_sub1080;
  assign c_sub1080 = (a1079 & b_inv1079) | (a1079 & c1079) | (b_inv1079 & c1079);
  wire s1080, sub1080, and1080, or1080;
  wire b_inv1080;
  assign b_inv1080 = ~b1080;
  assign s1080  = a1080 ^ b1080 ^ c1080;
  assign sub1080 = a1080 ^ b_inv1080 ^ c1080;
  assign and1080 = a1080 & b1080;
  assign or1080  = a1080 | b1080;
  assign c1081 = (a1080 & b1080) | (a1080 & c1080) | (b1080 & c1080);
  wire c_sub1081;
  assign c_sub1081 = (a1080 & b_inv1080) | (a1080 & c1080) | (b_inv1080 & c1080);
  wire s1081, sub1081, and1081, or1081;
  wire b_inv1081;
  assign b_inv1081 = ~b1081;
  assign s1081  = a1081 ^ b1081 ^ c1081;
  assign sub1081 = a1081 ^ b_inv1081 ^ c1081;
  assign and1081 = a1081 & b1081;
  assign or1081  = a1081 | b1081;
  assign c1082 = (a1081 & b1081) | (a1081 & c1081) | (b1081 & c1081);
  wire c_sub1082;
  assign c_sub1082 = (a1081 & b_inv1081) | (a1081 & c1081) | (b_inv1081 & c1081);
  wire s1082, sub1082, and1082, or1082;
  wire b_inv1082;
  assign b_inv1082 = ~b1082;
  assign s1082  = a1082 ^ b1082 ^ c1082;
  assign sub1082 = a1082 ^ b_inv1082 ^ c1082;
  assign and1082 = a1082 & b1082;
  assign or1082  = a1082 | b1082;
  assign c1083 = (a1082 & b1082) | (a1082 & c1082) | (b1082 & c1082);
  wire c_sub1083;
  assign c_sub1083 = (a1082 & b_inv1082) | (a1082 & c1082) | (b_inv1082 & c1082);
  wire s1083, sub1083, and1083, or1083;
  wire b_inv1083;
  assign b_inv1083 = ~b1083;
  assign s1083  = a1083 ^ b1083 ^ c1083;
  assign sub1083 = a1083 ^ b_inv1083 ^ c1083;
  assign and1083 = a1083 & b1083;
  assign or1083  = a1083 | b1083;
  assign c1084 = (a1083 & b1083) | (a1083 & c1083) | (b1083 & c1083);
  wire c_sub1084;
  assign c_sub1084 = (a1083 & b_inv1083) | (a1083 & c1083) | (b_inv1083 & c1083);
  wire s1084, sub1084, and1084, or1084;
  wire b_inv1084;
  assign b_inv1084 = ~b1084;
  assign s1084  = a1084 ^ b1084 ^ c1084;
  assign sub1084 = a1084 ^ b_inv1084 ^ c1084;
  assign and1084 = a1084 & b1084;
  assign or1084  = a1084 | b1084;
  assign c1085 = (a1084 & b1084) | (a1084 & c1084) | (b1084 & c1084);
  wire c_sub1085;
  assign c_sub1085 = (a1084 & b_inv1084) | (a1084 & c1084) | (b_inv1084 & c1084);
  wire s1085, sub1085, and1085, or1085;
  wire b_inv1085;
  assign b_inv1085 = ~b1085;
  assign s1085  = a1085 ^ b1085 ^ c1085;
  assign sub1085 = a1085 ^ b_inv1085 ^ c1085;
  assign and1085 = a1085 & b1085;
  assign or1085  = a1085 | b1085;
  assign c1086 = (a1085 & b1085) | (a1085 & c1085) | (b1085 & c1085);
  wire c_sub1086;
  assign c_sub1086 = (a1085 & b_inv1085) | (a1085 & c1085) | (b_inv1085 & c1085);
  wire s1086, sub1086, and1086, or1086;
  wire b_inv1086;
  assign b_inv1086 = ~b1086;
  assign s1086  = a1086 ^ b1086 ^ c1086;
  assign sub1086 = a1086 ^ b_inv1086 ^ c1086;
  assign and1086 = a1086 & b1086;
  assign or1086  = a1086 | b1086;
  assign c1087 = (a1086 & b1086) | (a1086 & c1086) | (b1086 & c1086);
  wire c_sub1087;
  assign c_sub1087 = (a1086 & b_inv1086) | (a1086 & c1086) | (b_inv1086 & c1086);
  wire s1087, sub1087, and1087, or1087;
  wire b_inv1087;
  assign b_inv1087 = ~b1087;
  assign s1087  = a1087 ^ b1087 ^ c1087;
  assign sub1087 = a1087 ^ b_inv1087 ^ c1087;
  assign and1087 = a1087 & b1087;
  assign or1087  = a1087 | b1087;
  assign c1088 = (a1087 & b1087) | (a1087 & c1087) | (b1087 & c1087);
  wire c_sub1088;
  assign c_sub1088 = (a1087 & b_inv1087) | (a1087 & c1087) | (b_inv1087 & c1087);
  wire s1088, sub1088, and1088, or1088;
  wire b_inv1088;
  assign b_inv1088 = ~b1088;
  assign s1088  = a1088 ^ b1088 ^ c1088;
  assign sub1088 = a1088 ^ b_inv1088 ^ c1088;
  assign and1088 = a1088 & b1088;
  assign or1088  = a1088 | b1088;
  assign c1089 = (a1088 & b1088) | (a1088 & c1088) | (b1088 & c1088);
  wire c_sub1089;
  assign c_sub1089 = (a1088 & b_inv1088) | (a1088 & c1088) | (b_inv1088 & c1088);
  wire s1089, sub1089, and1089, or1089;
  wire b_inv1089;
  assign b_inv1089 = ~b1089;
  assign s1089  = a1089 ^ b1089 ^ c1089;
  assign sub1089 = a1089 ^ b_inv1089 ^ c1089;
  assign and1089 = a1089 & b1089;
  assign or1089  = a1089 | b1089;
  assign c1090 = (a1089 & b1089) | (a1089 & c1089) | (b1089 & c1089);
  wire c_sub1090;
  assign c_sub1090 = (a1089 & b_inv1089) | (a1089 & c1089) | (b_inv1089 & c1089);
  wire s1090, sub1090, and1090, or1090;
  wire b_inv1090;
  assign b_inv1090 = ~b1090;
  assign s1090  = a1090 ^ b1090 ^ c1090;
  assign sub1090 = a1090 ^ b_inv1090 ^ c1090;
  assign and1090 = a1090 & b1090;
  assign or1090  = a1090 | b1090;
  assign c1091 = (a1090 & b1090) | (a1090 & c1090) | (b1090 & c1090);
  wire c_sub1091;
  assign c_sub1091 = (a1090 & b_inv1090) | (a1090 & c1090) | (b_inv1090 & c1090);
  wire s1091, sub1091, and1091, or1091;
  wire b_inv1091;
  assign b_inv1091 = ~b1091;
  assign s1091  = a1091 ^ b1091 ^ c1091;
  assign sub1091 = a1091 ^ b_inv1091 ^ c1091;
  assign and1091 = a1091 & b1091;
  assign or1091  = a1091 | b1091;
  assign c1092 = (a1091 & b1091) | (a1091 & c1091) | (b1091 & c1091);
  wire c_sub1092;
  assign c_sub1092 = (a1091 & b_inv1091) | (a1091 & c1091) | (b_inv1091 & c1091);
  wire s1092, sub1092, and1092, or1092;
  wire b_inv1092;
  assign b_inv1092 = ~b1092;
  assign s1092  = a1092 ^ b1092 ^ c1092;
  assign sub1092 = a1092 ^ b_inv1092 ^ c1092;
  assign and1092 = a1092 & b1092;
  assign or1092  = a1092 | b1092;
  assign c1093 = (a1092 & b1092) | (a1092 & c1092) | (b1092 & c1092);
  wire c_sub1093;
  assign c_sub1093 = (a1092 & b_inv1092) | (a1092 & c1092) | (b_inv1092 & c1092);
  wire s1093, sub1093, and1093, or1093;
  wire b_inv1093;
  assign b_inv1093 = ~b1093;
  assign s1093  = a1093 ^ b1093 ^ c1093;
  assign sub1093 = a1093 ^ b_inv1093 ^ c1093;
  assign and1093 = a1093 & b1093;
  assign or1093  = a1093 | b1093;
  assign c1094 = (a1093 & b1093) | (a1093 & c1093) | (b1093 & c1093);
  wire c_sub1094;
  assign c_sub1094 = (a1093 & b_inv1093) | (a1093 & c1093) | (b_inv1093 & c1093);
  wire s1094, sub1094, and1094, or1094;
  wire b_inv1094;
  assign b_inv1094 = ~b1094;
  assign s1094  = a1094 ^ b1094 ^ c1094;
  assign sub1094 = a1094 ^ b_inv1094 ^ c1094;
  assign and1094 = a1094 & b1094;
  assign or1094  = a1094 | b1094;
  assign c1095 = (a1094 & b1094) | (a1094 & c1094) | (b1094 & c1094);
  wire c_sub1095;
  assign c_sub1095 = (a1094 & b_inv1094) | (a1094 & c1094) | (b_inv1094 & c1094);
  wire s1095, sub1095, and1095, or1095;
  wire b_inv1095;
  assign b_inv1095 = ~b1095;
  assign s1095  = a1095 ^ b1095 ^ c1095;
  assign sub1095 = a1095 ^ b_inv1095 ^ c1095;
  assign and1095 = a1095 & b1095;
  assign or1095  = a1095 | b1095;
  assign c1096 = (a1095 & b1095) | (a1095 & c1095) | (b1095 & c1095);
  wire c_sub1096;
  assign c_sub1096 = (a1095 & b_inv1095) | (a1095 & c1095) | (b_inv1095 & c1095);
  wire s1096, sub1096, and1096, or1096;
  wire b_inv1096;
  assign b_inv1096 = ~b1096;
  assign s1096  = a1096 ^ b1096 ^ c1096;
  assign sub1096 = a1096 ^ b_inv1096 ^ c1096;
  assign and1096 = a1096 & b1096;
  assign or1096  = a1096 | b1096;
  assign c1097 = (a1096 & b1096) | (a1096 & c1096) | (b1096 & c1096);
  wire c_sub1097;
  assign c_sub1097 = (a1096 & b_inv1096) | (a1096 & c1096) | (b_inv1096 & c1096);
  wire s1097, sub1097, and1097, or1097;
  wire b_inv1097;
  assign b_inv1097 = ~b1097;
  assign s1097  = a1097 ^ b1097 ^ c1097;
  assign sub1097 = a1097 ^ b_inv1097 ^ c1097;
  assign and1097 = a1097 & b1097;
  assign or1097  = a1097 | b1097;
  assign c1098 = (a1097 & b1097) | (a1097 & c1097) | (b1097 & c1097);
  wire c_sub1098;
  assign c_sub1098 = (a1097 & b_inv1097) | (a1097 & c1097) | (b_inv1097 & c1097);
  wire s1098, sub1098, and1098, or1098;
  wire b_inv1098;
  assign b_inv1098 = ~b1098;
  assign s1098  = a1098 ^ b1098 ^ c1098;
  assign sub1098 = a1098 ^ b_inv1098 ^ c1098;
  assign and1098 = a1098 & b1098;
  assign or1098  = a1098 | b1098;
  assign c1099 = (a1098 & b1098) | (a1098 & c1098) | (b1098 & c1098);
  wire c_sub1099;
  assign c_sub1099 = (a1098 & b_inv1098) | (a1098 & c1098) | (b_inv1098 & c1098);
  wire s1099, sub1099, and1099, or1099;
  wire b_inv1099;
  assign b_inv1099 = ~b1099;
  assign s1099  = a1099 ^ b1099 ^ c1099;
  assign sub1099 = a1099 ^ b_inv1099 ^ c1099;
  assign and1099 = a1099 & b1099;
  assign or1099  = a1099 | b1099;
  assign c1100 = (a1099 & b1099) | (a1099 & c1099) | (b1099 & c1099);
  wire c_sub1100;
  assign c_sub1100 = (a1099 & b_inv1099) | (a1099 & c1099) | (b_inv1099 & c1099);
  wire s1100, sub1100, and1100, or1100;
  wire b_inv1100;
  assign b_inv1100 = ~b1100;
  assign s1100  = a1100 ^ b1100 ^ c1100;
  assign sub1100 = a1100 ^ b_inv1100 ^ c1100;
  assign and1100 = a1100 & b1100;
  assign or1100  = a1100 | b1100;
  assign c1101 = (a1100 & b1100) | (a1100 & c1100) | (b1100 & c1100);
  wire c_sub1101;
  assign c_sub1101 = (a1100 & b_inv1100) | (a1100 & c1100) | (b_inv1100 & c1100);
  wire s1101, sub1101, and1101, or1101;
  wire b_inv1101;
  assign b_inv1101 = ~b1101;
  assign s1101  = a1101 ^ b1101 ^ c1101;
  assign sub1101 = a1101 ^ b_inv1101 ^ c1101;
  assign and1101 = a1101 & b1101;
  assign or1101  = a1101 | b1101;
  assign c1102 = (a1101 & b1101) | (a1101 & c1101) | (b1101 & c1101);
  wire c_sub1102;
  assign c_sub1102 = (a1101 & b_inv1101) | (a1101 & c1101) | (b_inv1101 & c1101);
  wire s1102, sub1102, and1102, or1102;
  wire b_inv1102;
  assign b_inv1102 = ~b1102;
  assign s1102  = a1102 ^ b1102 ^ c1102;
  assign sub1102 = a1102 ^ b_inv1102 ^ c1102;
  assign and1102 = a1102 & b1102;
  assign or1102  = a1102 | b1102;
  assign c1103 = (a1102 & b1102) | (a1102 & c1102) | (b1102 & c1102);
  wire c_sub1103;
  assign c_sub1103 = (a1102 & b_inv1102) | (a1102 & c1102) | (b_inv1102 & c1102);
  wire s1103, sub1103, and1103, or1103;
  wire b_inv1103;
  assign b_inv1103 = ~b1103;
  assign s1103  = a1103 ^ b1103 ^ c1103;
  assign sub1103 = a1103 ^ b_inv1103 ^ c1103;
  assign and1103 = a1103 & b1103;
  assign or1103  = a1103 | b1103;
  assign c1104 = (a1103 & b1103) | (a1103 & c1103) | (b1103 & c1103);
  wire c_sub1104;
  assign c_sub1104 = (a1103 & b_inv1103) | (a1103 & c1103) | (b_inv1103 & c1103);
  wire s1104, sub1104, and1104, or1104;
  wire b_inv1104;
  assign b_inv1104 = ~b1104;
  assign s1104  = a1104 ^ b1104 ^ c1104;
  assign sub1104 = a1104 ^ b_inv1104 ^ c1104;
  assign and1104 = a1104 & b1104;
  assign or1104  = a1104 | b1104;
  assign c1105 = (a1104 & b1104) | (a1104 & c1104) | (b1104 & c1104);
  wire c_sub1105;
  assign c_sub1105 = (a1104 & b_inv1104) | (a1104 & c1104) | (b_inv1104 & c1104);
  wire s1105, sub1105, and1105, or1105;
  wire b_inv1105;
  assign b_inv1105 = ~b1105;
  assign s1105  = a1105 ^ b1105 ^ c1105;
  assign sub1105 = a1105 ^ b_inv1105 ^ c1105;
  assign and1105 = a1105 & b1105;
  assign or1105  = a1105 | b1105;
  assign c1106 = (a1105 & b1105) | (a1105 & c1105) | (b1105 & c1105);
  wire c_sub1106;
  assign c_sub1106 = (a1105 & b_inv1105) | (a1105 & c1105) | (b_inv1105 & c1105);
  wire s1106, sub1106, and1106, or1106;
  wire b_inv1106;
  assign b_inv1106 = ~b1106;
  assign s1106  = a1106 ^ b1106 ^ c1106;
  assign sub1106 = a1106 ^ b_inv1106 ^ c1106;
  assign and1106 = a1106 & b1106;
  assign or1106  = a1106 | b1106;
  assign c1107 = (a1106 & b1106) | (a1106 & c1106) | (b1106 & c1106);
  wire c_sub1107;
  assign c_sub1107 = (a1106 & b_inv1106) | (a1106 & c1106) | (b_inv1106 & c1106);
  wire s1107, sub1107, and1107, or1107;
  wire b_inv1107;
  assign b_inv1107 = ~b1107;
  assign s1107  = a1107 ^ b1107 ^ c1107;
  assign sub1107 = a1107 ^ b_inv1107 ^ c1107;
  assign and1107 = a1107 & b1107;
  assign or1107  = a1107 | b1107;
  assign c1108 = (a1107 & b1107) | (a1107 & c1107) | (b1107 & c1107);
  wire c_sub1108;
  assign c_sub1108 = (a1107 & b_inv1107) | (a1107 & c1107) | (b_inv1107 & c1107);
  wire s1108, sub1108, and1108, or1108;
  wire b_inv1108;
  assign b_inv1108 = ~b1108;
  assign s1108  = a1108 ^ b1108 ^ c1108;
  assign sub1108 = a1108 ^ b_inv1108 ^ c1108;
  assign and1108 = a1108 & b1108;
  assign or1108  = a1108 | b1108;
  assign c1109 = (a1108 & b1108) | (a1108 & c1108) | (b1108 & c1108);
  wire c_sub1109;
  assign c_sub1109 = (a1108 & b_inv1108) | (a1108 & c1108) | (b_inv1108 & c1108);
  wire s1109, sub1109, and1109, or1109;
  wire b_inv1109;
  assign b_inv1109 = ~b1109;
  assign s1109  = a1109 ^ b1109 ^ c1109;
  assign sub1109 = a1109 ^ b_inv1109 ^ c1109;
  assign and1109 = a1109 & b1109;
  assign or1109  = a1109 | b1109;
  assign c1110 = (a1109 & b1109) | (a1109 & c1109) | (b1109 & c1109);
  wire c_sub1110;
  assign c_sub1110 = (a1109 & b_inv1109) | (a1109 & c1109) | (b_inv1109 & c1109);
  wire s1110, sub1110, and1110, or1110;
  wire b_inv1110;
  assign b_inv1110 = ~b1110;
  assign s1110  = a1110 ^ b1110 ^ c1110;
  assign sub1110 = a1110 ^ b_inv1110 ^ c1110;
  assign and1110 = a1110 & b1110;
  assign or1110  = a1110 | b1110;
  assign c1111 = (a1110 & b1110) | (a1110 & c1110) | (b1110 & c1110);
  wire c_sub1111;
  assign c_sub1111 = (a1110 & b_inv1110) | (a1110 & c1110) | (b_inv1110 & c1110);
  wire s1111, sub1111, and1111, or1111;
  wire b_inv1111;
  assign b_inv1111 = ~b1111;
  assign s1111  = a1111 ^ b1111 ^ c1111;
  assign sub1111 = a1111 ^ b_inv1111 ^ c1111;
  assign and1111 = a1111 & b1111;
  assign or1111  = a1111 | b1111;
  assign c1112 = (a1111 & b1111) | (a1111 & c1111) | (b1111 & c1111);
  wire c_sub1112;
  assign c_sub1112 = (a1111 & b_inv1111) | (a1111 & c1111) | (b_inv1111 & c1111);
  wire s1112, sub1112, and1112, or1112;
  wire b_inv1112;
  assign b_inv1112 = ~b1112;
  assign s1112  = a1112 ^ b1112 ^ c1112;
  assign sub1112 = a1112 ^ b_inv1112 ^ c1112;
  assign and1112 = a1112 & b1112;
  assign or1112  = a1112 | b1112;
  assign c1113 = (a1112 & b1112) | (a1112 & c1112) | (b1112 & c1112);
  wire c_sub1113;
  assign c_sub1113 = (a1112 & b_inv1112) | (a1112 & c1112) | (b_inv1112 & c1112);
  wire s1113, sub1113, and1113, or1113;
  wire b_inv1113;
  assign b_inv1113 = ~b1113;
  assign s1113  = a1113 ^ b1113 ^ c1113;
  assign sub1113 = a1113 ^ b_inv1113 ^ c1113;
  assign and1113 = a1113 & b1113;
  assign or1113  = a1113 | b1113;
  assign c1114 = (a1113 & b1113) | (a1113 & c1113) | (b1113 & c1113);
  wire c_sub1114;
  assign c_sub1114 = (a1113 & b_inv1113) | (a1113 & c1113) | (b_inv1113 & c1113);
  wire s1114, sub1114, and1114, or1114;
  wire b_inv1114;
  assign b_inv1114 = ~b1114;
  assign s1114  = a1114 ^ b1114 ^ c1114;
  assign sub1114 = a1114 ^ b_inv1114 ^ c1114;
  assign and1114 = a1114 & b1114;
  assign or1114  = a1114 | b1114;
  assign c1115 = (a1114 & b1114) | (a1114 & c1114) | (b1114 & c1114);
  wire c_sub1115;
  assign c_sub1115 = (a1114 & b_inv1114) | (a1114 & c1114) | (b_inv1114 & c1114);
  wire s1115, sub1115, and1115, or1115;
  wire b_inv1115;
  assign b_inv1115 = ~b1115;
  assign s1115  = a1115 ^ b1115 ^ c1115;
  assign sub1115 = a1115 ^ b_inv1115 ^ c1115;
  assign and1115 = a1115 & b1115;
  assign or1115  = a1115 | b1115;
  assign c1116 = (a1115 & b1115) | (a1115 & c1115) | (b1115 & c1115);
  wire c_sub1116;
  assign c_sub1116 = (a1115 & b_inv1115) | (a1115 & c1115) | (b_inv1115 & c1115);
  wire s1116, sub1116, and1116, or1116;
  wire b_inv1116;
  assign b_inv1116 = ~b1116;
  assign s1116  = a1116 ^ b1116 ^ c1116;
  assign sub1116 = a1116 ^ b_inv1116 ^ c1116;
  assign and1116 = a1116 & b1116;
  assign or1116  = a1116 | b1116;
  assign c1117 = (a1116 & b1116) | (a1116 & c1116) | (b1116 & c1116);
  wire c_sub1117;
  assign c_sub1117 = (a1116 & b_inv1116) | (a1116 & c1116) | (b_inv1116 & c1116);
  wire s1117, sub1117, and1117, or1117;
  wire b_inv1117;
  assign b_inv1117 = ~b1117;
  assign s1117  = a1117 ^ b1117 ^ c1117;
  assign sub1117 = a1117 ^ b_inv1117 ^ c1117;
  assign and1117 = a1117 & b1117;
  assign or1117  = a1117 | b1117;
  assign c1118 = (a1117 & b1117) | (a1117 & c1117) | (b1117 & c1117);
  wire c_sub1118;
  assign c_sub1118 = (a1117 & b_inv1117) | (a1117 & c1117) | (b_inv1117 & c1117);
  wire s1118, sub1118, and1118, or1118;
  wire b_inv1118;
  assign b_inv1118 = ~b1118;
  assign s1118  = a1118 ^ b1118 ^ c1118;
  assign sub1118 = a1118 ^ b_inv1118 ^ c1118;
  assign and1118 = a1118 & b1118;
  assign or1118  = a1118 | b1118;
  assign c1119 = (a1118 & b1118) | (a1118 & c1118) | (b1118 & c1118);
  wire c_sub1119;
  assign c_sub1119 = (a1118 & b_inv1118) | (a1118 & c1118) | (b_inv1118 & c1118);
  wire s1119, sub1119, and1119, or1119;
  wire b_inv1119;
  assign b_inv1119 = ~b1119;
  assign s1119  = a1119 ^ b1119 ^ c1119;
  assign sub1119 = a1119 ^ b_inv1119 ^ c1119;
  assign and1119 = a1119 & b1119;
  assign or1119  = a1119 | b1119;
  assign c1120 = (a1119 & b1119) | (a1119 & c1119) | (b1119 & c1119);
  wire c_sub1120;
  assign c_sub1120 = (a1119 & b_inv1119) | (a1119 & c1119) | (b_inv1119 & c1119);
  wire s1120, sub1120, and1120, or1120;
  wire b_inv1120;
  assign b_inv1120 = ~b1120;
  assign s1120  = a1120 ^ b1120 ^ c1120;
  assign sub1120 = a1120 ^ b_inv1120 ^ c1120;
  assign and1120 = a1120 & b1120;
  assign or1120  = a1120 | b1120;
  assign c1121 = (a1120 & b1120) | (a1120 & c1120) | (b1120 & c1120);
  wire c_sub1121;
  assign c_sub1121 = (a1120 & b_inv1120) | (a1120 & c1120) | (b_inv1120 & c1120);
  wire s1121, sub1121, and1121, or1121;
  wire b_inv1121;
  assign b_inv1121 = ~b1121;
  assign s1121  = a1121 ^ b1121 ^ c1121;
  assign sub1121 = a1121 ^ b_inv1121 ^ c1121;
  assign and1121 = a1121 & b1121;
  assign or1121  = a1121 | b1121;
  assign c1122 = (a1121 & b1121) | (a1121 & c1121) | (b1121 & c1121);
  wire c_sub1122;
  assign c_sub1122 = (a1121 & b_inv1121) | (a1121 & c1121) | (b_inv1121 & c1121);
  wire s1122, sub1122, and1122, or1122;
  wire b_inv1122;
  assign b_inv1122 = ~b1122;
  assign s1122  = a1122 ^ b1122 ^ c1122;
  assign sub1122 = a1122 ^ b_inv1122 ^ c1122;
  assign and1122 = a1122 & b1122;
  assign or1122  = a1122 | b1122;
  assign c1123 = (a1122 & b1122) | (a1122 & c1122) | (b1122 & c1122);
  wire c_sub1123;
  assign c_sub1123 = (a1122 & b_inv1122) | (a1122 & c1122) | (b_inv1122 & c1122);
  wire s1123, sub1123, and1123, or1123;
  wire b_inv1123;
  assign b_inv1123 = ~b1123;
  assign s1123  = a1123 ^ b1123 ^ c1123;
  assign sub1123 = a1123 ^ b_inv1123 ^ c1123;
  assign and1123 = a1123 & b1123;
  assign or1123  = a1123 | b1123;
  assign c1124 = (a1123 & b1123) | (a1123 & c1123) | (b1123 & c1123);
  wire c_sub1124;
  assign c_sub1124 = (a1123 & b_inv1123) | (a1123 & c1123) | (b_inv1123 & c1123);
  wire s1124, sub1124, and1124, or1124;
  wire b_inv1124;
  assign b_inv1124 = ~b1124;
  assign s1124  = a1124 ^ b1124 ^ c1124;
  assign sub1124 = a1124 ^ b_inv1124 ^ c1124;
  assign and1124 = a1124 & b1124;
  assign or1124  = a1124 | b1124;
  assign c1125 = (a1124 & b1124) | (a1124 & c1124) | (b1124 & c1124);
  wire c_sub1125;
  assign c_sub1125 = (a1124 & b_inv1124) | (a1124 & c1124) | (b_inv1124 & c1124);
  wire s1125, sub1125, and1125, or1125;
  wire b_inv1125;
  assign b_inv1125 = ~b1125;
  assign s1125  = a1125 ^ b1125 ^ c1125;
  assign sub1125 = a1125 ^ b_inv1125 ^ c1125;
  assign and1125 = a1125 & b1125;
  assign or1125  = a1125 | b1125;
  assign c1126 = (a1125 & b1125) | (a1125 & c1125) | (b1125 & c1125);
  wire c_sub1126;
  assign c_sub1126 = (a1125 & b_inv1125) | (a1125 & c1125) | (b_inv1125 & c1125);
  wire s1126, sub1126, and1126, or1126;
  wire b_inv1126;
  assign b_inv1126 = ~b1126;
  assign s1126  = a1126 ^ b1126 ^ c1126;
  assign sub1126 = a1126 ^ b_inv1126 ^ c1126;
  assign and1126 = a1126 & b1126;
  assign or1126  = a1126 | b1126;
  assign c1127 = (a1126 & b1126) | (a1126 & c1126) | (b1126 & c1126);
  wire c_sub1127;
  assign c_sub1127 = (a1126 & b_inv1126) | (a1126 & c1126) | (b_inv1126 & c1126);
  wire s1127, sub1127, and1127, or1127;
  wire b_inv1127;
  assign b_inv1127 = ~b1127;
  assign s1127  = a1127 ^ b1127 ^ c1127;
  assign sub1127 = a1127 ^ b_inv1127 ^ c1127;
  assign and1127 = a1127 & b1127;
  assign or1127  = a1127 | b1127;
  assign c1128 = (a1127 & b1127) | (a1127 & c1127) | (b1127 & c1127);
  wire c_sub1128;
  assign c_sub1128 = (a1127 & b_inv1127) | (a1127 & c1127) | (b_inv1127 & c1127);
  wire s1128, sub1128, and1128, or1128;
  wire b_inv1128;
  assign b_inv1128 = ~b1128;
  assign s1128  = a1128 ^ b1128 ^ c1128;
  assign sub1128 = a1128 ^ b_inv1128 ^ c1128;
  assign and1128 = a1128 & b1128;
  assign or1128  = a1128 | b1128;
  assign c1129 = (a1128 & b1128) | (a1128 & c1128) | (b1128 & c1128);
  wire c_sub1129;
  assign c_sub1129 = (a1128 & b_inv1128) | (a1128 & c1128) | (b_inv1128 & c1128);
  wire s1129, sub1129, and1129, or1129;
  wire b_inv1129;
  assign b_inv1129 = ~b1129;
  assign s1129  = a1129 ^ b1129 ^ c1129;
  assign sub1129 = a1129 ^ b_inv1129 ^ c1129;
  assign and1129 = a1129 & b1129;
  assign or1129  = a1129 | b1129;
  assign c1130 = (a1129 & b1129) | (a1129 & c1129) | (b1129 & c1129);
  wire c_sub1130;
  assign c_sub1130 = (a1129 & b_inv1129) | (a1129 & c1129) | (b_inv1129 & c1129);
  wire s1130, sub1130, and1130, or1130;
  wire b_inv1130;
  assign b_inv1130 = ~b1130;
  assign s1130  = a1130 ^ b1130 ^ c1130;
  assign sub1130 = a1130 ^ b_inv1130 ^ c1130;
  assign and1130 = a1130 & b1130;
  assign or1130  = a1130 | b1130;
  assign c1131 = (a1130 & b1130) | (a1130 & c1130) | (b1130 & c1130);
  wire c_sub1131;
  assign c_sub1131 = (a1130 & b_inv1130) | (a1130 & c1130) | (b_inv1130 & c1130);
  wire s1131, sub1131, and1131, or1131;
  wire b_inv1131;
  assign b_inv1131 = ~b1131;
  assign s1131  = a1131 ^ b1131 ^ c1131;
  assign sub1131 = a1131 ^ b_inv1131 ^ c1131;
  assign and1131 = a1131 & b1131;
  assign or1131  = a1131 | b1131;
  assign c1132 = (a1131 & b1131) | (a1131 & c1131) | (b1131 & c1131);
  wire c_sub1132;
  assign c_sub1132 = (a1131 & b_inv1131) | (a1131 & c1131) | (b_inv1131 & c1131);
  wire s1132, sub1132, and1132, or1132;
  wire b_inv1132;
  assign b_inv1132 = ~b1132;
  assign s1132  = a1132 ^ b1132 ^ c1132;
  assign sub1132 = a1132 ^ b_inv1132 ^ c1132;
  assign and1132 = a1132 & b1132;
  assign or1132  = a1132 | b1132;
  assign c1133 = (a1132 & b1132) | (a1132 & c1132) | (b1132 & c1132);
  wire c_sub1133;
  assign c_sub1133 = (a1132 & b_inv1132) | (a1132 & c1132) | (b_inv1132 & c1132);
  wire s1133, sub1133, and1133, or1133;
  wire b_inv1133;
  assign b_inv1133 = ~b1133;
  assign s1133  = a1133 ^ b1133 ^ c1133;
  assign sub1133 = a1133 ^ b_inv1133 ^ c1133;
  assign and1133 = a1133 & b1133;
  assign or1133  = a1133 | b1133;
  assign c1134 = (a1133 & b1133) | (a1133 & c1133) | (b1133 & c1133);
  wire c_sub1134;
  assign c_sub1134 = (a1133 & b_inv1133) | (a1133 & c1133) | (b_inv1133 & c1133);
  wire s1134, sub1134, and1134, or1134;
  wire b_inv1134;
  assign b_inv1134 = ~b1134;
  assign s1134  = a1134 ^ b1134 ^ c1134;
  assign sub1134 = a1134 ^ b_inv1134 ^ c1134;
  assign and1134 = a1134 & b1134;
  assign or1134  = a1134 | b1134;
  assign c1135 = (a1134 & b1134) | (a1134 & c1134) | (b1134 & c1134);
  wire c_sub1135;
  assign c_sub1135 = (a1134 & b_inv1134) | (a1134 & c1134) | (b_inv1134 & c1134);
  wire s1135, sub1135, and1135, or1135;
  wire b_inv1135;
  assign b_inv1135 = ~b1135;
  assign s1135  = a1135 ^ b1135 ^ c1135;
  assign sub1135 = a1135 ^ b_inv1135 ^ c1135;
  assign and1135 = a1135 & b1135;
  assign or1135  = a1135 | b1135;
  assign c1136 = (a1135 & b1135) | (a1135 & c1135) | (b1135 & c1135);
  wire c_sub1136;
  assign c_sub1136 = (a1135 & b_inv1135) | (a1135 & c1135) | (b_inv1135 & c1135);
  wire s1136, sub1136, and1136, or1136;
  wire b_inv1136;
  assign b_inv1136 = ~b1136;
  assign s1136  = a1136 ^ b1136 ^ c1136;
  assign sub1136 = a1136 ^ b_inv1136 ^ c1136;
  assign and1136 = a1136 & b1136;
  assign or1136  = a1136 | b1136;
  assign c1137 = (a1136 & b1136) | (a1136 & c1136) | (b1136 & c1136);
  wire c_sub1137;
  assign c_sub1137 = (a1136 & b_inv1136) | (a1136 & c1136) | (b_inv1136 & c1136);
  wire s1137, sub1137, and1137, or1137;
  wire b_inv1137;
  assign b_inv1137 = ~b1137;
  assign s1137  = a1137 ^ b1137 ^ c1137;
  assign sub1137 = a1137 ^ b_inv1137 ^ c1137;
  assign and1137 = a1137 & b1137;
  assign or1137  = a1137 | b1137;
  assign c1138 = (a1137 & b1137) | (a1137 & c1137) | (b1137 & c1137);
  wire c_sub1138;
  assign c_sub1138 = (a1137 & b_inv1137) | (a1137 & c1137) | (b_inv1137 & c1137);
  wire s1138, sub1138, and1138, or1138;
  wire b_inv1138;
  assign b_inv1138 = ~b1138;
  assign s1138  = a1138 ^ b1138 ^ c1138;
  assign sub1138 = a1138 ^ b_inv1138 ^ c1138;
  assign and1138 = a1138 & b1138;
  assign or1138  = a1138 | b1138;
  assign c1139 = (a1138 & b1138) | (a1138 & c1138) | (b1138 & c1138);
  wire c_sub1139;
  assign c_sub1139 = (a1138 & b_inv1138) | (a1138 & c1138) | (b_inv1138 & c1138);
  wire s1139, sub1139, and1139, or1139;
  wire b_inv1139;
  assign b_inv1139 = ~b1139;
  assign s1139  = a1139 ^ b1139 ^ c1139;
  assign sub1139 = a1139 ^ b_inv1139 ^ c1139;
  assign and1139 = a1139 & b1139;
  assign or1139  = a1139 | b1139;
  assign c1140 = (a1139 & b1139) | (a1139 & c1139) | (b1139 & c1139);
  wire c_sub1140;
  assign c_sub1140 = (a1139 & b_inv1139) | (a1139 & c1139) | (b_inv1139 & c1139);
  wire s1140, sub1140, and1140, or1140;
  wire b_inv1140;
  assign b_inv1140 = ~b1140;
  assign s1140  = a1140 ^ b1140 ^ c1140;
  assign sub1140 = a1140 ^ b_inv1140 ^ c1140;
  assign and1140 = a1140 & b1140;
  assign or1140  = a1140 | b1140;
  assign c1141 = (a1140 & b1140) | (a1140 & c1140) | (b1140 & c1140);
  wire c_sub1141;
  assign c_sub1141 = (a1140 & b_inv1140) | (a1140 & c1140) | (b_inv1140 & c1140);
  wire s1141, sub1141, and1141, or1141;
  wire b_inv1141;
  assign b_inv1141 = ~b1141;
  assign s1141  = a1141 ^ b1141 ^ c1141;
  assign sub1141 = a1141 ^ b_inv1141 ^ c1141;
  assign and1141 = a1141 & b1141;
  assign or1141  = a1141 | b1141;
  assign c1142 = (a1141 & b1141) | (a1141 & c1141) | (b1141 & c1141);
  wire c_sub1142;
  assign c_sub1142 = (a1141 & b_inv1141) | (a1141 & c1141) | (b_inv1141 & c1141);
  wire s1142, sub1142, and1142, or1142;
  wire b_inv1142;
  assign b_inv1142 = ~b1142;
  assign s1142  = a1142 ^ b1142 ^ c1142;
  assign sub1142 = a1142 ^ b_inv1142 ^ c1142;
  assign and1142 = a1142 & b1142;
  assign or1142  = a1142 | b1142;
  assign c1143 = (a1142 & b1142) | (a1142 & c1142) | (b1142 & c1142);
  wire c_sub1143;
  assign c_sub1143 = (a1142 & b_inv1142) | (a1142 & c1142) | (b_inv1142 & c1142);
  wire s1143, sub1143, and1143, or1143;
  wire b_inv1143;
  assign b_inv1143 = ~b1143;
  assign s1143  = a1143 ^ b1143 ^ c1143;
  assign sub1143 = a1143 ^ b_inv1143 ^ c1143;
  assign and1143 = a1143 & b1143;
  assign or1143  = a1143 | b1143;
  assign c1144 = (a1143 & b1143) | (a1143 & c1143) | (b1143 & c1143);
  wire c_sub1144;
  assign c_sub1144 = (a1143 & b_inv1143) | (a1143 & c1143) | (b_inv1143 & c1143);
  wire s1144, sub1144, and1144, or1144;
  wire b_inv1144;
  assign b_inv1144 = ~b1144;
  assign s1144  = a1144 ^ b1144 ^ c1144;
  assign sub1144 = a1144 ^ b_inv1144 ^ c1144;
  assign and1144 = a1144 & b1144;
  assign or1144  = a1144 | b1144;
  assign c1145 = (a1144 & b1144) | (a1144 & c1144) | (b1144 & c1144);
  wire c_sub1145;
  assign c_sub1145 = (a1144 & b_inv1144) | (a1144 & c1144) | (b_inv1144 & c1144);
  wire s1145, sub1145, and1145, or1145;
  wire b_inv1145;
  assign b_inv1145 = ~b1145;
  assign s1145  = a1145 ^ b1145 ^ c1145;
  assign sub1145 = a1145 ^ b_inv1145 ^ c1145;
  assign and1145 = a1145 & b1145;
  assign or1145  = a1145 | b1145;
  assign c1146 = (a1145 & b1145) | (a1145 & c1145) | (b1145 & c1145);
  wire c_sub1146;
  assign c_sub1146 = (a1145 & b_inv1145) | (a1145 & c1145) | (b_inv1145 & c1145);
  wire s1146, sub1146, and1146, or1146;
  wire b_inv1146;
  assign b_inv1146 = ~b1146;
  assign s1146  = a1146 ^ b1146 ^ c1146;
  assign sub1146 = a1146 ^ b_inv1146 ^ c1146;
  assign and1146 = a1146 & b1146;
  assign or1146  = a1146 | b1146;
  assign c1147 = (a1146 & b1146) | (a1146 & c1146) | (b1146 & c1146);
  wire c_sub1147;
  assign c_sub1147 = (a1146 & b_inv1146) | (a1146 & c1146) | (b_inv1146 & c1146);
  wire s1147, sub1147, and1147, or1147;
  wire b_inv1147;
  assign b_inv1147 = ~b1147;
  assign s1147  = a1147 ^ b1147 ^ c1147;
  assign sub1147 = a1147 ^ b_inv1147 ^ c1147;
  assign and1147 = a1147 & b1147;
  assign or1147  = a1147 | b1147;
  assign c1148 = (a1147 & b1147) | (a1147 & c1147) | (b1147 & c1147);
  wire c_sub1148;
  assign c_sub1148 = (a1147 & b_inv1147) | (a1147 & c1147) | (b_inv1147 & c1147);
  wire s1148, sub1148, and1148, or1148;
  wire b_inv1148;
  assign b_inv1148 = ~b1148;
  assign s1148  = a1148 ^ b1148 ^ c1148;
  assign sub1148 = a1148 ^ b_inv1148 ^ c1148;
  assign and1148 = a1148 & b1148;
  assign or1148  = a1148 | b1148;
  assign c1149 = (a1148 & b1148) | (a1148 & c1148) | (b1148 & c1148);
  wire c_sub1149;
  assign c_sub1149 = (a1148 & b_inv1148) | (a1148 & c1148) | (b_inv1148 & c1148);
  wire s1149, sub1149, and1149, or1149;
  wire b_inv1149;
  assign b_inv1149 = ~b1149;
  assign s1149  = a1149 ^ b1149 ^ c1149;
  assign sub1149 = a1149 ^ b_inv1149 ^ c1149;
  assign and1149 = a1149 & b1149;
  assign or1149  = a1149 | b1149;
  assign c1150 = (a1149 & b1149) | (a1149 & c1149) | (b1149 & c1149);
  wire c_sub1150;
  assign c_sub1150 = (a1149 & b_inv1149) | (a1149 & c1149) | (b_inv1149 & c1149);
  wire s1150, sub1150, and1150, or1150;
  wire b_inv1150;
  assign b_inv1150 = ~b1150;
  assign s1150  = a1150 ^ b1150 ^ c1150;
  assign sub1150 = a1150 ^ b_inv1150 ^ c1150;
  assign and1150 = a1150 & b1150;
  assign or1150  = a1150 | b1150;
  assign c1151 = (a1150 & b1150) | (a1150 & c1150) | (b1150 & c1150);
  wire c_sub1151;
  assign c_sub1151 = (a1150 & b_inv1150) | (a1150 & c1150) | (b_inv1150 & c1150);
  wire s1151, sub1151, and1151, or1151;
  wire b_inv1151;
  assign b_inv1151 = ~b1151;
  assign s1151  = a1151 ^ b1151 ^ c1151;
  assign sub1151 = a1151 ^ b_inv1151 ^ c1151;
  assign and1151 = a1151 & b1151;
  assign or1151  = a1151 | b1151;
  assign c1152 = (a1151 & b1151) | (a1151 & c1151) | (b1151 & c1151);
  wire c_sub1152;
  assign c_sub1152 = (a1151 & b_inv1151) | (a1151 & c1151) | (b_inv1151 & c1151);
  wire s1152, sub1152, and1152, or1152;
  wire b_inv1152;
  assign b_inv1152 = ~b1152;
  assign s1152  = a1152 ^ b1152 ^ c1152;
  assign sub1152 = a1152 ^ b_inv1152 ^ c1152;
  assign and1152 = a1152 & b1152;
  assign or1152  = a1152 | b1152;
  assign c1153 = (a1152 & b1152) | (a1152 & c1152) | (b1152 & c1152);
  wire c_sub1153;
  assign c_sub1153 = (a1152 & b_inv1152) | (a1152 & c1152) | (b_inv1152 & c1152);
  wire s1153, sub1153, and1153, or1153;
  wire b_inv1153;
  assign b_inv1153 = ~b1153;
  assign s1153  = a1153 ^ b1153 ^ c1153;
  assign sub1153 = a1153 ^ b_inv1153 ^ c1153;
  assign and1153 = a1153 & b1153;
  assign or1153  = a1153 | b1153;
  assign c1154 = (a1153 & b1153) | (a1153 & c1153) | (b1153 & c1153);
  wire c_sub1154;
  assign c_sub1154 = (a1153 & b_inv1153) | (a1153 & c1153) | (b_inv1153 & c1153);
  wire s1154, sub1154, and1154, or1154;
  wire b_inv1154;
  assign b_inv1154 = ~b1154;
  assign s1154  = a1154 ^ b1154 ^ c1154;
  assign sub1154 = a1154 ^ b_inv1154 ^ c1154;
  assign and1154 = a1154 & b1154;
  assign or1154  = a1154 | b1154;
  assign c1155 = (a1154 & b1154) | (a1154 & c1154) | (b1154 & c1154);
  wire c_sub1155;
  assign c_sub1155 = (a1154 & b_inv1154) | (a1154 & c1154) | (b_inv1154 & c1154);
  wire s1155, sub1155, and1155, or1155;
  wire b_inv1155;
  assign b_inv1155 = ~b1155;
  assign s1155  = a1155 ^ b1155 ^ c1155;
  assign sub1155 = a1155 ^ b_inv1155 ^ c1155;
  assign and1155 = a1155 & b1155;
  assign or1155  = a1155 | b1155;
  assign c1156 = (a1155 & b1155) | (a1155 & c1155) | (b1155 & c1155);
  wire c_sub1156;
  assign c_sub1156 = (a1155 & b_inv1155) | (a1155 & c1155) | (b_inv1155 & c1155);
  wire s1156, sub1156, and1156, or1156;
  wire b_inv1156;
  assign b_inv1156 = ~b1156;
  assign s1156  = a1156 ^ b1156 ^ c1156;
  assign sub1156 = a1156 ^ b_inv1156 ^ c1156;
  assign and1156 = a1156 & b1156;
  assign or1156  = a1156 | b1156;
  assign c1157 = (a1156 & b1156) | (a1156 & c1156) | (b1156 & c1156);
  wire c_sub1157;
  assign c_sub1157 = (a1156 & b_inv1156) | (a1156 & c1156) | (b_inv1156 & c1156);
  wire s1157, sub1157, and1157, or1157;
  wire b_inv1157;
  assign b_inv1157 = ~b1157;
  assign s1157  = a1157 ^ b1157 ^ c1157;
  assign sub1157 = a1157 ^ b_inv1157 ^ c1157;
  assign and1157 = a1157 & b1157;
  assign or1157  = a1157 | b1157;
  assign c1158 = (a1157 & b1157) | (a1157 & c1157) | (b1157 & c1157);
  wire c_sub1158;
  assign c_sub1158 = (a1157 & b_inv1157) | (a1157 & c1157) | (b_inv1157 & c1157);
  wire s1158, sub1158, and1158, or1158;
  wire b_inv1158;
  assign b_inv1158 = ~b1158;
  assign s1158  = a1158 ^ b1158 ^ c1158;
  assign sub1158 = a1158 ^ b_inv1158 ^ c1158;
  assign and1158 = a1158 & b1158;
  assign or1158  = a1158 | b1158;
  assign c1159 = (a1158 & b1158) | (a1158 & c1158) | (b1158 & c1158);
  wire c_sub1159;
  assign c_sub1159 = (a1158 & b_inv1158) | (a1158 & c1158) | (b_inv1158 & c1158);
  wire s1159, sub1159, and1159, or1159;
  wire b_inv1159;
  assign b_inv1159 = ~b1159;
  assign s1159  = a1159 ^ b1159 ^ c1159;
  assign sub1159 = a1159 ^ b_inv1159 ^ c1159;
  assign and1159 = a1159 & b1159;
  assign or1159  = a1159 | b1159;
  assign c1160 = (a1159 & b1159) | (a1159 & c1159) | (b1159 & c1159);
  wire c_sub1160;
  assign c_sub1160 = (a1159 & b_inv1159) | (a1159 & c1159) | (b_inv1159 & c1159);
  wire s1160, sub1160, and1160, or1160;
  wire b_inv1160;
  assign b_inv1160 = ~b1160;
  assign s1160  = a1160 ^ b1160 ^ c1160;
  assign sub1160 = a1160 ^ b_inv1160 ^ c1160;
  assign and1160 = a1160 & b1160;
  assign or1160  = a1160 | b1160;
  assign c1161 = (a1160 & b1160) | (a1160 & c1160) | (b1160 & c1160);
  wire c_sub1161;
  assign c_sub1161 = (a1160 & b_inv1160) | (a1160 & c1160) | (b_inv1160 & c1160);
  wire s1161, sub1161, and1161, or1161;
  wire b_inv1161;
  assign b_inv1161 = ~b1161;
  assign s1161  = a1161 ^ b1161 ^ c1161;
  assign sub1161 = a1161 ^ b_inv1161 ^ c1161;
  assign and1161 = a1161 & b1161;
  assign or1161  = a1161 | b1161;
  assign c1162 = (a1161 & b1161) | (a1161 & c1161) | (b1161 & c1161);
  wire c_sub1162;
  assign c_sub1162 = (a1161 & b_inv1161) | (a1161 & c1161) | (b_inv1161 & c1161);
  wire s1162, sub1162, and1162, or1162;
  wire b_inv1162;
  assign b_inv1162 = ~b1162;
  assign s1162  = a1162 ^ b1162 ^ c1162;
  assign sub1162 = a1162 ^ b_inv1162 ^ c1162;
  assign and1162 = a1162 & b1162;
  assign or1162  = a1162 | b1162;
  assign c1163 = (a1162 & b1162) | (a1162 & c1162) | (b1162 & c1162);
  wire c_sub1163;
  assign c_sub1163 = (a1162 & b_inv1162) | (a1162 & c1162) | (b_inv1162 & c1162);
  wire s1163, sub1163, and1163, or1163;
  wire b_inv1163;
  assign b_inv1163 = ~b1163;
  assign s1163  = a1163 ^ b1163 ^ c1163;
  assign sub1163 = a1163 ^ b_inv1163 ^ c1163;
  assign and1163 = a1163 & b1163;
  assign or1163  = a1163 | b1163;
  assign c1164 = (a1163 & b1163) | (a1163 & c1163) | (b1163 & c1163);
  wire c_sub1164;
  assign c_sub1164 = (a1163 & b_inv1163) | (a1163 & c1163) | (b_inv1163 & c1163);
  wire s1164, sub1164, and1164, or1164;
  wire b_inv1164;
  assign b_inv1164 = ~b1164;
  assign s1164  = a1164 ^ b1164 ^ c1164;
  assign sub1164 = a1164 ^ b_inv1164 ^ c1164;
  assign and1164 = a1164 & b1164;
  assign or1164  = a1164 | b1164;
  assign c1165 = (a1164 & b1164) | (a1164 & c1164) | (b1164 & c1164);
  wire c_sub1165;
  assign c_sub1165 = (a1164 & b_inv1164) | (a1164 & c1164) | (b_inv1164 & c1164);
  wire s1165, sub1165, and1165, or1165;
  wire b_inv1165;
  assign b_inv1165 = ~b1165;
  assign s1165  = a1165 ^ b1165 ^ c1165;
  assign sub1165 = a1165 ^ b_inv1165 ^ c1165;
  assign and1165 = a1165 & b1165;
  assign or1165  = a1165 | b1165;
  assign c1166 = (a1165 & b1165) | (a1165 & c1165) | (b1165 & c1165);
  wire c_sub1166;
  assign c_sub1166 = (a1165 & b_inv1165) | (a1165 & c1165) | (b_inv1165 & c1165);
  wire s1166, sub1166, and1166, or1166;
  wire b_inv1166;
  assign b_inv1166 = ~b1166;
  assign s1166  = a1166 ^ b1166 ^ c1166;
  assign sub1166 = a1166 ^ b_inv1166 ^ c1166;
  assign and1166 = a1166 & b1166;
  assign or1166  = a1166 | b1166;
  assign c1167 = (a1166 & b1166) | (a1166 & c1166) | (b1166 & c1166);
  wire c_sub1167;
  assign c_sub1167 = (a1166 & b_inv1166) | (a1166 & c1166) | (b_inv1166 & c1166);
  wire s1167, sub1167, and1167, or1167;
  wire b_inv1167;
  assign b_inv1167 = ~b1167;
  assign s1167  = a1167 ^ b1167 ^ c1167;
  assign sub1167 = a1167 ^ b_inv1167 ^ c1167;
  assign and1167 = a1167 & b1167;
  assign or1167  = a1167 | b1167;
  assign c1168 = (a1167 & b1167) | (a1167 & c1167) | (b1167 & c1167);
  wire c_sub1168;
  assign c_sub1168 = (a1167 & b_inv1167) | (a1167 & c1167) | (b_inv1167 & c1167);
  wire s1168, sub1168, and1168, or1168;
  wire b_inv1168;
  assign b_inv1168 = ~b1168;
  assign s1168  = a1168 ^ b1168 ^ c1168;
  assign sub1168 = a1168 ^ b_inv1168 ^ c1168;
  assign and1168 = a1168 & b1168;
  assign or1168  = a1168 | b1168;
  assign c1169 = (a1168 & b1168) | (a1168 & c1168) | (b1168 & c1168);
  wire c_sub1169;
  assign c_sub1169 = (a1168 & b_inv1168) | (a1168 & c1168) | (b_inv1168 & c1168);
  wire s1169, sub1169, and1169, or1169;
  wire b_inv1169;
  assign b_inv1169 = ~b1169;
  assign s1169  = a1169 ^ b1169 ^ c1169;
  assign sub1169 = a1169 ^ b_inv1169 ^ c1169;
  assign and1169 = a1169 & b1169;
  assign or1169  = a1169 | b1169;
  assign c1170 = (a1169 & b1169) | (a1169 & c1169) | (b1169 & c1169);
  wire c_sub1170;
  assign c_sub1170 = (a1169 & b_inv1169) | (a1169 & c1169) | (b_inv1169 & c1169);
  wire s1170, sub1170, and1170, or1170;
  wire b_inv1170;
  assign b_inv1170 = ~b1170;
  assign s1170  = a1170 ^ b1170 ^ c1170;
  assign sub1170 = a1170 ^ b_inv1170 ^ c1170;
  assign and1170 = a1170 & b1170;
  assign or1170  = a1170 | b1170;
  assign c1171 = (a1170 & b1170) | (a1170 & c1170) | (b1170 & c1170);
  wire c_sub1171;
  assign c_sub1171 = (a1170 & b_inv1170) | (a1170 & c1170) | (b_inv1170 & c1170);
  wire s1171, sub1171, and1171, or1171;
  wire b_inv1171;
  assign b_inv1171 = ~b1171;
  assign s1171  = a1171 ^ b1171 ^ c1171;
  assign sub1171 = a1171 ^ b_inv1171 ^ c1171;
  assign and1171 = a1171 & b1171;
  assign or1171  = a1171 | b1171;
  assign c1172 = (a1171 & b1171) | (a1171 & c1171) | (b1171 & c1171);
  wire c_sub1172;
  assign c_sub1172 = (a1171 & b_inv1171) | (a1171 & c1171) | (b_inv1171 & c1171);
  wire s1172, sub1172, and1172, or1172;
  wire b_inv1172;
  assign b_inv1172 = ~b1172;
  assign s1172  = a1172 ^ b1172 ^ c1172;
  assign sub1172 = a1172 ^ b_inv1172 ^ c1172;
  assign and1172 = a1172 & b1172;
  assign or1172  = a1172 | b1172;
  assign c1173 = (a1172 & b1172) | (a1172 & c1172) | (b1172 & c1172);
  wire c_sub1173;
  assign c_sub1173 = (a1172 & b_inv1172) | (a1172 & c1172) | (b_inv1172 & c1172);
  wire s1173, sub1173, and1173, or1173;
  wire b_inv1173;
  assign b_inv1173 = ~b1173;
  assign s1173  = a1173 ^ b1173 ^ c1173;
  assign sub1173 = a1173 ^ b_inv1173 ^ c1173;
  assign and1173 = a1173 & b1173;
  assign or1173  = a1173 | b1173;
  assign c1174 = (a1173 & b1173) | (a1173 & c1173) | (b1173 & c1173);
  wire c_sub1174;
  assign c_sub1174 = (a1173 & b_inv1173) | (a1173 & c1173) | (b_inv1173 & c1173);
  wire s1174, sub1174, and1174, or1174;
  wire b_inv1174;
  assign b_inv1174 = ~b1174;
  assign s1174  = a1174 ^ b1174 ^ c1174;
  assign sub1174 = a1174 ^ b_inv1174 ^ c1174;
  assign and1174 = a1174 & b1174;
  assign or1174  = a1174 | b1174;
  assign c1175 = (a1174 & b1174) | (a1174 & c1174) | (b1174 & c1174);
  wire c_sub1175;
  assign c_sub1175 = (a1174 & b_inv1174) | (a1174 & c1174) | (b_inv1174 & c1174);
  wire s1175, sub1175, and1175, or1175;
  wire b_inv1175;
  assign b_inv1175 = ~b1175;
  assign s1175  = a1175 ^ b1175 ^ c1175;
  assign sub1175 = a1175 ^ b_inv1175 ^ c1175;
  assign and1175 = a1175 & b1175;
  assign or1175  = a1175 | b1175;
  assign c1176 = (a1175 & b1175) | (a1175 & c1175) | (b1175 & c1175);
  wire c_sub1176;
  assign c_sub1176 = (a1175 & b_inv1175) | (a1175 & c1175) | (b_inv1175 & c1175);
  wire s1176, sub1176, and1176, or1176;
  wire b_inv1176;
  assign b_inv1176 = ~b1176;
  assign s1176  = a1176 ^ b1176 ^ c1176;
  assign sub1176 = a1176 ^ b_inv1176 ^ c1176;
  assign and1176 = a1176 & b1176;
  assign or1176  = a1176 | b1176;
  assign c1177 = (a1176 & b1176) | (a1176 & c1176) | (b1176 & c1176);
  wire c_sub1177;
  assign c_sub1177 = (a1176 & b_inv1176) | (a1176 & c1176) | (b_inv1176 & c1176);
  wire s1177, sub1177, and1177, or1177;
  wire b_inv1177;
  assign b_inv1177 = ~b1177;
  assign s1177  = a1177 ^ b1177 ^ c1177;
  assign sub1177 = a1177 ^ b_inv1177 ^ c1177;
  assign and1177 = a1177 & b1177;
  assign or1177  = a1177 | b1177;
  assign c1178 = (a1177 & b1177) | (a1177 & c1177) | (b1177 & c1177);
  wire c_sub1178;
  assign c_sub1178 = (a1177 & b_inv1177) | (a1177 & c1177) | (b_inv1177 & c1177);
  wire s1178, sub1178, and1178, or1178;
  wire b_inv1178;
  assign b_inv1178 = ~b1178;
  assign s1178  = a1178 ^ b1178 ^ c1178;
  assign sub1178 = a1178 ^ b_inv1178 ^ c1178;
  assign and1178 = a1178 & b1178;
  assign or1178  = a1178 | b1178;
  assign c1179 = (a1178 & b1178) | (a1178 & c1178) | (b1178 & c1178);
  wire c_sub1179;
  assign c_sub1179 = (a1178 & b_inv1178) | (a1178 & c1178) | (b_inv1178 & c1178);
  wire s1179, sub1179, and1179, or1179;
  wire b_inv1179;
  assign b_inv1179 = ~b1179;
  assign s1179  = a1179 ^ b1179 ^ c1179;
  assign sub1179 = a1179 ^ b_inv1179 ^ c1179;
  assign and1179 = a1179 & b1179;
  assign or1179  = a1179 | b1179;
  assign c1180 = (a1179 & b1179) | (a1179 & c1179) | (b1179 & c1179);
  wire c_sub1180;
  assign c_sub1180 = (a1179 & b_inv1179) | (a1179 & c1179) | (b_inv1179 & c1179);
  wire s1180, sub1180, and1180, or1180;
  wire b_inv1180;
  assign b_inv1180 = ~b1180;
  assign s1180  = a1180 ^ b1180 ^ c1180;
  assign sub1180 = a1180 ^ b_inv1180 ^ c1180;
  assign and1180 = a1180 & b1180;
  assign or1180  = a1180 | b1180;
  assign c1181 = (a1180 & b1180) | (a1180 & c1180) | (b1180 & c1180);
  wire c_sub1181;
  assign c_sub1181 = (a1180 & b_inv1180) | (a1180 & c1180) | (b_inv1180 & c1180);
  wire s1181, sub1181, and1181, or1181;
  wire b_inv1181;
  assign b_inv1181 = ~b1181;
  assign s1181  = a1181 ^ b1181 ^ c1181;
  assign sub1181 = a1181 ^ b_inv1181 ^ c1181;
  assign and1181 = a1181 & b1181;
  assign or1181  = a1181 | b1181;
  assign c1182 = (a1181 & b1181) | (a1181 & c1181) | (b1181 & c1181);
  wire c_sub1182;
  assign c_sub1182 = (a1181 & b_inv1181) | (a1181 & c1181) | (b_inv1181 & c1181);
  wire s1182, sub1182, and1182, or1182;
  wire b_inv1182;
  assign b_inv1182 = ~b1182;
  assign s1182  = a1182 ^ b1182 ^ c1182;
  assign sub1182 = a1182 ^ b_inv1182 ^ c1182;
  assign and1182 = a1182 & b1182;
  assign or1182  = a1182 | b1182;
  assign c1183 = (a1182 & b1182) | (a1182 & c1182) | (b1182 & c1182);
  wire c_sub1183;
  assign c_sub1183 = (a1182 & b_inv1182) | (a1182 & c1182) | (b_inv1182 & c1182);
  wire s1183, sub1183, and1183, or1183;
  wire b_inv1183;
  assign b_inv1183 = ~b1183;
  assign s1183  = a1183 ^ b1183 ^ c1183;
  assign sub1183 = a1183 ^ b_inv1183 ^ c1183;
  assign and1183 = a1183 & b1183;
  assign or1183  = a1183 | b1183;
  assign c1184 = (a1183 & b1183) | (a1183 & c1183) | (b1183 & c1183);
  wire c_sub1184;
  assign c_sub1184 = (a1183 & b_inv1183) | (a1183 & c1183) | (b_inv1183 & c1183);
  wire s1184, sub1184, and1184, or1184;
  wire b_inv1184;
  assign b_inv1184 = ~b1184;
  assign s1184  = a1184 ^ b1184 ^ c1184;
  assign sub1184 = a1184 ^ b_inv1184 ^ c1184;
  assign and1184 = a1184 & b1184;
  assign or1184  = a1184 | b1184;
  assign c1185 = (a1184 & b1184) | (a1184 & c1184) | (b1184 & c1184);
  wire c_sub1185;
  assign c_sub1185 = (a1184 & b_inv1184) | (a1184 & c1184) | (b_inv1184 & c1184);
  wire s1185, sub1185, and1185, or1185;
  wire b_inv1185;
  assign b_inv1185 = ~b1185;
  assign s1185  = a1185 ^ b1185 ^ c1185;
  assign sub1185 = a1185 ^ b_inv1185 ^ c1185;
  assign and1185 = a1185 & b1185;
  assign or1185  = a1185 | b1185;
  assign c1186 = (a1185 & b1185) | (a1185 & c1185) | (b1185 & c1185);
  wire c_sub1186;
  assign c_sub1186 = (a1185 & b_inv1185) | (a1185 & c1185) | (b_inv1185 & c1185);
  wire s1186, sub1186, and1186, or1186;
  wire b_inv1186;
  assign b_inv1186 = ~b1186;
  assign s1186  = a1186 ^ b1186 ^ c1186;
  assign sub1186 = a1186 ^ b_inv1186 ^ c1186;
  assign and1186 = a1186 & b1186;
  assign or1186  = a1186 | b1186;
  assign c1187 = (a1186 & b1186) | (a1186 & c1186) | (b1186 & c1186);
  wire c_sub1187;
  assign c_sub1187 = (a1186 & b_inv1186) | (a1186 & c1186) | (b_inv1186 & c1186);
  wire s1187, sub1187, and1187, or1187;
  wire b_inv1187;
  assign b_inv1187 = ~b1187;
  assign s1187  = a1187 ^ b1187 ^ c1187;
  assign sub1187 = a1187 ^ b_inv1187 ^ c1187;
  assign and1187 = a1187 & b1187;
  assign or1187  = a1187 | b1187;
  assign c1188 = (a1187 & b1187) | (a1187 & c1187) | (b1187 & c1187);
  wire c_sub1188;
  assign c_sub1188 = (a1187 & b_inv1187) | (a1187 & c1187) | (b_inv1187 & c1187);
  wire s1188, sub1188, and1188, or1188;
  wire b_inv1188;
  assign b_inv1188 = ~b1188;
  assign s1188  = a1188 ^ b1188 ^ c1188;
  assign sub1188 = a1188 ^ b_inv1188 ^ c1188;
  assign and1188 = a1188 & b1188;
  assign or1188  = a1188 | b1188;
  assign c1189 = (a1188 & b1188) | (a1188 & c1188) | (b1188 & c1188);
  wire c_sub1189;
  assign c_sub1189 = (a1188 & b_inv1188) | (a1188 & c1188) | (b_inv1188 & c1188);
  wire s1189, sub1189, and1189, or1189;
  wire b_inv1189;
  assign b_inv1189 = ~b1189;
  assign s1189  = a1189 ^ b1189 ^ c1189;
  assign sub1189 = a1189 ^ b_inv1189 ^ c1189;
  assign and1189 = a1189 & b1189;
  assign or1189  = a1189 | b1189;
  assign c1190 = (a1189 & b1189) | (a1189 & c1189) | (b1189 & c1189);
  wire c_sub1190;
  assign c_sub1190 = (a1189 & b_inv1189) | (a1189 & c1189) | (b_inv1189 & c1189);
  wire s1190, sub1190, and1190, or1190;
  wire b_inv1190;
  assign b_inv1190 = ~b1190;
  assign s1190  = a1190 ^ b1190 ^ c1190;
  assign sub1190 = a1190 ^ b_inv1190 ^ c1190;
  assign and1190 = a1190 & b1190;
  assign or1190  = a1190 | b1190;
  assign c1191 = (a1190 & b1190) | (a1190 & c1190) | (b1190 & c1190);
  wire c_sub1191;
  assign c_sub1191 = (a1190 & b_inv1190) | (a1190 & c1190) | (b_inv1190 & c1190);
  wire s1191, sub1191, and1191, or1191;
  wire b_inv1191;
  assign b_inv1191 = ~b1191;
  assign s1191  = a1191 ^ b1191 ^ c1191;
  assign sub1191 = a1191 ^ b_inv1191 ^ c1191;
  assign and1191 = a1191 & b1191;
  assign or1191  = a1191 | b1191;
  assign c1192 = (a1191 & b1191) | (a1191 & c1191) | (b1191 & c1191);
  wire c_sub1192;
  assign c_sub1192 = (a1191 & b_inv1191) | (a1191 & c1191) | (b_inv1191 & c1191);
  wire s1192, sub1192, and1192, or1192;
  wire b_inv1192;
  assign b_inv1192 = ~b1192;
  assign s1192  = a1192 ^ b1192 ^ c1192;
  assign sub1192 = a1192 ^ b_inv1192 ^ c1192;
  assign and1192 = a1192 & b1192;
  assign or1192  = a1192 | b1192;
  assign c1193 = (a1192 & b1192) | (a1192 & c1192) | (b1192 & c1192);
  wire c_sub1193;
  assign c_sub1193 = (a1192 & b_inv1192) | (a1192 & c1192) | (b_inv1192 & c1192);
  wire s1193, sub1193, and1193, or1193;
  wire b_inv1193;
  assign b_inv1193 = ~b1193;
  assign s1193  = a1193 ^ b1193 ^ c1193;
  assign sub1193 = a1193 ^ b_inv1193 ^ c1193;
  assign and1193 = a1193 & b1193;
  assign or1193  = a1193 | b1193;
  assign c1194 = (a1193 & b1193) | (a1193 & c1193) | (b1193 & c1193);
  wire c_sub1194;
  assign c_sub1194 = (a1193 & b_inv1193) | (a1193 & c1193) | (b_inv1193 & c1193);
  wire s1194, sub1194, and1194, or1194;
  wire b_inv1194;
  assign b_inv1194 = ~b1194;
  assign s1194  = a1194 ^ b1194 ^ c1194;
  assign sub1194 = a1194 ^ b_inv1194 ^ c1194;
  assign and1194 = a1194 & b1194;
  assign or1194  = a1194 | b1194;
  assign c1195 = (a1194 & b1194) | (a1194 & c1194) | (b1194 & c1194);
  wire c_sub1195;
  assign c_sub1195 = (a1194 & b_inv1194) | (a1194 & c1194) | (b_inv1194 & c1194);
  wire s1195, sub1195, and1195, or1195;
  wire b_inv1195;
  assign b_inv1195 = ~b1195;
  assign s1195  = a1195 ^ b1195 ^ c1195;
  assign sub1195 = a1195 ^ b_inv1195 ^ c1195;
  assign and1195 = a1195 & b1195;
  assign or1195  = a1195 | b1195;
  assign c1196 = (a1195 & b1195) | (a1195 & c1195) | (b1195 & c1195);
  wire c_sub1196;
  assign c_sub1196 = (a1195 & b_inv1195) | (a1195 & c1195) | (b_inv1195 & c1195);
  wire s1196, sub1196, and1196, or1196;
  wire b_inv1196;
  assign b_inv1196 = ~b1196;
  assign s1196  = a1196 ^ b1196 ^ c1196;
  assign sub1196 = a1196 ^ b_inv1196 ^ c1196;
  assign and1196 = a1196 & b1196;
  assign or1196  = a1196 | b1196;
  assign c1197 = (a1196 & b1196) | (a1196 & c1196) | (b1196 & c1196);
  wire c_sub1197;
  assign c_sub1197 = (a1196 & b_inv1196) | (a1196 & c1196) | (b_inv1196 & c1196);
  wire s1197, sub1197, and1197, or1197;
  wire b_inv1197;
  assign b_inv1197 = ~b1197;
  assign s1197  = a1197 ^ b1197 ^ c1197;
  assign sub1197 = a1197 ^ b_inv1197 ^ c1197;
  assign and1197 = a1197 & b1197;
  assign or1197  = a1197 | b1197;
  assign c1198 = (a1197 & b1197) | (a1197 & c1197) | (b1197 & c1197);
  wire c_sub1198;
  assign c_sub1198 = (a1197 & b_inv1197) | (a1197 & c1197) | (b_inv1197 & c1197);
  wire s1198, sub1198, and1198, or1198;
  wire b_inv1198;
  assign b_inv1198 = ~b1198;
  assign s1198  = a1198 ^ b1198 ^ c1198;
  assign sub1198 = a1198 ^ b_inv1198 ^ c1198;
  assign and1198 = a1198 & b1198;
  assign or1198  = a1198 | b1198;
  assign c1199 = (a1198 & b1198) | (a1198 & c1198) | (b1198 & c1198);
  wire c_sub1199;
  assign c_sub1199 = (a1198 & b_inv1198) | (a1198 & c1198) | (b_inv1198 & c1198);
  wire s1199, sub1199, and1199, or1199;
  wire b_inv1199;
  assign b_inv1199 = ~b1199;
  assign s1199  = a1199 ^ b1199 ^ c1199;
  assign sub1199 = a1199 ^ b_inv1199 ^ c1199;
  assign and1199 = a1199 & b1199;
  assign or1199  = a1199 | b1199;
  assign c1200 = (a1199 & b1199) | (a1199 & c1199) | (b1199 & c1199);
  wire c_sub1200;
  assign c_sub1200 = (a1199 & b_inv1199) | (a1199 & c1199) | (b_inv1199 & c1199);
  wire s1200, sub1200, and1200, or1200;
  wire b_inv1200;
  assign b_inv1200 = ~b1200;
  assign s1200  = a1200 ^ b1200 ^ c1200;
  assign sub1200 = a1200 ^ b_inv1200 ^ c1200;
  assign and1200 = a1200 & b1200;
  assign or1200  = a1200 | b1200;
  assign c1201 = (a1200 & b1200) | (a1200 & c1200) | (b1200 & c1200);
  wire c_sub1201;
  assign c_sub1201 = (a1200 & b_inv1200) | (a1200 & c1200) | (b_inv1200 & c1200);
  wire s1201, sub1201, and1201, or1201;
  wire b_inv1201;
  assign b_inv1201 = ~b1201;
  assign s1201  = a1201 ^ b1201 ^ c1201;
  assign sub1201 = a1201 ^ b_inv1201 ^ c1201;
  assign and1201 = a1201 & b1201;
  assign or1201  = a1201 | b1201;
  assign c1202 = (a1201 & b1201) | (a1201 & c1201) | (b1201 & c1201);
  wire c_sub1202;
  assign c_sub1202 = (a1201 & b_inv1201) | (a1201 & c1201) | (b_inv1201 & c1201);
  wire s1202, sub1202, and1202, or1202;
  wire b_inv1202;
  assign b_inv1202 = ~b1202;
  assign s1202  = a1202 ^ b1202 ^ c1202;
  assign sub1202 = a1202 ^ b_inv1202 ^ c1202;
  assign and1202 = a1202 & b1202;
  assign or1202  = a1202 | b1202;
  assign c1203 = (a1202 & b1202) | (a1202 & c1202) | (b1202 & c1202);
  wire c_sub1203;
  assign c_sub1203 = (a1202 & b_inv1202) | (a1202 & c1202) | (b_inv1202 & c1202);
  wire s1203, sub1203, and1203, or1203;
  wire b_inv1203;
  assign b_inv1203 = ~b1203;
  assign s1203  = a1203 ^ b1203 ^ c1203;
  assign sub1203 = a1203 ^ b_inv1203 ^ c1203;
  assign and1203 = a1203 & b1203;
  assign or1203  = a1203 | b1203;
  assign c1204 = (a1203 & b1203) | (a1203 & c1203) | (b1203 & c1203);
  wire c_sub1204;
  assign c_sub1204 = (a1203 & b_inv1203) | (a1203 & c1203) | (b_inv1203 & c1203);
  wire s1204, sub1204, and1204, or1204;
  wire b_inv1204;
  assign b_inv1204 = ~b1204;
  assign s1204  = a1204 ^ b1204 ^ c1204;
  assign sub1204 = a1204 ^ b_inv1204 ^ c1204;
  assign and1204 = a1204 & b1204;
  assign or1204  = a1204 | b1204;
  assign c1205 = (a1204 & b1204) | (a1204 & c1204) | (b1204 & c1204);
  wire c_sub1205;
  assign c_sub1205 = (a1204 & b_inv1204) | (a1204 & c1204) | (b_inv1204 & c1204);
  wire s1205, sub1205, and1205, or1205;
  wire b_inv1205;
  assign b_inv1205 = ~b1205;
  assign s1205  = a1205 ^ b1205 ^ c1205;
  assign sub1205 = a1205 ^ b_inv1205 ^ c1205;
  assign and1205 = a1205 & b1205;
  assign or1205  = a1205 | b1205;
  assign c1206 = (a1205 & b1205) | (a1205 & c1205) | (b1205 & c1205);
  wire c_sub1206;
  assign c_sub1206 = (a1205 & b_inv1205) | (a1205 & c1205) | (b_inv1205 & c1205);
  wire s1206, sub1206, and1206, or1206;
  wire b_inv1206;
  assign b_inv1206 = ~b1206;
  assign s1206  = a1206 ^ b1206 ^ c1206;
  assign sub1206 = a1206 ^ b_inv1206 ^ c1206;
  assign and1206 = a1206 & b1206;
  assign or1206  = a1206 | b1206;
  assign c1207 = (a1206 & b1206) | (a1206 & c1206) | (b1206 & c1206);
  wire c_sub1207;
  assign c_sub1207 = (a1206 & b_inv1206) | (a1206 & c1206) | (b_inv1206 & c1206);
  wire s1207, sub1207, and1207, or1207;
  wire b_inv1207;
  assign b_inv1207 = ~b1207;
  assign s1207  = a1207 ^ b1207 ^ c1207;
  assign sub1207 = a1207 ^ b_inv1207 ^ c1207;
  assign and1207 = a1207 & b1207;
  assign or1207  = a1207 | b1207;
  assign c1208 = (a1207 & b1207) | (a1207 & c1207) | (b1207 & c1207);
  wire c_sub1208;
  assign c_sub1208 = (a1207 & b_inv1207) | (a1207 & c1207) | (b_inv1207 & c1207);
  wire s1208, sub1208, and1208, or1208;
  wire b_inv1208;
  assign b_inv1208 = ~b1208;
  assign s1208  = a1208 ^ b1208 ^ c1208;
  assign sub1208 = a1208 ^ b_inv1208 ^ c1208;
  assign and1208 = a1208 & b1208;
  assign or1208  = a1208 | b1208;
  assign c1209 = (a1208 & b1208) | (a1208 & c1208) | (b1208 & c1208);
  wire c_sub1209;
  assign c_sub1209 = (a1208 & b_inv1208) | (a1208 & c1208) | (b_inv1208 & c1208);
  wire s1209, sub1209, and1209, or1209;
  wire b_inv1209;
  assign b_inv1209 = ~b1209;
  assign s1209  = a1209 ^ b1209 ^ c1209;
  assign sub1209 = a1209 ^ b_inv1209 ^ c1209;
  assign and1209 = a1209 & b1209;
  assign or1209  = a1209 | b1209;
  assign c1210 = (a1209 & b1209) | (a1209 & c1209) | (b1209 & c1209);
  wire c_sub1210;
  assign c_sub1210 = (a1209 & b_inv1209) | (a1209 & c1209) | (b_inv1209 & c1209);
  wire s1210, sub1210, and1210, or1210;
  wire b_inv1210;
  assign b_inv1210 = ~b1210;
  assign s1210  = a1210 ^ b1210 ^ c1210;
  assign sub1210 = a1210 ^ b_inv1210 ^ c1210;
  assign and1210 = a1210 & b1210;
  assign or1210  = a1210 | b1210;
  assign c1211 = (a1210 & b1210) | (a1210 & c1210) | (b1210 & c1210);
  wire c_sub1211;
  assign c_sub1211 = (a1210 & b_inv1210) | (a1210 & c1210) | (b_inv1210 & c1210);
  wire s1211, sub1211, and1211, or1211;
  wire b_inv1211;
  assign b_inv1211 = ~b1211;
  assign s1211  = a1211 ^ b1211 ^ c1211;
  assign sub1211 = a1211 ^ b_inv1211 ^ c1211;
  assign and1211 = a1211 & b1211;
  assign or1211  = a1211 | b1211;
  assign c1212 = (a1211 & b1211) | (a1211 & c1211) | (b1211 & c1211);
  wire c_sub1212;
  assign c_sub1212 = (a1211 & b_inv1211) | (a1211 & c1211) | (b_inv1211 & c1211);
  wire s1212, sub1212, and1212, or1212;
  wire b_inv1212;
  assign b_inv1212 = ~b1212;
  assign s1212  = a1212 ^ b1212 ^ c1212;
  assign sub1212 = a1212 ^ b_inv1212 ^ c1212;
  assign and1212 = a1212 & b1212;
  assign or1212  = a1212 | b1212;
  assign c1213 = (a1212 & b1212) | (a1212 & c1212) | (b1212 & c1212);
  wire c_sub1213;
  assign c_sub1213 = (a1212 & b_inv1212) | (a1212 & c1212) | (b_inv1212 & c1212);
  wire s1213, sub1213, and1213, or1213;
  wire b_inv1213;
  assign b_inv1213 = ~b1213;
  assign s1213  = a1213 ^ b1213 ^ c1213;
  assign sub1213 = a1213 ^ b_inv1213 ^ c1213;
  assign and1213 = a1213 & b1213;
  assign or1213  = a1213 | b1213;
  assign c1214 = (a1213 & b1213) | (a1213 & c1213) | (b1213 & c1213);
  wire c_sub1214;
  assign c_sub1214 = (a1213 & b_inv1213) | (a1213 & c1213) | (b_inv1213 & c1213);
  wire s1214, sub1214, and1214, or1214;
  wire b_inv1214;
  assign b_inv1214 = ~b1214;
  assign s1214  = a1214 ^ b1214 ^ c1214;
  assign sub1214 = a1214 ^ b_inv1214 ^ c1214;
  assign and1214 = a1214 & b1214;
  assign or1214  = a1214 | b1214;
  assign c1215 = (a1214 & b1214) | (a1214 & c1214) | (b1214 & c1214);
  wire c_sub1215;
  assign c_sub1215 = (a1214 & b_inv1214) | (a1214 & c1214) | (b_inv1214 & c1214);
  wire s1215, sub1215, and1215, or1215;
  wire b_inv1215;
  assign b_inv1215 = ~b1215;
  assign s1215  = a1215 ^ b1215 ^ c1215;
  assign sub1215 = a1215 ^ b_inv1215 ^ c1215;
  assign and1215 = a1215 & b1215;
  assign or1215  = a1215 | b1215;
  assign c1216 = (a1215 & b1215) | (a1215 & c1215) | (b1215 & c1215);
  wire c_sub1216;
  assign c_sub1216 = (a1215 & b_inv1215) | (a1215 & c1215) | (b_inv1215 & c1215);
  wire s1216, sub1216, and1216, or1216;
  wire b_inv1216;
  assign b_inv1216 = ~b1216;
  assign s1216  = a1216 ^ b1216 ^ c1216;
  assign sub1216 = a1216 ^ b_inv1216 ^ c1216;
  assign and1216 = a1216 & b1216;
  assign or1216  = a1216 | b1216;
  assign c1217 = (a1216 & b1216) | (a1216 & c1216) | (b1216 & c1216);
  wire c_sub1217;
  assign c_sub1217 = (a1216 & b_inv1216) | (a1216 & c1216) | (b_inv1216 & c1216);
  wire s1217, sub1217, and1217, or1217;
  wire b_inv1217;
  assign b_inv1217 = ~b1217;
  assign s1217  = a1217 ^ b1217 ^ c1217;
  assign sub1217 = a1217 ^ b_inv1217 ^ c1217;
  assign and1217 = a1217 & b1217;
  assign or1217  = a1217 | b1217;
  assign c1218 = (a1217 & b1217) | (a1217 & c1217) | (b1217 & c1217);
  wire c_sub1218;
  assign c_sub1218 = (a1217 & b_inv1217) | (a1217 & c1217) | (b_inv1217 & c1217);
  wire s1218, sub1218, and1218, or1218;
  wire b_inv1218;
  assign b_inv1218 = ~b1218;
  assign s1218  = a1218 ^ b1218 ^ c1218;
  assign sub1218 = a1218 ^ b_inv1218 ^ c1218;
  assign and1218 = a1218 & b1218;
  assign or1218  = a1218 | b1218;
  assign c1219 = (a1218 & b1218) | (a1218 & c1218) | (b1218 & c1218);
  wire c_sub1219;
  assign c_sub1219 = (a1218 & b_inv1218) | (a1218 & c1218) | (b_inv1218 & c1218);
  wire s1219, sub1219, and1219, or1219;
  wire b_inv1219;
  assign b_inv1219 = ~b1219;
  assign s1219  = a1219 ^ b1219 ^ c1219;
  assign sub1219 = a1219 ^ b_inv1219 ^ c1219;
  assign and1219 = a1219 & b1219;
  assign or1219  = a1219 | b1219;
  assign c1220 = (a1219 & b1219) | (a1219 & c1219) | (b1219 & c1219);
  wire c_sub1220;
  assign c_sub1220 = (a1219 & b_inv1219) | (a1219 & c1219) | (b_inv1219 & c1219);
  wire s1220, sub1220, and1220, or1220;
  wire b_inv1220;
  assign b_inv1220 = ~b1220;
  assign s1220  = a1220 ^ b1220 ^ c1220;
  assign sub1220 = a1220 ^ b_inv1220 ^ c1220;
  assign and1220 = a1220 & b1220;
  assign or1220  = a1220 | b1220;
  assign c1221 = (a1220 & b1220) | (a1220 & c1220) | (b1220 & c1220);
  wire c_sub1221;
  assign c_sub1221 = (a1220 & b_inv1220) | (a1220 & c1220) | (b_inv1220 & c1220);
  wire s1221, sub1221, and1221, or1221;
  wire b_inv1221;
  assign b_inv1221 = ~b1221;
  assign s1221  = a1221 ^ b1221 ^ c1221;
  assign sub1221 = a1221 ^ b_inv1221 ^ c1221;
  assign and1221 = a1221 & b1221;
  assign or1221  = a1221 | b1221;
  assign c1222 = (a1221 & b1221) | (a1221 & c1221) | (b1221 & c1221);
  wire c_sub1222;
  assign c_sub1222 = (a1221 & b_inv1221) | (a1221 & c1221) | (b_inv1221 & c1221);
  wire s1222, sub1222, and1222, or1222;
  wire b_inv1222;
  assign b_inv1222 = ~b1222;
  assign s1222  = a1222 ^ b1222 ^ c1222;
  assign sub1222 = a1222 ^ b_inv1222 ^ c1222;
  assign and1222 = a1222 & b1222;
  assign or1222  = a1222 | b1222;
  assign c1223 = (a1222 & b1222) | (a1222 & c1222) | (b1222 & c1222);
  wire c_sub1223;
  assign c_sub1223 = (a1222 & b_inv1222) | (a1222 & c1222) | (b_inv1222 & c1222);
  wire s1223, sub1223, and1223, or1223;
  wire b_inv1223;
  assign b_inv1223 = ~b1223;
  assign s1223  = a1223 ^ b1223 ^ c1223;
  assign sub1223 = a1223 ^ b_inv1223 ^ c1223;
  assign and1223 = a1223 & b1223;
  assign or1223  = a1223 | b1223;
  assign c1224 = (a1223 & b1223) | (a1223 & c1223) | (b1223 & c1223);
  wire c_sub1224;
  assign c_sub1224 = (a1223 & b_inv1223) | (a1223 & c1223) | (b_inv1223 & c1223);
  wire s1224, sub1224, and1224, or1224;
  wire b_inv1224;
  assign b_inv1224 = ~b1224;
  assign s1224  = a1224 ^ b1224 ^ c1224;
  assign sub1224 = a1224 ^ b_inv1224 ^ c1224;
  assign and1224 = a1224 & b1224;
  assign or1224  = a1224 | b1224;
  assign c1225 = (a1224 & b1224) | (a1224 & c1224) | (b1224 & c1224);
  wire c_sub1225;
  assign c_sub1225 = (a1224 & b_inv1224) | (a1224 & c1224) | (b_inv1224 & c1224);
  wire s1225, sub1225, and1225, or1225;
  wire b_inv1225;
  assign b_inv1225 = ~b1225;
  assign s1225  = a1225 ^ b1225 ^ c1225;
  assign sub1225 = a1225 ^ b_inv1225 ^ c1225;
  assign and1225 = a1225 & b1225;
  assign or1225  = a1225 | b1225;
  assign c1226 = (a1225 & b1225) | (a1225 & c1225) | (b1225 & c1225);
  wire c_sub1226;
  assign c_sub1226 = (a1225 & b_inv1225) | (a1225 & c1225) | (b_inv1225 & c1225);
  wire s1226, sub1226, and1226, or1226;
  wire b_inv1226;
  assign b_inv1226 = ~b1226;
  assign s1226  = a1226 ^ b1226 ^ c1226;
  assign sub1226 = a1226 ^ b_inv1226 ^ c1226;
  assign and1226 = a1226 & b1226;
  assign or1226  = a1226 | b1226;
  assign c1227 = (a1226 & b1226) | (a1226 & c1226) | (b1226 & c1226);
  wire c_sub1227;
  assign c_sub1227 = (a1226 & b_inv1226) | (a1226 & c1226) | (b_inv1226 & c1226);
  wire s1227, sub1227, and1227, or1227;
  wire b_inv1227;
  assign b_inv1227 = ~b1227;
  assign s1227  = a1227 ^ b1227 ^ c1227;
  assign sub1227 = a1227 ^ b_inv1227 ^ c1227;
  assign and1227 = a1227 & b1227;
  assign or1227  = a1227 | b1227;
  assign c1228 = (a1227 & b1227) | (a1227 & c1227) | (b1227 & c1227);
  wire c_sub1228;
  assign c_sub1228 = (a1227 & b_inv1227) | (a1227 & c1227) | (b_inv1227 & c1227);
  wire s1228, sub1228, and1228, or1228;
  wire b_inv1228;
  assign b_inv1228 = ~b1228;
  assign s1228  = a1228 ^ b1228 ^ c1228;
  assign sub1228 = a1228 ^ b_inv1228 ^ c1228;
  assign and1228 = a1228 & b1228;
  assign or1228  = a1228 | b1228;
  assign c1229 = (a1228 & b1228) | (a1228 & c1228) | (b1228 & c1228);
  wire c_sub1229;
  assign c_sub1229 = (a1228 & b_inv1228) | (a1228 & c1228) | (b_inv1228 & c1228);
  wire s1229, sub1229, and1229, or1229;
  wire b_inv1229;
  assign b_inv1229 = ~b1229;
  assign s1229  = a1229 ^ b1229 ^ c1229;
  assign sub1229 = a1229 ^ b_inv1229 ^ c1229;
  assign and1229 = a1229 & b1229;
  assign or1229  = a1229 | b1229;
  assign c1230 = (a1229 & b1229) | (a1229 & c1229) | (b1229 & c1229);
  wire c_sub1230;
  assign c_sub1230 = (a1229 & b_inv1229) | (a1229 & c1229) | (b_inv1229 & c1229);
  wire s1230, sub1230, and1230, or1230;
  wire b_inv1230;
  assign b_inv1230 = ~b1230;
  assign s1230  = a1230 ^ b1230 ^ c1230;
  assign sub1230 = a1230 ^ b_inv1230 ^ c1230;
  assign and1230 = a1230 & b1230;
  assign or1230  = a1230 | b1230;
  assign c1231 = (a1230 & b1230) | (a1230 & c1230) | (b1230 & c1230);
  wire c_sub1231;
  assign c_sub1231 = (a1230 & b_inv1230) | (a1230 & c1230) | (b_inv1230 & c1230);
  wire s1231, sub1231, and1231, or1231;
  wire b_inv1231;
  assign b_inv1231 = ~b1231;
  assign s1231  = a1231 ^ b1231 ^ c1231;
  assign sub1231 = a1231 ^ b_inv1231 ^ c1231;
  assign and1231 = a1231 & b1231;
  assign or1231  = a1231 | b1231;
  assign c1232 = (a1231 & b1231) | (a1231 & c1231) | (b1231 & c1231);
  wire c_sub1232;
  assign c_sub1232 = (a1231 & b_inv1231) | (a1231 & c1231) | (b_inv1231 & c1231);
  wire s1232, sub1232, and1232, or1232;
  wire b_inv1232;
  assign b_inv1232 = ~b1232;
  assign s1232  = a1232 ^ b1232 ^ c1232;
  assign sub1232 = a1232 ^ b_inv1232 ^ c1232;
  assign and1232 = a1232 & b1232;
  assign or1232  = a1232 | b1232;
  assign c1233 = (a1232 & b1232) | (a1232 & c1232) | (b1232 & c1232);
  wire c_sub1233;
  assign c_sub1233 = (a1232 & b_inv1232) | (a1232 & c1232) | (b_inv1232 & c1232);
  wire s1233, sub1233, and1233, or1233;
  wire b_inv1233;
  assign b_inv1233 = ~b1233;
  assign s1233  = a1233 ^ b1233 ^ c1233;
  assign sub1233 = a1233 ^ b_inv1233 ^ c1233;
  assign and1233 = a1233 & b1233;
  assign or1233  = a1233 | b1233;
  assign c1234 = (a1233 & b1233) | (a1233 & c1233) | (b1233 & c1233);
  wire c_sub1234;
  assign c_sub1234 = (a1233 & b_inv1233) | (a1233 & c1233) | (b_inv1233 & c1233);
  wire s1234, sub1234, and1234, or1234;
  wire b_inv1234;
  assign b_inv1234 = ~b1234;
  assign s1234  = a1234 ^ b1234 ^ c1234;
  assign sub1234 = a1234 ^ b_inv1234 ^ c1234;
  assign and1234 = a1234 & b1234;
  assign or1234  = a1234 | b1234;
  assign c1235 = (a1234 & b1234) | (a1234 & c1234) | (b1234 & c1234);
  wire c_sub1235;
  assign c_sub1235 = (a1234 & b_inv1234) | (a1234 & c1234) | (b_inv1234 & c1234);
  wire s1235, sub1235, and1235, or1235;
  wire b_inv1235;
  assign b_inv1235 = ~b1235;
  assign s1235  = a1235 ^ b1235 ^ c1235;
  assign sub1235 = a1235 ^ b_inv1235 ^ c1235;
  assign and1235 = a1235 & b1235;
  assign or1235  = a1235 | b1235;
  assign c1236 = (a1235 & b1235) | (a1235 & c1235) | (b1235 & c1235);
  wire c_sub1236;
  assign c_sub1236 = (a1235 & b_inv1235) | (a1235 & c1235) | (b_inv1235 & c1235);
  wire s1236, sub1236, and1236, or1236;
  wire b_inv1236;
  assign b_inv1236 = ~b1236;
  assign s1236  = a1236 ^ b1236 ^ c1236;
  assign sub1236 = a1236 ^ b_inv1236 ^ c1236;
  assign and1236 = a1236 & b1236;
  assign or1236  = a1236 | b1236;
  assign c1237 = (a1236 & b1236) | (a1236 & c1236) | (b1236 & c1236);
  wire c_sub1237;
  assign c_sub1237 = (a1236 & b_inv1236) | (a1236 & c1236) | (b_inv1236 & c1236);
  wire s1237, sub1237, and1237, or1237;
  wire b_inv1237;
  assign b_inv1237 = ~b1237;
  assign s1237  = a1237 ^ b1237 ^ c1237;
  assign sub1237 = a1237 ^ b_inv1237 ^ c1237;
  assign and1237 = a1237 & b1237;
  assign or1237  = a1237 | b1237;
  assign c1238 = (a1237 & b1237) | (a1237 & c1237) | (b1237 & c1237);
  wire c_sub1238;
  assign c_sub1238 = (a1237 & b_inv1237) | (a1237 & c1237) | (b_inv1237 & c1237);
  wire s1238, sub1238, and1238, or1238;
  wire b_inv1238;
  assign b_inv1238 = ~b1238;
  assign s1238  = a1238 ^ b1238 ^ c1238;
  assign sub1238 = a1238 ^ b_inv1238 ^ c1238;
  assign and1238 = a1238 & b1238;
  assign or1238  = a1238 | b1238;
  assign c1239 = (a1238 & b1238) | (a1238 & c1238) | (b1238 & c1238);
  wire c_sub1239;
  assign c_sub1239 = (a1238 & b_inv1238) | (a1238 & c1238) | (b_inv1238 & c1238);
  wire s1239, sub1239, and1239, or1239;
  wire b_inv1239;
  assign b_inv1239 = ~b1239;
  assign s1239  = a1239 ^ b1239 ^ c1239;
  assign sub1239 = a1239 ^ b_inv1239 ^ c1239;
  assign and1239 = a1239 & b1239;
  assign or1239  = a1239 | b1239;
  assign c1240 = (a1239 & b1239) | (a1239 & c1239) | (b1239 & c1239);
  wire c_sub1240;
  assign c_sub1240 = (a1239 & b_inv1239) | (a1239 & c1239) | (b_inv1239 & c1239);
  wire s1240, sub1240, and1240, or1240;
  wire b_inv1240;
  assign b_inv1240 = ~b1240;
  assign s1240  = a1240 ^ b1240 ^ c1240;
  assign sub1240 = a1240 ^ b_inv1240 ^ c1240;
  assign and1240 = a1240 & b1240;
  assign or1240  = a1240 | b1240;
  assign c1241 = (a1240 & b1240) | (a1240 & c1240) | (b1240 & c1240);
  wire c_sub1241;
  assign c_sub1241 = (a1240 & b_inv1240) | (a1240 & c1240) | (b_inv1240 & c1240);
  wire s1241, sub1241, and1241, or1241;
  wire b_inv1241;
  assign b_inv1241 = ~b1241;
  assign s1241  = a1241 ^ b1241 ^ c1241;
  assign sub1241 = a1241 ^ b_inv1241 ^ c1241;
  assign and1241 = a1241 & b1241;
  assign or1241  = a1241 | b1241;
  assign c1242 = (a1241 & b1241) | (a1241 & c1241) | (b1241 & c1241);
  wire c_sub1242;
  assign c_sub1242 = (a1241 & b_inv1241) | (a1241 & c1241) | (b_inv1241 & c1241);
  wire s1242, sub1242, and1242, or1242;
  wire b_inv1242;
  assign b_inv1242 = ~b1242;
  assign s1242  = a1242 ^ b1242 ^ c1242;
  assign sub1242 = a1242 ^ b_inv1242 ^ c1242;
  assign and1242 = a1242 & b1242;
  assign or1242  = a1242 | b1242;
  assign c1243 = (a1242 & b1242) | (a1242 & c1242) | (b1242 & c1242);
  wire c_sub1243;
  assign c_sub1243 = (a1242 & b_inv1242) | (a1242 & c1242) | (b_inv1242 & c1242);
  wire s1243, sub1243, and1243, or1243;
  wire b_inv1243;
  assign b_inv1243 = ~b1243;
  assign s1243  = a1243 ^ b1243 ^ c1243;
  assign sub1243 = a1243 ^ b_inv1243 ^ c1243;
  assign and1243 = a1243 & b1243;
  assign or1243  = a1243 | b1243;
  assign c1244 = (a1243 & b1243) | (a1243 & c1243) | (b1243 & c1243);
  wire c_sub1244;
  assign c_sub1244 = (a1243 & b_inv1243) | (a1243 & c1243) | (b_inv1243 & c1243);
  wire s1244, sub1244, and1244, or1244;
  wire b_inv1244;
  assign b_inv1244 = ~b1244;
  assign s1244  = a1244 ^ b1244 ^ c1244;
  assign sub1244 = a1244 ^ b_inv1244 ^ c1244;
  assign and1244 = a1244 & b1244;
  assign or1244  = a1244 | b1244;
  assign c1245 = (a1244 & b1244) | (a1244 & c1244) | (b1244 & c1244);
  wire c_sub1245;
  assign c_sub1245 = (a1244 & b_inv1244) | (a1244 & c1244) | (b_inv1244 & c1244);
  wire s1245, sub1245, and1245, or1245;
  wire b_inv1245;
  assign b_inv1245 = ~b1245;
  assign s1245  = a1245 ^ b1245 ^ c1245;
  assign sub1245 = a1245 ^ b_inv1245 ^ c1245;
  assign and1245 = a1245 & b1245;
  assign or1245  = a1245 | b1245;
  assign c1246 = (a1245 & b1245) | (a1245 & c1245) | (b1245 & c1245);
  wire c_sub1246;
  assign c_sub1246 = (a1245 & b_inv1245) | (a1245 & c1245) | (b_inv1245 & c1245);
  wire s1246, sub1246, and1246, or1246;
  wire b_inv1246;
  assign b_inv1246 = ~b1246;
  assign s1246  = a1246 ^ b1246 ^ c1246;
  assign sub1246 = a1246 ^ b_inv1246 ^ c1246;
  assign and1246 = a1246 & b1246;
  assign or1246  = a1246 | b1246;
  assign c1247 = (a1246 & b1246) | (a1246 & c1246) | (b1246 & c1246);
  wire c_sub1247;
  assign c_sub1247 = (a1246 & b_inv1246) | (a1246 & c1246) | (b_inv1246 & c1246);
  wire s1247, sub1247, and1247, or1247;
  wire b_inv1247;
  assign b_inv1247 = ~b1247;
  assign s1247  = a1247 ^ b1247 ^ c1247;
  assign sub1247 = a1247 ^ b_inv1247 ^ c1247;
  assign and1247 = a1247 & b1247;
  assign or1247  = a1247 | b1247;
  assign c1248 = (a1247 & b1247) | (a1247 & c1247) | (b1247 & c1247);
  wire c_sub1248;
  assign c_sub1248 = (a1247 & b_inv1247) | (a1247 & c1247) | (b_inv1247 & c1247);
  wire s1248, sub1248, and1248, or1248;
  wire b_inv1248;
  assign b_inv1248 = ~b1248;
  assign s1248  = a1248 ^ b1248 ^ c1248;
  assign sub1248 = a1248 ^ b_inv1248 ^ c1248;
  assign and1248 = a1248 & b1248;
  assign or1248  = a1248 | b1248;
  assign c1249 = (a1248 & b1248) | (a1248 & c1248) | (b1248 & c1248);
  wire c_sub1249;
  assign c_sub1249 = (a1248 & b_inv1248) | (a1248 & c1248) | (b_inv1248 & c1248);
  wire s1249, sub1249, and1249, or1249;
  wire b_inv1249;
  assign b_inv1249 = ~b1249;
  assign s1249  = a1249 ^ b1249 ^ c1249;
  assign sub1249 = a1249 ^ b_inv1249 ^ c1249;
  assign and1249 = a1249 & b1249;
  assign or1249  = a1249 | b1249;
  assign c1250 = (a1249 & b1249) | (a1249 & c1249) | (b1249 & c1249);
  wire c_sub1250;
  assign c_sub1250 = (a1249 & b_inv1249) | (a1249 & c1249) | (b_inv1249 & c1249);
  wire s1250, sub1250, and1250, or1250;
  wire b_inv1250;
  assign b_inv1250 = ~b1250;
  assign s1250  = a1250 ^ b1250 ^ c1250;
  assign sub1250 = a1250 ^ b_inv1250 ^ c1250;
  assign and1250 = a1250 & b1250;
  assign or1250  = a1250 | b1250;
  assign c1251 = (a1250 & b1250) | (a1250 & c1250) | (b1250 & c1250);
  wire c_sub1251;
  assign c_sub1251 = (a1250 & b_inv1250) | (a1250 & c1250) | (b_inv1250 & c1250);
  wire s1251, sub1251, and1251, or1251;
  wire b_inv1251;
  assign b_inv1251 = ~b1251;
  assign s1251  = a1251 ^ b1251 ^ c1251;
  assign sub1251 = a1251 ^ b_inv1251 ^ c1251;
  assign and1251 = a1251 & b1251;
  assign or1251  = a1251 | b1251;
  assign c1252 = (a1251 & b1251) | (a1251 & c1251) | (b1251 & c1251);
  wire c_sub1252;
  assign c_sub1252 = (a1251 & b_inv1251) | (a1251 & c1251) | (b_inv1251 & c1251);
  wire s1252, sub1252, and1252, or1252;
  wire b_inv1252;
  assign b_inv1252 = ~b1252;
  assign s1252  = a1252 ^ b1252 ^ c1252;
  assign sub1252 = a1252 ^ b_inv1252 ^ c1252;
  assign and1252 = a1252 & b1252;
  assign or1252  = a1252 | b1252;
  assign c1253 = (a1252 & b1252) | (a1252 & c1252) | (b1252 & c1252);
  wire c_sub1253;
  assign c_sub1253 = (a1252 & b_inv1252) | (a1252 & c1252) | (b_inv1252 & c1252);
  wire s1253, sub1253, and1253, or1253;
  wire b_inv1253;
  assign b_inv1253 = ~b1253;
  assign s1253  = a1253 ^ b1253 ^ c1253;
  assign sub1253 = a1253 ^ b_inv1253 ^ c1253;
  assign and1253 = a1253 & b1253;
  assign or1253  = a1253 | b1253;
  assign c1254 = (a1253 & b1253) | (a1253 & c1253) | (b1253 & c1253);
  wire c_sub1254;
  assign c_sub1254 = (a1253 & b_inv1253) | (a1253 & c1253) | (b_inv1253 & c1253);
  wire s1254, sub1254, and1254, or1254;
  wire b_inv1254;
  assign b_inv1254 = ~b1254;
  assign s1254  = a1254 ^ b1254 ^ c1254;
  assign sub1254 = a1254 ^ b_inv1254 ^ c1254;
  assign and1254 = a1254 & b1254;
  assign or1254  = a1254 | b1254;
  assign c1255 = (a1254 & b1254) | (a1254 & c1254) | (b1254 & c1254);
  wire c_sub1255;
  assign c_sub1255 = (a1254 & b_inv1254) | (a1254 & c1254) | (b_inv1254 & c1254);
  wire s1255, sub1255, and1255, or1255;
  wire b_inv1255;
  assign b_inv1255 = ~b1255;
  assign s1255  = a1255 ^ b1255 ^ c1255;
  assign sub1255 = a1255 ^ b_inv1255 ^ c1255;
  assign and1255 = a1255 & b1255;
  assign or1255  = a1255 | b1255;
  assign c1256 = (a1255 & b1255) | (a1255 & c1255) | (b1255 & c1255);
  wire c_sub1256;
  assign c_sub1256 = (a1255 & b_inv1255) | (a1255 & c1255) | (b_inv1255 & c1255);
  wire s1256, sub1256, and1256, or1256;
  wire b_inv1256;
  assign b_inv1256 = ~b1256;
  assign s1256  = a1256 ^ b1256 ^ c1256;
  assign sub1256 = a1256 ^ b_inv1256 ^ c1256;
  assign and1256 = a1256 & b1256;
  assign or1256  = a1256 | b1256;
  assign c1257 = (a1256 & b1256) | (a1256 & c1256) | (b1256 & c1256);
  wire c_sub1257;
  assign c_sub1257 = (a1256 & b_inv1256) | (a1256 & c1256) | (b_inv1256 & c1256);
  wire s1257, sub1257, and1257, or1257;
  wire b_inv1257;
  assign b_inv1257 = ~b1257;
  assign s1257  = a1257 ^ b1257 ^ c1257;
  assign sub1257 = a1257 ^ b_inv1257 ^ c1257;
  assign and1257 = a1257 & b1257;
  assign or1257  = a1257 | b1257;
  assign c1258 = (a1257 & b1257) | (a1257 & c1257) | (b1257 & c1257);
  wire c_sub1258;
  assign c_sub1258 = (a1257 & b_inv1257) | (a1257 & c1257) | (b_inv1257 & c1257);
  wire s1258, sub1258, and1258, or1258;
  wire b_inv1258;
  assign b_inv1258 = ~b1258;
  assign s1258  = a1258 ^ b1258 ^ c1258;
  assign sub1258 = a1258 ^ b_inv1258 ^ c1258;
  assign and1258 = a1258 & b1258;
  assign or1258  = a1258 | b1258;
  assign c1259 = (a1258 & b1258) | (a1258 & c1258) | (b1258 & c1258);
  wire c_sub1259;
  assign c_sub1259 = (a1258 & b_inv1258) | (a1258 & c1258) | (b_inv1258 & c1258);
  wire s1259, sub1259, and1259, or1259;
  wire b_inv1259;
  assign b_inv1259 = ~b1259;
  assign s1259  = a1259 ^ b1259 ^ c1259;
  assign sub1259 = a1259 ^ b_inv1259 ^ c1259;
  assign and1259 = a1259 & b1259;
  assign or1259  = a1259 | b1259;
  assign c1260 = (a1259 & b1259) | (a1259 & c1259) | (b1259 & c1259);
  wire c_sub1260;
  assign c_sub1260 = (a1259 & b_inv1259) | (a1259 & c1259) | (b_inv1259 & c1259);
  wire s1260, sub1260, and1260, or1260;
  wire b_inv1260;
  assign b_inv1260 = ~b1260;
  assign s1260  = a1260 ^ b1260 ^ c1260;
  assign sub1260 = a1260 ^ b_inv1260 ^ c1260;
  assign and1260 = a1260 & b1260;
  assign or1260  = a1260 | b1260;
  assign c1261 = (a1260 & b1260) | (a1260 & c1260) | (b1260 & c1260);
  wire c_sub1261;
  assign c_sub1261 = (a1260 & b_inv1260) | (a1260 & c1260) | (b_inv1260 & c1260);
  wire s1261, sub1261, and1261, or1261;
  wire b_inv1261;
  assign b_inv1261 = ~b1261;
  assign s1261  = a1261 ^ b1261 ^ c1261;
  assign sub1261 = a1261 ^ b_inv1261 ^ c1261;
  assign and1261 = a1261 & b1261;
  assign or1261  = a1261 | b1261;
  assign c1262 = (a1261 & b1261) | (a1261 & c1261) | (b1261 & c1261);
  wire c_sub1262;
  assign c_sub1262 = (a1261 & b_inv1261) | (a1261 & c1261) | (b_inv1261 & c1261);
  wire s1262, sub1262, and1262, or1262;
  wire b_inv1262;
  assign b_inv1262 = ~b1262;
  assign s1262  = a1262 ^ b1262 ^ c1262;
  assign sub1262 = a1262 ^ b_inv1262 ^ c1262;
  assign and1262 = a1262 & b1262;
  assign or1262  = a1262 | b1262;
  assign c1263 = (a1262 & b1262) | (a1262 & c1262) | (b1262 & c1262);
  wire c_sub1263;
  assign c_sub1263 = (a1262 & b_inv1262) | (a1262 & c1262) | (b_inv1262 & c1262);
  wire s1263, sub1263, and1263, or1263;
  wire b_inv1263;
  assign b_inv1263 = ~b1263;
  assign s1263  = a1263 ^ b1263 ^ c1263;
  assign sub1263 = a1263 ^ b_inv1263 ^ c1263;
  assign and1263 = a1263 & b1263;
  assign or1263  = a1263 | b1263;
  assign c1264 = (a1263 & b1263) | (a1263 & c1263) | (b1263 & c1263);
  wire c_sub1264;
  assign c_sub1264 = (a1263 & b_inv1263) | (a1263 & c1263) | (b_inv1263 & c1263);
  wire s1264, sub1264, and1264, or1264;
  wire b_inv1264;
  assign b_inv1264 = ~b1264;
  assign s1264  = a1264 ^ b1264 ^ c1264;
  assign sub1264 = a1264 ^ b_inv1264 ^ c1264;
  assign and1264 = a1264 & b1264;
  assign or1264  = a1264 | b1264;
  assign c1265 = (a1264 & b1264) | (a1264 & c1264) | (b1264 & c1264);
  wire c_sub1265;
  assign c_sub1265 = (a1264 & b_inv1264) | (a1264 & c1264) | (b_inv1264 & c1264);
  wire s1265, sub1265, and1265, or1265;
  wire b_inv1265;
  assign b_inv1265 = ~b1265;
  assign s1265  = a1265 ^ b1265 ^ c1265;
  assign sub1265 = a1265 ^ b_inv1265 ^ c1265;
  assign and1265 = a1265 & b1265;
  assign or1265  = a1265 | b1265;
  assign c1266 = (a1265 & b1265) | (a1265 & c1265) | (b1265 & c1265);
  wire c_sub1266;
  assign c_sub1266 = (a1265 & b_inv1265) | (a1265 & c1265) | (b_inv1265 & c1265);
  wire s1266, sub1266, and1266, or1266;
  wire b_inv1266;
  assign b_inv1266 = ~b1266;
  assign s1266  = a1266 ^ b1266 ^ c1266;
  assign sub1266 = a1266 ^ b_inv1266 ^ c1266;
  assign and1266 = a1266 & b1266;
  assign or1266  = a1266 | b1266;
  assign c1267 = (a1266 & b1266) | (a1266 & c1266) | (b1266 & c1266);
  wire c_sub1267;
  assign c_sub1267 = (a1266 & b_inv1266) | (a1266 & c1266) | (b_inv1266 & c1266);
  wire s1267, sub1267, and1267, or1267;
  wire b_inv1267;
  assign b_inv1267 = ~b1267;
  assign s1267  = a1267 ^ b1267 ^ c1267;
  assign sub1267 = a1267 ^ b_inv1267 ^ c1267;
  assign and1267 = a1267 & b1267;
  assign or1267  = a1267 | b1267;
  assign c1268 = (a1267 & b1267) | (a1267 & c1267) | (b1267 & c1267);
  wire c_sub1268;
  assign c_sub1268 = (a1267 & b_inv1267) | (a1267 & c1267) | (b_inv1267 & c1267);
  wire s1268, sub1268, and1268, or1268;
  wire b_inv1268;
  assign b_inv1268 = ~b1268;
  assign s1268  = a1268 ^ b1268 ^ c1268;
  assign sub1268 = a1268 ^ b_inv1268 ^ c1268;
  assign and1268 = a1268 & b1268;
  assign or1268  = a1268 | b1268;
  assign c1269 = (a1268 & b1268) | (a1268 & c1268) | (b1268 & c1268);
  wire c_sub1269;
  assign c_sub1269 = (a1268 & b_inv1268) | (a1268 & c1268) | (b_inv1268 & c1268);
  wire s1269, sub1269, and1269, or1269;
  wire b_inv1269;
  assign b_inv1269 = ~b1269;
  assign s1269  = a1269 ^ b1269 ^ c1269;
  assign sub1269 = a1269 ^ b_inv1269 ^ c1269;
  assign and1269 = a1269 & b1269;
  assign or1269  = a1269 | b1269;
  assign c1270 = (a1269 & b1269) | (a1269 & c1269) | (b1269 & c1269);
  wire c_sub1270;
  assign c_sub1270 = (a1269 & b_inv1269) | (a1269 & c1269) | (b_inv1269 & c1269);
  wire s1270, sub1270, and1270, or1270;
  wire b_inv1270;
  assign b_inv1270 = ~b1270;
  assign s1270  = a1270 ^ b1270 ^ c1270;
  assign sub1270 = a1270 ^ b_inv1270 ^ c1270;
  assign and1270 = a1270 & b1270;
  assign or1270  = a1270 | b1270;
  assign c1271 = (a1270 & b1270) | (a1270 & c1270) | (b1270 & c1270);
  wire c_sub1271;
  assign c_sub1271 = (a1270 & b_inv1270) | (a1270 & c1270) | (b_inv1270 & c1270);
  wire s1271, sub1271, and1271, or1271;
  wire b_inv1271;
  assign b_inv1271 = ~b1271;
  assign s1271  = a1271 ^ b1271 ^ c1271;
  assign sub1271 = a1271 ^ b_inv1271 ^ c1271;
  assign and1271 = a1271 & b1271;
  assign or1271  = a1271 | b1271;
  assign c1272 = (a1271 & b1271) | (a1271 & c1271) | (b1271 & c1271);
  wire c_sub1272;
  assign c_sub1272 = (a1271 & b_inv1271) | (a1271 & c1271) | (b_inv1271 & c1271);
  wire s1272, sub1272, and1272, or1272;
  wire b_inv1272;
  assign b_inv1272 = ~b1272;
  assign s1272  = a1272 ^ b1272 ^ c1272;
  assign sub1272 = a1272 ^ b_inv1272 ^ c1272;
  assign and1272 = a1272 & b1272;
  assign or1272  = a1272 | b1272;
  assign c1273 = (a1272 & b1272) | (a1272 & c1272) | (b1272 & c1272);
  wire c_sub1273;
  assign c_sub1273 = (a1272 & b_inv1272) | (a1272 & c1272) | (b_inv1272 & c1272);
  wire s1273, sub1273, and1273, or1273;
  wire b_inv1273;
  assign b_inv1273 = ~b1273;
  assign s1273  = a1273 ^ b1273 ^ c1273;
  assign sub1273 = a1273 ^ b_inv1273 ^ c1273;
  assign and1273 = a1273 & b1273;
  assign or1273  = a1273 | b1273;
  assign c1274 = (a1273 & b1273) | (a1273 & c1273) | (b1273 & c1273);
  wire c_sub1274;
  assign c_sub1274 = (a1273 & b_inv1273) | (a1273 & c1273) | (b_inv1273 & c1273);
  wire s1274, sub1274, and1274, or1274;
  wire b_inv1274;
  assign b_inv1274 = ~b1274;
  assign s1274  = a1274 ^ b1274 ^ c1274;
  assign sub1274 = a1274 ^ b_inv1274 ^ c1274;
  assign and1274 = a1274 & b1274;
  assign or1274  = a1274 | b1274;
  assign c1275 = (a1274 & b1274) | (a1274 & c1274) | (b1274 & c1274);
  wire c_sub1275;
  assign c_sub1275 = (a1274 & b_inv1274) | (a1274 & c1274) | (b_inv1274 & c1274);
  wire s1275, sub1275, and1275, or1275;
  wire b_inv1275;
  assign b_inv1275 = ~b1275;
  assign s1275  = a1275 ^ b1275 ^ c1275;
  assign sub1275 = a1275 ^ b_inv1275 ^ c1275;
  assign and1275 = a1275 & b1275;
  assign or1275  = a1275 | b1275;
  assign c1276 = (a1275 & b1275) | (a1275 & c1275) | (b1275 & c1275);
  wire c_sub1276;
  assign c_sub1276 = (a1275 & b_inv1275) | (a1275 & c1275) | (b_inv1275 & c1275);
  wire s1276, sub1276, and1276, or1276;
  wire b_inv1276;
  assign b_inv1276 = ~b1276;
  assign s1276  = a1276 ^ b1276 ^ c1276;
  assign sub1276 = a1276 ^ b_inv1276 ^ c1276;
  assign and1276 = a1276 & b1276;
  assign or1276  = a1276 | b1276;
  assign c1277 = (a1276 & b1276) | (a1276 & c1276) | (b1276 & c1276);
  wire c_sub1277;
  assign c_sub1277 = (a1276 & b_inv1276) | (a1276 & c1276) | (b_inv1276 & c1276);
  wire s1277, sub1277, and1277, or1277;
  wire b_inv1277;
  assign b_inv1277 = ~b1277;
  assign s1277  = a1277 ^ b1277 ^ c1277;
  assign sub1277 = a1277 ^ b_inv1277 ^ c1277;
  assign and1277 = a1277 & b1277;
  assign or1277  = a1277 | b1277;
  assign c1278 = (a1277 & b1277) | (a1277 & c1277) | (b1277 & c1277);
  wire c_sub1278;
  assign c_sub1278 = (a1277 & b_inv1277) | (a1277 & c1277) | (b_inv1277 & c1277);
  wire s1278, sub1278, and1278, or1278;
  wire b_inv1278;
  assign b_inv1278 = ~b1278;
  assign s1278  = a1278 ^ b1278 ^ c1278;
  assign sub1278 = a1278 ^ b_inv1278 ^ c1278;
  assign and1278 = a1278 & b1278;
  assign or1278  = a1278 | b1278;
  assign c1279 = (a1278 & b1278) | (a1278 & c1278) | (b1278 & c1278);
  wire c_sub1279;
  assign c_sub1279 = (a1278 & b_inv1278) | (a1278 & c1278) | (b_inv1278 & c1278);
  wire s1279, sub1279, and1279, or1279;
  wire b_inv1279;
  assign b_inv1279 = ~b1279;
  assign s1279  = a1279 ^ b1279 ^ c1279;
  assign sub1279 = a1279 ^ b_inv1279 ^ c1279;
  assign and1279 = a1279 & b1279;
  assign or1279  = a1279 | b1279;
  assign c1280 = (a1279 & b1279) | (a1279 & c1279) | (b1279 & c1279);
  wire c_sub1280;
  assign c_sub1280 = (a1279 & b_inv1279) | (a1279 & c1279) | (b_inv1279 & c1279);
  wire s1280, sub1280, and1280, or1280;
  wire b_inv1280;
  assign b_inv1280 = ~b1280;
  assign s1280  = a1280 ^ b1280 ^ c1280;
  assign sub1280 = a1280 ^ b_inv1280 ^ c1280;
  assign and1280 = a1280 & b1280;
  assign or1280  = a1280 | b1280;
  assign c1281 = (a1280 & b1280) | (a1280 & c1280) | (b1280 & c1280);
  wire c_sub1281;
  assign c_sub1281 = (a1280 & b_inv1280) | (a1280 & c1280) | (b_inv1280 & c1280);
  wire s1281, sub1281, and1281, or1281;
  wire b_inv1281;
  assign b_inv1281 = ~b1281;
  assign s1281  = a1281 ^ b1281 ^ c1281;
  assign sub1281 = a1281 ^ b_inv1281 ^ c1281;
  assign and1281 = a1281 & b1281;
  assign or1281  = a1281 | b1281;
  assign c1282 = (a1281 & b1281) | (a1281 & c1281) | (b1281 & c1281);
  wire c_sub1282;
  assign c_sub1282 = (a1281 & b_inv1281) | (a1281 & c1281) | (b_inv1281 & c1281);
  wire s1282, sub1282, and1282, or1282;
  wire b_inv1282;
  assign b_inv1282 = ~b1282;
  assign s1282  = a1282 ^ b1282 ^ c1282;
  assign sub1282 = a1282 ^ b_inv1282 ^ c1282;
  assign and1282 = a1282 & b1282;
  assign or1282  = a1282 | b1282;
  assign c1283 = (a1282 & b1282) | (a1282 & c1282) | (b1282 & c1282);
  wire c_sub1283;
  assign c_sub1283 = (a1282 & b_inv1282) | (a1282 & c1282) | (b_inv1282 & c1282);
  wire s1283, sub1283, and1283, or1283;
  wire b_inv1283;
  assign b_inv1283 = ~b1283;
  assign s1283  = a1283 ^ b1283 ^ c1283;
  assign sub1283 = a1283 ^ b_inv1283 ^ c1283;
  assign and1283 = a1283 & b1283;
  assign or1283  = a1283 | b1283;
  assign c1284 = (a1283 & b1283) | (a1283 & c1283) | (b1283 & c1283);
  wire c_sub1284;
  assign c_sub1284 = (a1283 & b_inv1283) | (a1283 & c1283) | (b_inv1283 & c1283);
  wire s1284, sub1284, and1284, or1284;
  wire b_inv1284;
  assign b_inv1284 = ~b1284;
  assign s1284  = a1284 ^ b1284 ^ c1284;
  assign sub1284 = a1284 ^ b_inv1284 ^ c1284;
  assign and1284 = a1284 & b1284;
  assign or1284  = a1284 | b1284;
  assign c1285 = (a1284 & b1284) | (a1284 & c1284) | (b1284 & c1284);
  wire c_sub1285;
  assign c_sub1285 = (a1284 & b_inv1284) | (a1284 & c1284) | (b_inv1284 & c1284);
  wire s1285, sub1285, and1285, or1285;
  wire b_inv1285;
  assign b_inv1285 = ~b1285;
  assign s1285  = a1285 ^ b1285 ^ c1285;
  assign sub1285 = a1285 ^ b_inv1285 ^ c1285;
  assign and1285 = a1285 & b1285;
  assign or1285  = a1285 | b1285;
  assign c1286 = (a1285 & b1285) | (a1285 & c1285) | (b1285 & c1285);
  wire c_sub1286;
  assign c_sub1286 = (a1285 & b_inv1285) | (a1285 & c1285) | (b_inv1285 & c1285);
  wire s1286, sub1286, and1286, or1286;
  wire b_inv1286;
  assign b_inv1286 = ~b1286;
  assign s1286  = a1286 ^ b1286 ^ c1286;
  assign sub1286 = a1286 ^ b_inv1286 ^ c1286;
  assign and1286 = a1286 & b1286;
  assign or1286  = a1286 | b1286;
  assign c1287 = (a1286 & b1286) | (a1286 & c1286) | (b1286 & c1286);
  wire c_sub1287;
  assign c_sub1287 = (a1286 & b_inv1286) | (a1286 & c1286) | (b_inv1286 & c1286);
  wire s1287, sub1287, and1287, or1287;
  wire b_inv1287;
  assign b_inv1287 = ~b1287;
  assign s1287  = a1287 ^ b1287 ^ c1287;
  assign sub1287 = a1287 ^ b_inv1287 ^ c1287;
  assign and1287 = a1287 & b1287;
  assign or1287  = a1287 | b1287;
  assign c1288 = (a1287 & b1287) | (a1287 & c1287) | (b1287 & c1287);
  wire c_sub1288;
  assign c_sub1288 = (a1287 & b_inv1287) | (a1287 & c1287) | (b_inv1287 & c1287);
  wire s1288, sub1288, and1288, or1288;
  wire b_inv1288;
  assign b_inv1288 = ~b1288;
  assign s1288  = a1288 ^ b1288 ^ c1288;
  assign sub1288 = a1288 ^ b_inv1288 ^ c1288;
  assign and1288 = a1288 & b1288;
  assign or1288  = a1288 | b1288;
  assign c1289 = (a1288 & b1288) | (a1288 & c1288) | (b1288 & c1288);
  wire c_sub1289;
  assign c_sub1289 = (a1288 & b_inv1288) | (a1288 & c1288) | (b_inv1288 & c1288);
  wire s1289, sub1289, and1289, or1289;
  wire b_inv1289;
  assign b_inv1289 = ~b1289;
  assign s1289  = a1289 ^ b1289 ^ c1289;
  assign sub1289 = a1289 ^ b_inv1289 ^ c1289;
  assign and1289 = a1289 & b1289;
  assign or1289  = a1289 | b1289;
  assign c1290 = (a1289 & b1289) | (a1289 & c1289) | (b1289 & c1289);
  wire c_sub1290;
  assign c_sub1290 = (a1289 & b_inv1289) | (a1289 & c1289) | (b_inv1289 & c1289);
  wire s1290, sub1290, and1290, or1290;
  wire b_inv1290;
  assign b_inv1290 = ~b1290;
  assign s1290  = a1290 ^ b1290 ^ c1290;
  assign sub1290 = a1290 ^ b_inv1290 ^ c1290;
  assign and1290 = a1290 & b1290;
  assign or1290  = a1290 | b1290;
  assign c1291 = (a1290 & b1290) | (a1290 & c1290) | (b1290 & c1290);
  wire c_sub1291;
  assign c_sub1291 = (a1290 & b_inv1290) | (a1290 & c1290) | (b_inv1290 & c1290);
  wire s1291, sub1291, and1291, or1291;
  wire b_inv1291;
  assign b_inv1291 = ~b1291;
  assign s1291  = a1291 ^ b1291 ^ c1291;
  assign sub1291 = a1291 ^ b_inv1291 ^ c1291;
  assign and1291 = a1291 & b1291;
  assign or1291  = a1291 | b1291;
  assign c1292 = (a1291 & b1291) | (a1291 & c1291) | (b1291 & c1291);
  wire c_sub1292;
  assign c_sub1292 = (a1291 & b_inv1291) | (a1291 & c1291) | (b_inv1291 & c1291);
  wire s1292, sub1292, and1292, or1292;
  wire b_inv1292;
  assign b_inv1292 = ~b1292;
  assign s1292  = a1292 ^ b1292 ^ c1292;
  assign sub1292 = a1292 ^ b_inv1292 ^ c1292;
  assign and1292 = a1292 & b1292;
  assign or1292  = a1292 | b1292;
  assign c1293 = (a1292 & b1292) | (a1292 & c1292) | (b1292 & c1292);
  wire c_sub1293;
  assign c_sub1293 = (a1292 & b_inv1292) | (a1292 & c1292) | (b_inv1292 & c1292);
  wire s1293, sub1293, and1293, or1293;
  wire b_inv1293;
  assign b_inv1293 = ~b1293;
  assign s1293  = a1293 ^ b1293 ^ c1293;
  assign sub1293 = a1293 ^ b_inv1293 ^ c1293;
  assign and1293 = a1293 & b1293;
  assign or1293  = a1293 | b1293;
  assign c1294 = (a1293 & b1293) | (a1293 & c1293) | (b1293 & c1293);
  wire c_sub1294;
  assign c_sub1294 = (a1293 & b_inv1293) | (a1293 & c1293) | (b_inv1293 & c1293);
  wire s1294, sub1294, and1294, or1294;
  wire b_inv1294;
  assign b_inv1294 = ~b1294;
  assign s1294  = a1294 ^ b1294 ^ c1294;
  assign sub1294 = a1294 ^ b_inv1294 ^ c1294;
  assign and1294 = a1294 & b1294;
  assign or1294  = a1294 | b1294;
  assign c1295 = (a1294 & b1294) | (a1294 & c1294) | (b1294 & c1294);
  wire c_sub1295;
  assign c_sub1295 = (a1294 & b_inv1294) | (a1294 & c1294) | (b_inv1294 & c1294);
  wire s1295, sub1295, and1295, or1295;
  wire b_inv1295;
  assign b_inv1295 = ~b1295;
  assign s1295  = a1295 ^ b1295 ^ c1295;
  assign sub1295 = a1295 ^ b_inv1295 ^ c1295;
  assign and1295 = a1295 & b1295;
  assign or1295  = a1295 | b1295;
  assign c1296 = (a1295 & b1295) | (a1295 & c1295) | (b1295 & c1295);
  wire c_sub1296;
  assign c_sub1296 = (a1295 & b_inv1295) | (a1295 & c1295) | (b_inv1295 & c1295);
  wire s1296, sub1296, and1296, or1296;
  wire b_inv1296;
  assign b_inv1296 = ~b1296;
  assign s1296  = a1296 ^ b1296 ^ c1296;
  assign sub1296 = a1296 ^ b_inv1296 ^ c1296;
  assign and1296 = a1296 & b1296;
  assign or1296  = a1296 | b1296;
  assign c1297 = (a1296 & b1296) | (a1296 & c1296) | (b1296 & c1296);
  wire c_sub1297;
  assign c_sub1297 = (a1296 & b_inv1296) | (a1296 & c1296) | (b_inv1296 & c1296);
  wire s1297, sub1297, and1297, or1297;
  wire b_inv1297;
  assign b_inv1297 = ~b1297;
  assign s1297  = a1297 ^ b1297 ^ c1297;
  assign sub1297 = a1297 ^ b_inv1297 ^ c1297;
  assign and1297 = a1297 & b1297;
  assign or1297  = a1297 | b1297;
  assign c1298 = (a1297 & b1297) | (a1297 & c1297) | (b1297 & c1297);
  wire c_sub1298;
  assign c_sub1298 = (a1297 & b_inv1297) | (a1297 & c1297) | (b_inv1297 & c1297);
  wire s1298, sub1298, and1298, or1298;
  wire b_inv1298;
  assign b_inv1298 = ~b1298;
  assign s1298  = a1298 ^ b1298 ^ c1298;
  assign sub1298 = a1298 ^ b_inv1298 ^ c1298;
  assign and1298 = a1298 & b1298;
  assign or1298  = a1298 | b1298;
  assign c1299 = (a1298 & b1298) | (a1298 & c1298) | (b1298 & c1298);
  wire c_sub1299;
  assign c_sub1299 = (a1298 & b_inv1298) | (a1298 & c1298) | (b_inv1298 & c1298);
  wire s1299, sub1299, and1299, or1299;
  wire b_inv1299;
  assign b_inv1299 = ~b1299;
  assign s1299  = a1299 ^ b1299 ^ c1299;
  assign sub1299 = a1299 ^ b_inv1299 ^ c1299;
  assign and1299 = a1299 & b1299;
  assign or1299  = a1299 | b1299;
  assign c1300 = (a1299 & b1299) | (a1299 & c1299) | (b1299 & c1299);
  wire c_sub1300;
  assign c_sub1300 = (a1299 & b_inv1299) | (a1299 & c1299) | (b_inv1299 & c1299);
  wire s1300, sub1300, and1300, or1300;
  wire b_inv1300;
  assign b_inv1300 = ~b1300;
  assign s1300  = a1300 ^ b1300 ^ c1300;
  assign sub1300 = a1300 ^ b_inv1300 ^ c1300;
  assign and1300 = a1300 & b1300;
  assign or1300  = a1300 | b1300;
  assign c1301 = (a1300 & b1300) | (a1300 & c1300) | (b1300 & c1300);
  wire c_sub1301;
  assign c_sub1301 = (a1300 & b_inv1300) | (a1300 & c1300) | (b_inv1300 & c1300);
  wire s1301, sub1301, and1301, or1301;
  wire b_inv1301;
  assign b_inv1301 = ~b1301;
  assign s1301  = a1301 ^ b1301 ^ c1301;
  assign sub1301 = a1301 ^ b_inv1301 ^ c1301;
  assign and1301 = a1301 & b1301;
  assign or1301  = a1301 | b1301;
  assign c1302 = (a1301 & b1301) | (a1301 & c1301) | (b1301 & c1301);
  wire c_sub1302;
  assign c_sub1302 = (a1301 & b_inv1301) | (a1301 & c1301) | (b_inv1301 & c1301);
  wire s1302, sub1302, and1302, or1302;
  wire b_inv1302;
  assign b_inv1302 = ~b1302;
  assign s1302  = a1302 ^ b1302 ^ c1302;
  assign sub1302 = a1302 ^ b_inv1302 ^ c1302;
  assign and1302 = a1302 & b1302;
  assign or1302  = a1302 | b1302;
  assign c1303 = (a1302 & b1302) | (a1302 & c1302) | (b1302 & c1302);
  wire c_sub1303;
  assign c_sub1303 = (a1302 & b_inv1302) | (a1302 & c1302) | (b_inv1302 & c1302);
  wire s1303, sub1303, and1303, or1303;
  wire b_inv1303;
  assign b_inv1303 = ~b1303;
  assign s1303  = a1303 ^ b1303 ^ c1303;
  assign sub1303 = a1303 ^ b_inv1303 ^ c1303;
  assign and1303 = a1303 & b1303;
  assign or1303  = a1303 | b1303;
  assign c1304 = (a1303 & b1303) | (a1303 & c1303) | (b1303 & c1303);
  wire c_sub1304;
  assign c_sub1304 = (a1303 & b_inv1303) | (a1303 & c1303) | (b_inv1303 & c1303);
  wire s1304, sub1304, and1304, or1304;
  wire b_inv1304;
  assign b_inv1304 = ~b1304;
  assign s1304  = a1304 ^ b1304 ^ c1304;
  assign sub1304 = a1304 ^ b_inv1304 ^ c1304;
  assign and1304 = a1304 & b1304;
  assign or1304  = a1304 | b1304;
  assign c1305 = (a1304 & b1304) | (a1304 & c1304) | (b1304 & c1304);
  wire c_sub1305;
  assign c_sub1305 = (a1304 & b_inv1304) | (a1304 & c1304) | (b_inv1304 & c1304);
  wire s1305, sub1305, and1305, or1305;
  wire b_inv1305;
  assign b_inv1305 = ~b1305;
  assign s1305  = a1305 ^ b1305 ^ c1305;
  assign sub1305 = a1305 ^ b_inv1305 ^ c1305;
  assign and1305 = a1305 & b1305;
  assign or1305  = a1305 | b1305;
  assign c1306 = (a1305 & b1305) | (a1305 & c1305) | (b1305 & c1305);
  wire c_sub1306;
  assign c_sub1306 = (a1305 & b_inv1305) | (a1305 & c1305) | (b_inv1305 & c1305);
  wire s1306, sub1306, and1306, or1306;
  wire b_inv1306;
  assign b_inv1306 = ~b1306;
  assign s1306  = a1306 ^ b1306 ^ c1306;
  assign sub1306 = a1306 ^ b_inv1306 ^ c1306;
  assign and1306 = a1306 & b1306;
  assign or1306  = a1306 | b1306;
  assign c1307 = (a1306 & b1306) | (a1306 & c1306) | (b1306 & c1306);
  wire c_sub1307;
  assign c_sub1307 = (a1306 & b_inv1306) | (a1306 & c1306) | (b_inv1306 & c1306);
  wire s1307, sub1307, and1307, or1307;
  wire b_inv1307;
  assign b_inv1307 = ~b1307;
  assign s1307  = a1307 ^ b1307 ^ c1307;
  assign sub1307 = a1307 ^ b_inv1307 ^ c1307;
  assign and1307 = a1307 & b1307;
  assign or1307  = a1307 | b1307;
  assign c1308 = (a1307 & b1307) | (a1307 & c1307) | (b1307 & c1307);
  wire c_sub1308;
  assign c_sub1308 = (a1307 & b_inv1307) | (a1307 & c1307) | (b_inv1307 & c1307);
  wire s1308, sub1308, and1308, or1308;
  wire b_inv1308;
  assign b_inv1308 = ~b1308;
  assign s1308  = a1308 ^ b1308 ^ c1308;
  assign sub1308 = a1308 ^ b_inv1308 ^ c1308;
  assign and1308 = a1308 & b1308;
  assign or1308  = a1308 | b1308;
  assign c1309 = (a1308 & b1308) | (a1308 & c1308) | (b1308 & c1308);
  wire c_sub1309;
  assign c_sub1309 = (a1308 & b_inv1308) | (a1308 & c1308) | (b_inv1308 & c1308);
  wire s1309, sub1309, and1309, or1309;
  wire b_inv1309;
  assign b_inv1309 = ~b1309;
  assign s1309  = a1309 ^ b1309 ^ c1309;
  assign sub1309 = a1309 ^ b_inv1309 ^ c1309;
  assign and1309 = a1309 & b1309;
  assign or1309  = a1309 | b1309;
  assign c1310 = (a1309 & b1309) | (a1309 & c1309) | (b1309 & c1309);
  wire c_sub1310;
  assign c_sub1310 = (a1309 & b_inv1309) | (a1309 & c1309) | (b_inv1309 & c1309);
  wire s1310, sub1310, and1310, or1310;
  wire b_inv1310;
  assign b_inv1310 = ~b1310;
  assign s1310  = a1310 ^ b1310 ^ c1310;
  assign sub1310 = a1310 ^ b_inv1310 ^ c1310;
  assign and1310 = a1310 & b1310;
  assign or1310  = a1310 | b1310;
  assign c1311 = (a1310 & b1310) | (a1310 & c1310) | (b1310 & c1310);
  wire c_sub1311;
  assign c_sub1311 = (a1310 & b_inv1310) | (a1310 & c1310) | (b_inv1310 & c1310);
  wire s1311, sub1311, and1311, or1311;
  wire b_inv1311;
  assign b_inv1311 = ~b1311;
  assign s1311  = a1311 ^ b1311 ^ c1311;
  assign sub1311 = a1311 ^ b_inv1311 ^ c1311;
  assign and1311 = a1311 & b1311;
  assign or1311  = a1311 | b1311;
  assign c1312 = (a1311 & b1311) | (a1311 & c1311) | (b1311 & c1311);
  wire c_sub1312;
  assign c_sub1312 = (a1311 & b_inv1311) | (a1311 & c1311) | (b_inv1311 & c1311);
  wire s1312, sub1312, and1312, or1312;
  wire b_inv1312;
  assign b_inv1312 = ~b1312;
  assign s1312  = a1312 ^ b1312 ^ c1312;
  assign sub1312 = a1312 ^ b_inv1312 ^ c1312;
  assign and1312 = a1312 & b1312;
  assign or1312  = a1312 | b1312;
  assign c1313 = (a1312 & b1312) | (a1312 & c1312) | (b1312 & c1312);
  wire c_sub1313;
  assign c_sub1313 = (a1312 & b_inv1312) | (a1312 & c1312) | (b_inv1312 & c1312);
  wire s1313, sub1313, and1313, or1313;
  wire b_inv1313;
  assign b_inv1313 = ~b1313;
  assign s1313  = a1313 ^ b1313 ^ c1313;
  assign sub1313 = a1313 ^ b_inv1313 ^ c1313;
  assign and1313 = a1313 & b1313;
  assign or1313  = a1313 | b1313;
  assign c1314 = (a1313 & b1313) | (a1313 & c1313) | (b1313 & c1313);
  wire c_sub1314;
  assign c_sub1314 = (a1313 & b_inv1313) | (a1313 & c1313) | (b_inv1313 & c1313);
  wire s1314, sub1314, and1314, or1314;
  wire b_inv1314;
  assign b_inv1314 = ~b1314;
  assign s1314  = a1314 ^ b1314 ^ c1314;
  assign sub1314 = a1314 ^ b_inv1314 ^ c1314;
  assign and1314 = a1314 & b1314;
  assign or1314  = a1314 | b1314;
  assign c1315 = (a1314 & b1314) | (a1314 & c1314) | (b1314 & c1314);
  wire c_sub1315;
  assign c_sub1315 = (a1314 & b_inv1314) | (a1314 & c1314) | (b_inv1314 & c1314);
  wire s1315, sub1315, and1315, or1315;
  wire b_inv1315;
  assign b_inv1315 = ~b1315;
  assign s1315  = a1315 ^ b1315 ^ c1315;
  assign sub1315 = a1315 ^ b_inv1315 ^ c1315;
  assign and1315 = a1315 & b1315;
  assign or1315  = a1315 | b1315;
  assign c1316 = (a1315 & b1315) | (a1315 & c1315) | (b1315 & c1315);
  wire c_sub1316;
  assign c_sub1316 = (a1315 & b_inv1315) | (a1315 & c1315) | (b_inv1315 & c1315);
  wire s1316, sub1316, and1316, or1316;
  wire b_inv1316;
  assign b_inv1316 = ~b1316;
  assign s1316  = a1316 ^ b1316 ^ c1316;
  assign sub1316 = a1316 ^ b_inv1316 ^ c1316;
  assign and1316 = a1316 & b1316;
  assign or1316  = a1316 | b1316;
  assign c1317 = (a1316 & b1316) | (a1316 & c1316) | (b1316 & c1316);
  wire c_sub1317;
  assign c_sub1317 = (a1316 & b_inv1316) | (a1316 & c1316) | (b_inv1316 & c1316);
  wire s1317, sub1317, and1317, or1317;
  wire b_inv1317;
  assign b_inv1317 = ~b1317;
  assign s1317  = a1317 ^ b1317 ^ c1317;
  assign sub1317 = a1317 ^ b_inv1317 ^ c1317;
  assign and1317 = a1317 & b1317;
  assign or1317  = a1317 | b1317;
  assign c1318 = (a1317 & b1317) | (a1317 & c1317) | (b1317 & c1317);
  wire c_sub1318;
  assign c_sub1318 = (a1317 & b_inv1317) | (a1317 & c1317) | (b_inv1317 & c1317);
  wire s1318, sub1318, and1318, or1318;
  wire b_inv1318;
  assign b_inv1318 = ~b1318;
  assign s1318  = a1318 ^ b1318 ^ c1318;
  assign sub1318 = a1318 ^ b_inv1318 ^ c1318;
  assign and1318 = a1318 & b1318;
  assign or1318  = a1318 | b1318;
  assign c1319 = (a1318 & b1318) | (a1318 & c1318) | (b1318 & c1318);
  wire c_sub1319;
  assign c_sub1319 = (a1318 & b_inv1318) | (a1318 & c1318) | (b_inv1318 & c1318);
  wire s1319, sub1319, and1319, or1319;
  wire b_inv1319;
  assign b_inv1319 = ~b1319;
  assign s1319  = a1319 ^ b1319 ^ c1319;
  assign sub1319 = a1319 ^ b_inv1319 ^ c1319;
  assign and1319 = a1319 & b1319;
  assign or1319  = a1319 | b1319;
  assign c1320 = (a1319 & b1319) | (a1319 & c1319) | (b1319 & c1319);
  wire c_sub1320;
  assign c_sub1320 = (a1319 & b_inv1319) | (a1319 & c1319) | (b_inv1319 & c1319);
  wire s1320, sub1320, and1320, or1320;
  wire b_inv1320;
  assign b_inv1320 = ~b1320;
  assign s1320  = a1320 ^ b1320 ^ c1320;
  assign sub1320 = a1320 ^ b_inv1320 ^ c1320;
  assign and1320 = a1320 & b1320;
  assign or1320  = a1320 | b1320;
  assign c1321 = (a1320 & b1320) | (a1320 & c1320) | (b1320 & c1320);
  wire c_sub1321;
  assign c_sub1321 = (a1320 & b_inv1320) | (a1320 & c1320) | (b_inv1320 & c1320);
  wire s1321, sub1321, and1321, or1321;
  wire b_inv1321;
  assign b_inv1321 = ~b1321;
  assign s1321  = a1321 ^ b1321 ^ c1321;
  assign sub1321 = a1321 ^ b_inv1321 ^ c1321;
  assign and1321 = a1321 & b1321;
  assign or1321  = a1321 | b1321;
  assign c1322 = (a1321 & b1321) | (a1321 & c1321) | (b1321 & c1321);
  wire c_sub1322;
  assign c_sub1322 = (a1321 & b_inv1321) | (a1321 & c1321) | (b_inv1321 & c1321);
  wire s1322, sub1322, and1322, or1322;
  wire b_inv1322;
  assign b_inv1322 = ~b1322;
  assign s1322  = a1322 ^ b1322 ^ c1322;
  assign sub1322 = a1322 ^ b_inv1322 ^ c1322;
  assign and1322 = a1322 & b1322;
  assign or1322  = a1322 | b1322;
  assign c1323 = (a1322 & b1322) | (a1322 & c1322) | (b1322 & c1322);
  wire c_sub1323;
  assign c_sub1323 = (a1322 & b_inv1322) | (a1322 & c1322) | (b_inv1322 & c1322);
  wire s1323, sub1323, and1323, or1323;
  wire b_inv1323;
  assign b_inv1323 = ~b1323;
  assign s1323  = a1323 ^ b1323 ^ c1323;
  assign sub1323 = a1323 ^ b_inv1323 ^ c1323;
  assign and1323 = a1323 & b1323;
  assign or1323  = a1323 | b1323;
  assign c1324 = (a1323 & b1323) | (a1323 & c1323) | (b1323 & c1323);
  wire c_sub1324;
  assign c_sub1324 = (a1323 & b_inv1323) | (a1323 & c1323) | (b_inv1323 & c1323);
  wire s1324, sub1324, and1324, or1324;
  wire b_inv1324;
  assign b_inv1324 = ~b1324;
  assign s1324  = a1324 ^ b1324 ^ c1324;
  assign sub1324 = a1324 ^ b_inv1324 ^ c1324;
  assign and1324 = a1324 & b1324;
  assign or1324  = a1324 | b1324;
  assign c1325 = (a1324 & b1324) | (a1324 & c1324) | (b1324 & c1324);
  wire c_sub1325;
  assign c_sub1325 = (a1324 & b_inv1324) | (a1324 & c1324) | (b_inv1324 & c1324);
  wire s1325, sub1325, and1325, or1325;
  wire b_inv1325;
  assign b_inv1325 = ~b1325;
  assign s1325  = a1325 ^ b1325 ^ c1325;
  assign sub1325 = a1325 ^ b_inv1325 ^ c1325;
  assign and1325 = a1325 & b1325;
  assign or1325  = a1325 | b1325;
  assign c1326 = (a1325 & b1325) | (a1325 & c1325) | (b1325 & c1325);
  wire c_sub1326;
  assign c_sub1326 = (a1325 & b_inv1325) | (a1325 & c1325) | (b_inv1325 & c1325);
  wire s1326, sub1326, and1326, or1326;
  wire b_inv1326;
  assign b_inv1326 = ~b1326;
  assign s1326  = a1326 ^ b1326 ^ c1326;
  assign sub1326 = a1326 ^ b_inv1326 ^ c1326;
  assign and1326 = a1326 & b1326;
  assign or1326  = a1326 | b1326;
  assign c1327 = (a1326 & b1326) | (a1326 & c1326) | (b1326 & c1326);
  wire c_sub1327;
  assign c_sub1327 = (a1326 & b_inv1326) | (a1326 & c1326) | (b_inv1326 & c1326);
  wire s1327, sub1327, and1327, or1327;
  wire b_inv1327;
  assign b_inv1327 = ~b1327;
  assign s1327  = a1327 ^ b1327 ^ c1327;
  assign sub1327 = a1327 ^ b_inv1327 ^ c1327;
  assign and1327 = a1327 & b1327;
  assign or1327  = a1327 | b1327;
  assign c1328 = (a1327 & b1327) | (a1327 & c1327) | (b1327 & c1327);
  wire c_sub1328;
  assign c_sub1328 = (a1327 & b_inv1327) | (a1327 & c1327) | (b_inv1327 & c1327);
  wire s1328, sub1328, and1328, or1328;
  wire b_inv1328;
  assign b_inv1328 = ~b1328;
  assign s1328  = a1328 ^ b1328 ^ c1328;
  assign sub1328 = a1328 ^ b_inv1328 ^ c1328;
  assign and1328 = a1328 & b1328;
  assign or1328  = a1328 | b1328;
  assign c1329 = (a1328 & b1328) | (a1328 & c1328) | (b1328 & c1328);
  wire c_sub1329;
  assign c_sub1329 = (a1328 & b_inv1328) | (a1328 & c1328) | (b_inv1328 & c1328);
  wire s1329, sub1329, and1329, or1329;
  wire b_inv1329;
  assign b_inv1329 = ~b1329;
  assign s1329  = a1329 ^ b1329 ^ c1329;
  assign sub1329 = a1329 ^ b_inv1329 ^ c1329;
  assign and1329 = a1329 & b1329;
  assign or1329  = a1329 | b1329;
  assign c1330 = (a1329 & b1329) | (a1329 & c1329) | (b1329 & c1329);
  wire c_sub1330;
  assign c_sub1330 = (a1329 & b_inv1329) | (a1329 & c1329) | (b_inv1329 & c1329);
  wire s1330, sub1330, and1330, or1330;
  wire b_inv1330;
  assign b_inv1330 = ~b1330;
  assign s1330  = a1330 ^ b1330 ^ c1330;
  assign sub1330 = a1330 ^ b_inv1330 ^ c1330;
  assign and1330 = a1330 & b1330;
  assign or1330  = a1330 | b1330;
  assign c1331 = (a1330 & b1330) | (a1330 & c1330) | (b1330 & c1330);
  wire c_sub1331;
  assign c_sub1331 = (a1330 & b_inv1330) | (a1330 & c1330) | (b_inv1330 & c1330);
  wire s1331, sub1331, and1331, or1331;
  wire b_inv1331;
  assign b_inv1331 = ~b1331;
  assign s1331  = a1331 ^ b1331 ^ c1331;
  assign sub1331 = a1331 ^ b_inv1331 ^ c1331;
  assign and1331 = a1331 & b1331;
  assign or1331  = a1331 | b1331;
  assign c1332 = (a1331 & b1331) | (a1331 & c1331) | (b1331 & c1331);
  wire c_sub1332;
  assign c_sub1332 = (a1331 & b_inv1331) | (a1331 & c1331) | (b_inv1331 & c1331);
  wire s1332, sub1332, and1332, or1332;
  wire b_inv1332;
  assign b_inv1332 = ~b1332;
  assign s1332  = a1332 ^ b1332 ^ c1332;
  assign sub1332 = a1332 ^ b_inv1332 ^ c1332;
  assign and1332 = a1332 & b1332;
  assign or1332  = a1332 | b1332;
  assign c1333 = (a1332 & b1332) | (a1332 & c1332) | (b1332 & c1332);
  wire c_sub1333;
  assign c_sub1333 = (a1332 & b_inv1332) | (a1332 & c1332) | (b_inv1332 & c1332);
  wire s1333, sub1333, and1333, or1333;
  wire b_inv1333;
  assign b_inv1333 = ~b1333;
  assign s1333  = a1333 ^ b1333 ^ c1333;
  assign sub1333 = a1333 ^ b_inv1333 ^ c1333;
  assign and1333 = a1333 & b1333;
  assign or1333  = a1333 | b1333;
  assign c1334 = (a1333 & b1333) | (a1333 & c1333) | (b1333 & c1333);
  wire c_sub1334;
  assign c_sub1334 = (a1333 & b_inv1333) | (a1333 & c1333) | (b_inv1333 & c1333);
  wire s1334, sub1334, and1334, or1334;
  wire b_inv1334;
  assign b_inv1334 = ~b1334;
  assign s1334  = a1334 ^ b1334 ^ c1334;
  assign sub1334 = a1334 ^ b_inv1334 ^ c1334;
  assign and1334 = a1334 & b1334;
  assign or1334  = a1334 | b1334;
  assign c1335 = (a1334 & b1334) | (a1334 & c1334) | (b1334 & c1334);
  wire c_sub1335;
  assign c_sub1335 = (a1334 & b_inv1334) | (a1334 & c1334) | (b_inv1334 & c1334);
  wire s1335, sub1335, and1335, or1335;
  wire b_inv1335;
  assign b_inv1335 = ~b1335;
  assign s1335  = a1335 ^ b1335 ^ c1335;
  assign sub1335 = a1335 ^ b_inv1335 ^ c1335;
  assign and1335 = a1335 & b1335;
  assign or1335  = a1335 | b1335;
  assign c1336 = (a1335 & b1335) | (a1335 & c1335) | (b1335 & c1335);
  wire c_sub1336;
  assign c_sub1336 = (a1335 & b_inv1335) | (a1335 & c1335) | (b_inv1335 & c1335);
  wire s1336, sub1336, and1336, or1336;
  wire b_inv1336;
  assign b_inv1336 = ~b1336;
  assign s1336  = a1336 ^ b1336 ^ c1336;
  assign sub1336 = a1336 ^ b_inv1336 ^ c1336;
  assign and1336 = a1336 & b1336;
  assign or1336  = a1336 | b1336;
  assign c1337 = (a1336 & b1336) | (a1336 & c1336) | (b1336 & c1336);
  wire c_sub1337;
  assign c_sub1337 = (a1336 & b_inv1336) | (a1336 & c1336) | (b_inv1336 & c1336);
  wire s1337, sub1337, and1337, or1337;
  wire b_inv1337;
  assign b_inv1337 = ~b1337;
  assign s1337  = a1337 ^ b1337 ^ c1337;
  assign sub1337 = a1337 ^ b_inv1337 ^ c1337;
  assign and1337 = a1337 & b1337;
  assign or1337  = a1337 | b1337;
  assign c1338 = (a1337 & b1337) | (a1337 & c1337) | (b1337 & c1337);
  wire c_sub1338;
  assign c_sub1338 = (a1337 & b_inv1337) | (a1337 & c1337) | (b_inv1337 & c1337);
  wire s1338, sub1338, and1338, or1338;
  wire b_inv1338;
  assign b_inv1338 = ~b1338;
  assign s1338  = a1338 ^ b1338 ^ c1338;
  assign sub1338 = a1338 ^ b_inv1338 ^ c1338;
  assign and1338 = a1338 & b1338;
  assign or1338  = a1338 | b1338;
  assign c1339 = (a1338 & b1338) | (a1338 & c1338) | (b1338 & c1338);
  wire c_sub1339;
  assign c_sub1339 = (a1338 & b_inv1338) | (a1338 & c1338) | (b_inv1338 & c1338);
  wire s1339, sub1339, and1339, or1339;
  wire b_inv1339;
  assign b_inv1339 = ~b1339;
  assign s1339  = a1339 ^ b1339 ^ c1339;
  assign sub1339 = a1339 ^ b_inv1339 ^ c1339;
  assign and1339 = a1339 & b1339;
  assign or1339  = a1339 | b1339;
  assign c1340 = (a1339 & b1339) | (a1339 & c1339) | (b1339 & c1339);
  wire c_sub1340;
  assign c_sub1340 = (a1339 & b_inv1339) | (a1339 & c1339) | (b_inv1339 & c1339);
  wire s1340, sub1340, and1340, or1340;
  wire b_inv1340;
  assign b_inv1340 = ~b1340;
  assign s1340  = a1340 ^ b1340 ^ c1340;
  assign sub1340 = a1340 ^ b_inv1340 ^ c1340;
  assign and1340 = a1340 & b1340;
  assign or1340  = a1340 | b1340;
  assign c1341 = (a1340 & b1340) | (a1340 & c1340) | (b1340 & c1340);
  wire c_sub1341;
  assign c_sub1341 = (a1340 & b_inv1340) | (a1340 & c1340) | (b_inv1340 & c1340);
  wire s1341, sub1341, and1341, or1341;
  wire b_inv1341;
  assign b_inv1341 = ~b1341;
  assign s1341  = a1341 ^ b1341 ^ c1341;
  assign sub1341 = a1341 ^ b_inv1341 ^ c1341;
  assign and1341 = a1341 & b1341;
  assign or1341  = a1341 | b1341;
  assign c1342 = (a1341 & b1341) | (a1341 & c1341) | (b1341 & c1341);
  wire c_sub1342;
  assign c_sub1342 = (a1341 & b_inv1341) | (a1341 & c1341) | (b_inv1341 & c1341);
  wire s1342, sub1342, and1342, or1342;
  wire b_inv1342;
  assign b_inv1342 = ~b1342;
  assign s1342  = a1342 ^ b1342 ^ c1342;
  assign sub1342 = a1342 ^ b_inv1342 ^ c1342;
  assign and1342 = a1342 & b1342;
  assign or1342  = a1342 | b1342;
  assign c1343 = (a1342 & b1342) | (a1342 & c1342) | (b1342 & c1342);
  wire c_sub1343;
  assign c_sub1343 = (a1342 & b_inv1342) | (a1342 & c1342) | (b_inv1342 & c1342);
  wire s1343, sub1343, and1343, or1343;
  wire b_inv1343;
  assign b_inv1343 = ~b1343;
  assign s1343  = a1343 ^ b1343 ^ c1343;
  assign sub1343 = a1343 ^ b_inv1343 ^ c1343;
  assign and1343 = a1343 & b1343;
  assign or1343  = a1343 | b1343;
  assign c1344 = (a1343 & b1343) | (a1343 & c1343) | (b1343 & c1343);
  wire c_sub1344;
  assign c_sub1344 = (a1343 & b_inv1343) | (a1343 & c1343) | (b_inv1343 & c1343);
  wire s1344, sub1344, and1344, or1344;
  wire b_inv1344;
  assign b_inv1344 = ~b1344;
  assign s1344  = a1344 ^ b1344 ^ c1344;
  assign sub1344 = a1344 ^ b_inv1344 ^ c1344;
  assign and1344 = a1344 & b1344;
  assign or1344  = a1344 | b1344;
  assign c1345 = (a1344 & b1344) | (a1344 & c1344) | (b1344 & c1344);
  wire c_sub1345;
  assign c_sub1345 = (a1344 & b_inv1344) | (a1344 & c1344) | (b_inv1344 & c1344);
  wire s1345, sub1345, and1345, or1345;
  wire b_inv1345;
  assign b_inv1345 = ~b1345;
  assign s1345  = a1345 ^ b1345 ^ c1345;
  assign sub1345 = a1345 ^ b_inv1345 ^ c1345;
  assign and1345 = a1345 & b1345;
  assign or1345  = a1345 | b1345;
  assign c1346 = (a1345 & b1345) | (a1345 & c1345) | (b1345 & c1345);
  wire c_sub1346;
  assign c_sub1346 = (a1345 & b_inv1345) | (a1345 & c1345) | (b_inv1345 & c1345);
  wire s1346, sub1346, and1346, or1346;
  wire b_inv1346;
  assign b_inv1346 = ~b1346;
  assign s1346  = a1346 ^ b1346 ^ c1346;
  assign sub1346 = a1346 ^ b_inv1346 ^ c1346;
  assign and1346 = a1346 & b1346;
  assign or1346  = a1346 | b1346;
  assign c1347 = (a1346 & b1346) | (a1346 & c1346) | (b1346 & c1346);
  wire c_sub1347;
  assign c_sub1347 = (a1346 & b_inv1346) | (a1346 & c1346) | (b_inv1346 & c1346);
  wire s1347, sub1347, and1347, or1347;
  wire b_inv1347;
  assign b_inv1347 = ~b1347;
  assign s1347  = a1347 ^ b1347 ^ c1347;
  assign sub1347 = a1347 ^ b_inv1347 ^ c1347;
  assign and1347 = a1347 & b1347;
  assign or1347  = a1347 | b1347;
  assign c1348 = (a1347 & b1347) | (a1347 & c1347) | (b1347 & c1347);
  wire c_sub1348;
  assign c_sub1348 = (a1347 & b_inv1347) | (a1347 & c1347) | (b_inv1347 & c1347);
  wire s1348, sub1348, and1348, or1348;
  wire b_inv1348;
  assign b_inv1348 = ~b1348;
  assign s1348  = a1348 ^ b1348 ^ c1348;
  assign sub1348 = a1348 ^ b_inv1348 ^ c1348;
  assign and1348 = a1348 & b1348;
  assign or1348  = a1348 | b1348;
  assign c1349 = (a1348 & b1348) | (a1348 & c1348) | (b1348 & c1348);
  wire c_sub1349;
  assign c_sub1349 = (a1348 & b_inv1348) | (a1348 & c1348) | (b_inv1348 & c1348);
  wire s1349, sub1349, and1349, or1349;
  wire b_inv1349;
  assign b_inv1349 = ~b1349;
  assign s1349  = a1349 ^ b1349 ^ c1349;
  assign sub1349 = a1349 ^ b_inv1349 ^ c1349;
  assign and1349 = a1349 & b1349;
  assign or1349  = a1349 | b1349;
  assign c1350 = (a1349 & b1349) | (a1349 & c1349) | (b1349 & c1349);
  wire c_sub1350;
  assign c_sub1350 = (a1349 & b_inv1349) | (a1349 & c1349) | (b_inv1349 & c1349);
  wire s1350, sub1350, and1350, or1350;
  wire b_inv1350;
  assign b_inv1350 = ~b1350;
  assign s1350  = a1350 ^ b1350 ^ c1350;
  assign sub1350 = a1350 ^ b_inv1350 ^ c1350;
  assign and1350 = a1350 & b1350;
  assign or1350  = a1350 | b1350;
  assign c1351 = (a1350 & b1350) | (a1350 & c1350) | (b1350 & c1350);
  wire c_sub1351;
  assign c_sub1351 = (a1350 & b_inv1350) | (a1350 & c1350) | (b_inv1350 & c1350);
  wire s1351, sub1351, and1351, or1351;
  wire b_inv1351;
  assign b_inv1351 = ~b1351;
  assign s1351  = a1351 ^ b1351 ^ c1351;
  assign sub1351 = a1351 ^ b_inv1351 ^ c1351;
  assign and1351 = a1351 & b1351;
  assign or1351  = a1351 | b1351;
  assign c1352 = (a1351 & b1351) | (a1351 & c1351) | (b1351 & c1351);
  wire c_sub1352;
  assign c_sub1352 = (a1351 & b_inv1351) | (a1351 & c1351) | (b_inv1351 & c1351);
  wire s1352, sub1352, and1352, or1352;
  wire b_inv1352;
  assign b_inv1352 = ~b1352;
  assign s1352  = a1352 ^ b1352 ^ c1352;
  assign sub1352 = a1352 ^ b_inv1352 ^ c1352;
  assign and1352 = a1352 & b1352;
  assign or1352  = a1352 | b1352;
  assign c1353 = (a1352 & b1352) | (a1352 & c1352) | (b1352 & c1352);
  wire c_sub1353;
  assign c_sub1353 = (a1352 & b_inv1352) | (a1352 & c1352) | (b_inv1352 & c1352);
  wire s1353, sub1353, and1353, or1353;
  wire b_inv1353;
  assign b_inv1353 = ~b1353;
  assign s1353  = a1353 ^ b1353 ^ c1353;
  assign sub1353 = a1353 ^ b_inv1353 ^ c1353;
  assign and1353 = a1353 & b1353;
  assign or1353  = a1353 | b1353;
  assign c1354 = (a1353 & b1353) | (a1353 & c1353) | (b1353 & c1353);
  wire c_sub1354;
  assign c_sub1354 = (a1353 & b_inv1353) | (a1353 & c1353) | (b_inv1353 & c1353);
  wire s1354, sub1354, and1354, or1354;
  wire b_inv1354;
  assign b_inv1354 = ~b1354;
  assign s1354  = a1354 ^ b1354 ^ c1354;
  assign sub1354 = a1354 ^ b_inv1354 ^ c1354;
  assign and1354 = a1354 & b1354;
  assign or1354  = a1354 | b1354;
  assign c1355 = (a1354 & b1354) | (a1354 & c1354) | (b1354 & c1354);
  wire c_sub1355;
  assign c_sub1355 = (a1354 & b_inv1354) | (a1354 & c1354) | (b_inv1354 & c1354);
  wire s1355, sub1355, and1355, or1355;
  wire b_inv1355;
  assign b_inv1355 = ~b1355;
  assign s1355  = a1355 ^ b1355 ^ c1355;
  assign sub1355 = a1355 ^ b_inv1355 ^ c1355;
  assign and1355 = a1355 & b1355;
  assign or1355  = a1355 | b1355;
  assign c1356 = (a1355 & b1355) | (a1355 & c1355) | (b1355 & c1355);
  wire c_sub1356;
  assign c_sub1356 = (a1355 & b_inv1355) | (a1355 & c1355) | (b_inv1355 & c1355);
  wire s1356, sub1356, and1356, or1356;
  wire b_inv1356;
  assign b_inv1356 = ~b1356;
  assign s1356  = a1356 ^ b1356 ^ c1356;
  assign sub1356 = a1356 ^ b_inv1356 ^ c1356;
  assign and1356 = a1356 & b1356;
  assign or1356  = a1356 | b1356;
  assign c1357 = (a1356 & b1356) | (a1356 & c1356) | (b1356 & c1356);
  wire c_sub1357;
  assign c_sub1357 = (a1356 & b_inv1356) | (a1356 & c1356) | (b_inv1356 & c1356);
  wire s1357, sub1357, and1357, or1357;
  wire b_inv1357;
  assign b_inv1357 = ~b1357;
  assign s1357  = a1357 ^ b1357 ^ c1357;
  assign sub1357 = a1357 ^ b_inv1357 ^ c1357;
  assign and1357 = a1357 & b1357;
  assign or1357  = a1357 | b1357;
  assign c1358 = (a1357 & b1357) | (a1357 & c1357) | (b1357 & c1357);
  wire c_sub1358;
  assign c_sub1358 = (a1357 & b_inv1357) | (a1357 & c1357) | (b_inv1357 & c1357);
  wire s1358, sub1358, and1358, or1358;
  wire b_inv1358;
  assign b_inv1358 = ~b1358;
  assign s1358  = a1358 ^ b1358 ^ c1358;
  assign sub1358 = a1358 ^ b_inv1358 ^ c1358;
  assign and1358 = a1358 & b1358;
  assign or1358  = a1358 | b1358;
  assign c1359 = (a1358 & b1358) | (a1358 & c1358) | (b1358 & c1358);
  wire c_sub1359;
  assign c_sub1359 = (a1358 & b_inv1358) | (a1358 & c1358) | (b_inv1358 & c1358);
  wire s1359, sub1359, and1359, or1359;
  wire b_inv1359;
  assign b_inv1359 = ~b1359;
  assign s1359  = a1359 ^ b1359 ^ c1359;
  assign sub1359 = a1359 ^ b_inv1359 ^ c1359;
  assign and1359 = a1359 & b1359;
  assign or1359  = a1359 | b1359;
  assign c1360 = (a1359 & b1359) | (a1359 & c1359) | (b1359 & c1359);
  wire c_sub1360;
  assign c_sub1360 = (a1359 & b_inv1359) | (a1359 & c1359) | (b_inv1359 & c1359);
  wire s1360, sub1360, and1360, or1360;
  wire b_inv1360;
  assign b_inv1360 = ~b1360;
  assign s1360  = a1360 ^ b1360 ^ c1360;
  assign sub1360 = a1360 ^ b_inv1360 ^ c1360;
  assign and1360 = a1360 & b1360;
  assign or1360  = a1360 | b1360;
  assign c1361 = (a1360 & b1360) | (a1360 & c1360) | (b1360 & c1360);
  wire c_sub1361;
  assign c_sub1361 = (a1360 & b_inv1360) | (a1360 & c1360) | (b_inv1360 & c1360);
  wire s1361, sub1361, and1361, or1361;
  wire b_inv1361;
  assign b_inv1361 = ~b1361;
  assign s1361  = a1361 ^ b1361 ^ c1361;
  assign sub1361 = a1361 ^ b_inv1361 ^ c1361;
  assign and1361 = a1361 & b1361;
  assign or1361  = a1361 | b1361;
  assign c1362 = (a1361 & b1361) | (a1361 & c1361) | (b1361 & c1361);
  wire c_sub1362;
  assign c_sub1362 = (a1361 & b_inv1361) | (a1361 & c1361) | (b_inv1361 & c1361);
  wire s1362, sub1362, and1362, or1362;
  wire b_inv1362;
  assign b_inv1362 = ~b1362;
  assign s1362  = a1362 ^ b1362 ^ c1362;
  assign sub1362 = a1362 ^ b_inv1362 ^ c1362;
  assign and1362 = a1362 & b1362;
  assign or1362  = a1362 | b1362;
  assign c1363 = (a1362 & b1362) | (a1362 & c1362) | (b1362 & c1362);
  wire c_sub1363;
  assign c_sub1363 = (a1362 & b_inv1362) | (a1362 & c1362) | (b_inv1362 & c1362);
  wire s1363, sub1363, and1363, or1363;
  wire b_inv1363;
  assign b_inv1363 = ~b1363;
  assign s1363  = a1363 ^ b1363 ^ c1363;
  assign sub1363 = a1363 ^ b_inv1363 ^ c1363;
  assign and1363 = a1363 & b1363;
  assign or1363  = a1363 | b1363;
  assign c1364 = (a1363 & b1363) | (a1363 & c1363) | (b1363 & c1363);
  wire c_sub1364;
  assign c_sub1364 = (a1363 & b_inv1363) | (a1363 & c1363) | (b_inv1363 & c1363);
  wire s1364, sub1364, and1364, or1364;
  wire b_inv1364;
  assign b_inv1364 = ~b1364;
  assign s1364  = a1364 ^ b1364 ^ c1364;
  assign sub1364 = a1364 ^ b_inv1364 ^ c1364;
  assign and1364 = a1364 & b1364;
  assign or1364  = a1364 | b1364;
  assign c1365 = (a1364 & b1364) | (a1364 & c1364) | (b1364 & c1364);
  wire c_sub1365;
  assign c_sub1365 = (a1364 & b_inv1364) | (a1364 & c1364) | (b_inv1364 & c1364);
  wire s1365, sub1365, and1365, or1365;
  wire b_inv1365;
  assign b_inv1365 = ~b1365;
  assign s1365  = a1365 ^ b1365 ^ c1365;
  assign sub1365 = a1365 ^ b_inv1365 ^ c1365;
  assign and1365 = a1365 & b1365;
  assign or1365  = a1365 | b1365;
  assign c1366 = (a1365 & b1365) | (a1365 & c1365) | (b1365 & c1365);
  wire c_sub1366;
  assign c_sub1366 = (a1365 & b_inv1365) | (a1365 & c1365) | (b_inv1365 & c1365);
  wire s1366, sub1366, and1366, or1366;
  wire b_inv1366;
  assign b_inv1366 = ~b1366;
  assign s1366  = a1366 ^ b1366 ^ c1366;
  assign sub1366 = a1366 ^ b_inv1366 ^ c1366;
  assign and1366 = a1366 & b1366;
  assign or1366  = a1366 | b1366;
  assign c1367 = (a1366 & b1366) | (a1366 & c1366) | (b1366 & c1366);
  wire c_sub1367;
  assign c_sub1367 = (a1366 & b_inv1366) | (a1366 & c1366) | (b_inv1366 & c1366);
  wire s1367, sub1367, and1367, or1367;
  wire b_inv1367;
  assign b_inv1367 = ~b1367;
  assign s1367  = a1367 ^ b1367 ^ c1367;
  assign sub1367 = a1367 ^ b_inv1367 ^ c1367;
  assign and1367 = a1367 & b1367;
  assign or1367  = a1367 | b1367;
  assign c1368 = (a1367 & b1367) | (a1367 & c1367) | (b1367 & c1367);
  wire c_sub1368;
  assign c_sub1368 = (a1367 & b_inv1367) | (a1367 & c1367) | (b_inv1367 & c1367);
  wire s1368, sub1368, and1368, or1368;
  wire b_inv1368;
  assign b_inv1368 = ~b1368;
  assign s1368  = a1368 ^ b1368 ^ c1368;
  assign sub1368 = a1368 ^ b_inv1368 ^ c1368;
  assign and1368 = a1368 & b1368;
  assign or1368  = a1368 | b1368;
  assign c1369 = (a1368 & b1368) | (a1368 & c1368) | (b1368 & c1368);
  wire c_sub1369;
  assign c_sub1369 = (a1368 & b_inv1368) | (a1368 & c1368) | (b_inv1368 & c1368);
  wire s1369, sub1369, and1369, or1369;
  wire b_inv1369;
  assign b_inv1369 = ~b1369;
  assign s1369  = a1369 ^ b1369 ^ c1369;
  assign sub1369 = a1369 ^ b_inv1369 ^ c1369;
  assign and1369 = a1369 & b1369;
  assign or1369  = a1369 | b1369;
  assign c1370 = (a1369 & b1369) | (a1369 & c1369) | (b1369 & c1369);
  wire c_sub1370;
  assign c_sub1370 = (a1369 & b_inv1369) | (a1369 & c1369) | (b_inv1369 & c1369);
  wire s1370, sub1370, and1370, or1370;
  wire b_inv1370;
  assign b_inv1370 = ~b1370;
  assign s1370  = a1370 ^ b1370 ^ c1370;
  assign sub1370 = a1370 ^ b_inv1370 ^ c1370;
  assign and1370 = a1370 & b1370;
  assign or1370  = a1370 | b1370;
  assign c1371 = (a1370 & b1370) | (a1370 & c1370) | (b1370 & c1370);
  wire c_sub1371;
  assign c_sub1371 = (a1370 & b_inv1370) | (a1370 & c1370) | (b_inv1370 & c1370);
  wire s1371, sub1371, and1371, or1371;
  wire b_inv1371;
  assign b_inv1371 = ~b1371;
  assign s1371  = a1371 ^ b1371 ^ c1371;
  assign sub1371 = a1371 ^ b_inv1371 ^ c1371;
  assign and1371 = a1371 & b1371;
  assign or1371  = a1371 | b1371;
  assign c1372 = (a1371 & b1371) | (a1371 & c1371) | (b1371 & c1371);
  wire c_sub1372;
  assign c_sub1372 = (a1371 & b_inv1371) | (a1371 & c1371) | (b_inv1371 & c1371);
  wire s1372, sub1372, and1372, or1372;
  wire b_inv1372;
  assign b_inv1372 = ~b1372;
  assign s1372  = a1372 ^ b1372 ^ c1372;
  assign sub1372 = a1372 ^ b_inv1372 ^ c1372;
  assign and1372 = a1372 & b1372;
  assign or1372  = a1372 | b1372;
  assign c1373 = (a1372 & b1372) | (a1372 & c1372) | (b1372 & c1372);
  wire c_sub1373;
  assign c_sub1373 = (a1372 & b_inv1372) | (a1372 & c1372) | (b_inv1372 & c1372);
  wire s1373, sub1373, and1373, or1373;
  wire b_inv1373;
  assign b_inv1373 = ~b1373;
  assign s1373  = a1373 ^ b1373 ^ c1373;
  assign sub1373 = a1373 ^ b_inv1373 ^ c1373;
  assign and1373 = a1373 & b1373;
  assign or1373  = a1373 | b1373;
  assign c1374 = (a1373 & b1373) | (a1373 & c1373) | (b1373 & c1373);
  wire c_sub1374;
  assign c_sub1374 = (a1373 & b_inv1373) | (a1373 & c1373) | (b_inv1373 & c1373);
  wire s1374, sub1374, and1374, or1374;
  wire b_inv1374;
  assign b_inv1374 = ~b1374;
  assign s1374  = a1374 ^ b1374 ^ c1374;
  assign sub1374 = a1374 ^ b_inv1374 ^ c1374;
  assign and1374 = a1374 & b1374;
  assign or1374  = a1374 | b1374;
  assign c1375 = (a1374 & b1374) | (a1374 & c1374) | (b1374 & c1374);
  wire c_sub1375;
  assign c_sub1375 = (a1374 & b_inv1374) | (a1374 & c1374) | (b_inv1374 & c1374);
  wire s1375, sub1375, and1375, or1375;
  wire b_inv1375;
  assign b_inv1375 = ~b1375;
  assign s1375  = a1375 ^ b1375 ^ c1375;
  assign sub1375 = a1375 ^ b_inv1375 ^ c1375;
  assign and1375 = a1375 & b1375;
  assign or1375  = a1375 | b1375;
  assign c1376 = (a1375 & b1375) | (a1375 & c1375) | (b1375 & c1375);
  wire c_sub1376;
  assign c_sub1376 = (a1375 & b_inv1375) | (a1375 & c1375) | (b_inv1375 & c1375);
  wire s1376, sub1376, and1376, or1376;
  wire b_inv1376;
  assign b_inv1376 = ~b1376;
  assign s1376  = a1376 ^ b1376 ^ c1376;
  assign sub1376 = a1376 ^ b_inv1376 ^ c1376;
  assign and1376 = a1376 & b1376;
  assign or1376  = a1376 | b1376;
  assign c1377 = (a1376 & b1376) | (a1376 & c1376) | (b1376 & c1376);
  wire c_sub1377;
  assign c_sub1377 = (a1376 & b_inv1376) | (a1376 & c1376) | (b_inv1376 & c1376);
  wire s1377, sub1377, and1377, or1377;
  wire b_inv1377;
  assign b_inv1377 = ~b1377;
  assign s1377  = a1377 ^ b1377 ^ c1377;
  assign sub1377 = a1377 ^ b_inv1377 ^ c1377;
  assign and1377 = a1377 & b1377;
  assign or1377  = a1377 | b1377;
  assign c1378 = (a1377 & b1377) | (a1377 & c1377) | (b1377 & c1377);
  wire c_sub1378;
  assign c_sub1378 = (a1377 & b_inv1377) | (a1377 & c1377) | (b_inv1377 & c1377);
  wire s1378, sub1378, and1378, or1378;
  wire b_inv1378;
  assign b_inv1378 = ~b1378;
  assign s1378  = a1378 ^ b1378 ^ c1378;
  assign sub1378 = a1378 ^ b_inv1378 ^ c1378;
  assign and1378 = a1378 & b1378;
  assign or1378  = a1378 | b1378;
  assign c1379 = (a1378 & b1378) | (a1378 & c1378) | (b1378 & c1378);
  wire c_sub1379;
  assign c_sub1379 = (a1378 & b_inv1378) | (a1378 & c1378) | (b_inv1378 & c1378);
  wire s1379, sub1379, and1379, or1379;
  wire b_inv1379;
  assign b_inv1379 = ~b1379;
  assign s1379  = a1379 ^ b1379 ^ c1379;
  assign sub1379 = a1379 ^ b_inv1379 ^ c1379;
  assign and1379 = a1379 & b1379;
  assign or1379  = a1379 | b1379;
  assign c1380 = (a1379 & b1379) | (a1379 & c1379) | (b1379 & c1379);
  wire c_sub1380;
  assign c_sub1380 = (a1379 & b_inv1379) | (a1379 & c1379) | (b_inv1379 & c1379);
  wire s1380, sub1380, and1380, or1380;
  wire b_inv1380;
  assign b_inv1380 = ~b1380;
  assign s1380  = a1380 ^ b1380 ^ c1380;
  assign sub1380 = a1380 ^ b_inv1380 ^ c1380;
  assign and1380 = a1380 & b1380;
  assign or1380  = a1380 | b1380;
  assign c1381 = (a1380 & b1380) | (a1380 & c1380) | (b1380 & c1380);
  wire c_sub1381;
  assign c_sub1381 = (a1380 & b_inv1380) | (a1380 & c1380) | (b_inv1380 & c1380);
  wire s1381, sub1381, and1381, or1381;
  wire b_inv1381;
  assign b_inv1381 = ~b1381;
  assign s1381  = a1381 ^ b1381 ^ c1381;
  assign sub1381 = a1381 ^ b_inv1381 ^ c1381;
  assign and1381 = a1381 & b1381;
  assign or1381  = a1381 | b1381;
  assign c1382 = (a1381 & b1381) | (a1381 & c1381) | (b1381 & c1381);
  wire c_sub1382;
  assign c_sub1382 = (a1381 & b_inv1381) | (a1381 & c1381) | (b_inv1381 & c1381);
  wire s1382, sub1382, and1382, or1382;
  wire b_inv1382;
  assign b_inv1382 = ~b1382;
  assign s1382  = a1382 ^ b1382 ^ c1382;
  assign sub1382 = a1382 ^ b_inv1382 ^ c1382;
  assign and1382 = a1382 & b1382;
  assign or1382  = a1382 | b1382;
  assign c1383 = (a1382 & b1382) | (a1382 & c1382) | (b1382 & c1382);
  wire c_sub1383;
  assign c_sub1383 = (a1382 & b_inv1382) | (a1382 & c1382) | (b_inv1382 & c1382);
  wire s1383, sub1383, and1383, or1383;
  wire b_inv1383;
  assign b_inv1383 = ~b1383;
  assign s1383  = a1383 ^ b1383 ^ c1383;
  assign sub1383 = a1383 ^ b_inv1383 ^ c1383;
  assign and1383 = a1383 & b1383;
  assign or1383  = a1383 | b1383;
  assign c1384 = (a1383 & b1383) | (a1383 & c1383) | (b1383 & c1383);
  wire c_sub1384;
  assign c_sub1384 = (a1383 & b_inv1383) | (a1383 & c1383) | (b_inv1383 & c1383);
  wire s1384, sub1384, and1384, or1384;
  wire b_inv1384;
  assign b_inv1384 = ~b1384;
  assign s1384  = a1384 ^ b1384 ^ c1384;
  assign sub1384 = a1384 ^ b_inv1384 ^ c1384;
  assign and1384 = a1384 & b1384;
  assign or1384  = a1384 | b1384;
  assign c1385 = (a1384 & b1384) | (a1384 & c1384) | (b1384 & c1384);
  wire c_sub1385;
  assign c_sub1385 = (a1384 & b_inv1384) | (a1384 & c1384) | (b_inv1384 & c1384);
  wire s1385, sub1385, and1385, or1385;
  wire b_inv1385;
  assign b_inv1385 = ~b1385;
  assign s1385  = a1385 ^ b1385 ^ c1385;
  assign sub1385 = a1385 ^ b_inv1385 ^ c1385;
  assign and1385 = a1385 & b1385;
  assign or1385  = a1385 | b1385;
  assign c1386 = (a1385 & b1385) | (a1385 & c1385) | (b1385 & c1385);
  wire c_sub1386;
  assign c_sub1386 = (a1385 & b_inv1385) | (a1385 & c1385) | (b_inv1385 & c1385);
  wire s1386, sub1386, and1386, or1386;
  wire b_inv1386;
  assign b_inv1386 = ~b1386;
  assign s1386  = a1386 ^ b1386 ^ c1386;
  assign sub1386 = a1386 ^ b_inv1386 ^ c1386;
  assign and1386 = a1386 & b1386;
  assign or1386  = a1386 | b1386;
  assign c1387 = (a1386 & b1386) | (a1386 & c1386) | (b1386 & c1386);
  wire c_sub1387;
  assign c_sub1387 = (a1386 & b_inv1386) | (a1386 & c1386) | (b_inv1386 & c1386);
  wire s1387, sub1387, and1387, or1387;
  wire b_inv1387;
  assign b_inv1387 = ~b1387;
  assign s1387  = a1387 ^ b1387 ^ c1387;
  assign sub1387 = a1387 ^ b_inv1387 ^ c1387;
  assign and1387 = a1387 & b1387;
  assign or1387  = a1387 | b1387;
  assign c1388 = (a1387 & b1387) | (a1387 & c1387) | (b1387 & c1387);
  wire c_sub1388;
  assign c_sub1388 = (a1387 & b_inv1387) | (a1387 & c1387) | (b_inv1387 & c1387);
  wire s1388, sub1388, and1388, or1388;
  wire b_inv1388;
  assign b_inv1388 = ~b1388;
  assign s1388  = a1388 ^ b1388 ^ c1388;
  assign sub1388 = a1388 ^ b_inv1388 ^ c1388;
  assign and1388 = a1388 & b1388;
  assign or1388  = a1388 | b1388;
  assign c1389 = (a1388 & b1388) | (a1388 & c1388) | (b1388 & c1388);
  wire c_sub1389;
  assign c_sub1389 = (a1388 & b_inv1388) | (a1388 & c1388) | (b_inv1388 & c1388);
  wire s1389, sub1389, and1389, or1389;
  wire b_inv1389;
  assign b_inv1389 = ~b1389;
  assign s1389  = a1389 ^ b1389 ^ c1389;
  assign sub1389 = a1389 ^ b_inv1389 ^ c1389;
  assign and1389 = a1389 & b1389;
  assign or1389  = a1389 | b1389;
  assign c1390 = (a1389 & b1389) | (a1389 & c1389) | (b1389 & c1389);
  wire c_sub1390;
  assign c_sub1390 = (a1389 & b_inv1389) | (a1389 & c1389) | (b_inv1389 & c1389);
  wire s1390, sub1390, and1390, or1390;
  wire b_inv1390;
  assign b_inv1390 = ~b1390;
  assign s1390  = a1390 ^ b1390 ^ c1390;
  assign sub1390 = a1390 ^ b_inv1390 ^ c1390;
  assign and1390 = a1390 & b1390;
  assign or1390  = a1390 | b1390;
  assign c1391 = (a1390 & b1390) | (a1390 & c1390) | (b1390 & c1390);
  wire c_sub1391;
  assign c_sub1391 = (a1390 & b_inv1390) | (a1390 & c1390) | (b_inv1390 & c1390);
  wire s1391, sub1391, and1391, or1391;
  wire b_inv1391;
  assign b_inv1391 = ~b1391;
  assign s1391  = a1391 ^ b1391 ^ c1391;
  assign sub1391 = a1391 ^ b_inv1391 ^ c1391;
  assign and1391 = a1391 & b1391;
  assign or1391  = a1391 | b1391;
  assign c1392 = (a1391 & b1391) | (a1391 & c1391) | (b1391 & c1391);
  wire c_sub1392;
  assign c_sub1392 = (a1391 & b_inv1391) | (a1391 & c1391) | (b_inv1391 & c1391);
  wire s1392, sub1392, and1392, or1392;
  wire b_inv1392;
  assign b_inv1392 = ~b1392;
  assign s1392  = a1392 ^ b1392 ^ c1392;
  assign sub1392 = a1392 ^ b_inv1392 ^ c1392;
  assign and1392 = a1392 & b1392;
  assign or1392  = a1392 | b1392;
  assign c1393 = (a1392 & b1392) | (a1392 & c1392) | (b1392 & c1392);
  wire c_sub1393;
  assign c_sub1393 = (a1392 & b_inv1392) | (a1392 & c1392) | (b_inv1392 & c1392);
  wire s1393, sub1393, and1393, or1393;
  wire b_inv1393;
  assign b_inv1393 = ~b1393;
  assign s1393  = a1393 ^ b1393 ^ c1393;
  assign sub1393 = a1393 ^ b_inv1393 ^ c1393;
  assign and1393 = a1393 & b1393;
  assign or1393  = a1393 | b1393;
  assign c1394 = (a1393 & b1393) | (a1393 & c1393) | (b1393 & c1393);
  wire c_sub1394;
  assign c_sub1394 = (a1393 & b_inv1393) | (a1393 & c1393) | (b_inv1393 & c1393);
  wire s1394, sub1394, and1394, or1394;
  wire b_inv1394;
  assign b_inv1394 = ~b1394;
  assign s1394  = a1394 ^ b1394 ^ c1394;
  assign sub1394 = a1394 ^ b_inv1394 ^ c1394;
  assign and1394 = a1394 & b1394;
  assign or1394  = a1394 | b1394;
  assign c1395 = (a1394 & b1394) | (a1394 & c1394) | (b1394 & c1394);
  wire c_sub1395;
  assign c_sub1395 = (a1394 & b_inv1394) | (a1394 & c1394) | (b_inv1394 & c1394);
  wire s1395, sub1395, and1395, or1395;
  wire b_inv1395;
  assign b_inv1395 = ~b1395;
  assign s1395  = a1395 ^ b1395 ^ c1395;
  assign sub1395 = a1395 ^ b_inv1395 ^ c1395;
  assign and1395 = a1395 & b1395;
  assign or1395  = a1395 | b1395;
  assign c1396 = (a1395 & b1395) | (a1395 & c1395) | (b1395 & c1395);
  wire c_sub1396;
  assign c_sub1396 = (a1395 & b_inv1395) | (a1395 & c1395) | (b_inv1395 & c1395);
  wire s1396, sub1396, and1396, or1396;
  wire b_inv1396;
  assign b_inv1396 = ~b1396;
  assign s1396  = a1396 ^ b1396 ^ c1396;
  assign sub1396 = a1396 ^ b_inv1396 ^ c1396;
  assign and1396 = a1396 & b1396;
  assign or1396  = a1396 | b1396;
  assign c1397 = (a1396 & b1396) | (a1396 & c1396) | (b1396 & c1396);
  wire c_sub1397;
  assign c_sub1397 = (a1396 & b_inv1396) | (a1396 & c1396) | (b_inv1396 & c1396);
  wire s1397, sub1397, and1397, or1397;
  wire b_inv1397;
  assign b_inv1397 = ~b1397;
  assign s1397  = a1397 ^ b1397 ^ c1397;
  assign sub1397 = a1397 ^ b_inv1397 ^ c1397;
  assign and1397 = a1397 & b1397;
  assign or1397  = a1397 | b1397;
  assign c1398 = (a1397 & b1397) | (a1397 & c1397) | (b1397 & c1397);
  wire c_sub1398;
  assign c_sub1398 = (a1397 & b_inv1397) | (a1397 & c1397) | (b_inv1397 & c1397);
  wire s1398, sub1398, and1398, or1398;
  wire b_inv1398;
  assign b_inv1398 = ~b1398;
  assign s1398  = a1398 ^ b1398 ^ c1398;
  assign sub1398 = a1398 ^ b_inv1398 ^ c1398;
  assign and1398 = a1398 & b1398;
  assign or1398  = a1398 | b1398;
  assign c1399 = (a1398 & b1398) | (a1398 & c1398) | (b1398 & c1398);
  wire c_sub1399;
  assign c_sub1399 = (a1398 & b_inv1398) | (a1398 & c1398) | (b_inv1398 & c1398);
  wire s1399, sub1399, and1399, or1399;
  wire b_inv1399;
  assign b_inv1399 = ~b1399;
  assign s1399  = a1399 ^ b1399 ^ c1399;
  assign sub1399 = a1399 ^ b_inv1399 ^ c1399;
  assign and1399 = a1399 & b1399;
  assign or1399  = a1399 | b1399;
  assign c1400 = (a1399 & b1399) | (a1399 & c1399) | (b1399 & c1399);
  wire c_sub1400;
  assign c_sub1400 = (a1399 & b_inv1399) | (a1399 & c1399) | (b_inv1399 & c1399);
  wire s1400, sub1400, and1400, or1400;
  wire b_inv1400;
  assign b_inv1400 = ~b1400;
  assign s1400  = a1400 ^ b1400 ^ c1400;
  assign sub1400 = a1400 ^ b_inv1400 ^ c1400;
  assign and1400 = a1400 & b1400;
  assign or1400  = a1400 | b1400;
  assign c1401 = (a1400 & b1400) | (a1400 & c1400) | (b1400 & c1400);
  wire c_sub1401;
  assign c_sub1401 = (a1400 & b_inv1400) | (a1400 & c1400) | (b_inv1400 & c1400);
  wire s1401, sub1401, and1401, or1401;
  wire b_inv1401;
  assign b_inv1401 = ~b1401;
  assign s1401  = a1401 ^ b1401 ^ c1401;
  assign sub1401 = a1401 ^ b_inv1401 ^ c1401;
  assign and1401 = a1401 & b1401;
  assign or1401  = a1401 | b1401;
  assign c1402 = (a1401 & b1401) | (a1401 & c1401) | (b1401 & c1401);
  wire c_sub1402;
  assign c_sub1402 = (a1401 & b_inv1401) | (a1401 & c1401) | (b_inv1401 & c1401);
  wire s1402, sub1402, and1402, or1402;
  wire b_inv1402;
  assign b_inv1402 = ~b1402;
  assign s1402  = a1402 ^ b1402 ^ c1402;
  assign sub1402 = a1402 ^ b_inv1402 ^ c1402;
  assign and1402 = a1402 & b1402;
  assign or1402  = a1402 | b1402;
  assign c1403 = (a1402 & b1402) | (a1402 & c1402) | (b1402 & c1402);
  wire c_sub1403;
  assign c_sub1403 = (a1402 & b_inv1402) | (a1402 & c1402) | (b_inv1402 & c1402);
  wire s1403, sub1403, and1403, or1403;
  wire b_inv1403;
  assign b_inv1403 = ~b1403;
  assign s1403  = a1403 ^ b1403 ^ c1403;
  assign sub1403 = a1403 ^ b_inv1403 ^ c1403;
  assign and1403 = a1403 & b1403;
  assign or1403  = a1403 | b1403;
  assign c1404 = (a1403 & b1403) | (a1403 & c1403) | (b1403 & c1403);
  wire c_sub1404;
  assign c_sub1404 = (a1403 & b_inv1403) | (a1403 & c1403) | (b_inv1403 & c1403);
  wire s1404, sub1404, and1404, or1404;
  wire b_inv1404;
  assign b_inv1404 = ~b1404;
  assign s1404  = a1404 ^ b1404 ^ c1404;
  assign sub1404 = a1404 ^ b_inv1404 ^ c1404;
  assign and1404 = a1404 & b1404;
  assign or1404  = a1404 | b1404;
  assign c1405 = (a1404 & b1404) | (a1404 & c1404) | (b1404 & c1404);
  wire c_sub1405;
  assign c_sub1405 = (a1404 & b_inv1404) | (a1404 & c1404) | (b_inv1404 & c1404);
  wire s1405, sub1405, and1405, or1405;
  wire b_inv1405;
  assign b_inv1405 = ~b1405;
  assign s1405  = a1405 ^ b1405 ^ c1405;
  assign sub1405 = a1405 ^ b_inv1405 ^ c1405;
  assign and1405 = a1405 & b1405;
  assign or1405  = a1405 | b1405;
  assign c1406 = (a1405 & b1405) | (a1405 & c1405) | (b1405 & c1405);
  wire c_sub1406;
  assign c_sub1406 = (a1405 & b_inv1405) | (a1405 & c1405) | (b_inv1405 & c1405);
  wire s1406, sub1406, and1406, or1406;
  wire b_inv1406;
  assign b_inv1406 = ~b1406;
  assign s1406  = a1406 ^ b1406 ^ c1406;
  assign sub1406 = a1406 ^ b_inv1406 ^ c1406;
  assign and1406 = a1406 & b1406;
  assign or1406  = a1406 | b1406;
  assign c1407 = (a1406 & b1406) | (a1406 & c1406) | (b1406 & c1406);
  wire c_sub1407;
  assign c_sub1407 = (a1406 & b_inv1406) | (a1406 & c1406) | (b_inv1406 & c1406);
  wire s1407, sub1407, and1407, or1407;
  wire b_inv1407;
  assign b_inv1407 = ~b1407;
  assign s1407  = a1407 ^ b1407 ^ c1407;
  assign sub1407 = a1407 ^ b_inv1407 ^ c1407;
  assign and1407 = a1407 & b1407;
  assign or1407  = a1407 | b1407;
  assign c1408 = (a1407 & b1407) | (a1407 & c1407) | (b1407 & c1407);
  wire c_sub1408;
  assign c_sub1408 = (a1407 & b_inv1407) | (a1407 & c1407) | (b_inv1407 & c1407);
  wire s1408, sub1408, and1408, or1408;
  wire b_inv1408;
  assign b_inv1408 = ~b1408;
  assign s1408  = a1408 ^ b1408 ^ c1408;
  assign sub1408 = a1408 ^ b_inv1408 ^ c1408;
  assign and1408 = a1408 & b1408;
  assign or1408  = a1408 | b1408;
  assign c1409 = (a1408 & b1408) | (a1408 & c1408) | (b1408 & c1408);
  wire c_sub1409;
  assign c_sub1409 = (a1408 & b_inv1408) | (a1408 & c1408) | (b_inv1408 & c1408);
  wire s1409, sub1409, and1409, or1409;
  wire b_inv1409;
  assign b_inv1409 = ~b1409;
  assign s1409  = a1409 ^ b1409 ^ c1409;
  assign sub1409 = a1409 ^ b_inv1409 ^ c1409;
  assign and1409 = a1409 & b1409;
  assign or1409  = a1409 | b1409;
  assign c1410 = (a1409 & b1409) | (a1409 & c1409) | (b1409 & c1409);
  wire c_sub1410;
  assign c_sub1410 = (a1409 & b_inv1409) | (a1409 & c1409) | (b_inv1409 & c1409);
  wire s1410, sub1410, and1410, or1410;
  wire b_inv1410;
  assign b_inv1410 = ~b1410;
  assign s1410  = a1410 ^ b1410 ^ c1410;
  assign sub1410 = a1410 ^ b_inv1410 ^ c1410;
  assign and1410 = a1410 & b1410;
  assign or1410  = a1410 | b1410;
  assign c1411 = (a1410 & b1410) | (a1410 & c1410) | (b1410 & c1410);
  wire c_sub1411;
  assign c_sub1411 = (a1410 & b_inv1410) | (a1410 & c1410) | (b_inv1410 & c1410);
  wire s1411, sub1411, and1411, or1411;
  wire b_inv1411;
  assign b_inv1411 = ~b1411;
  assign s1411  = a1411 ^ b1411 ^ c1411;
  assign sub1411 = a1411 ^ b_inv1411 ^ c1411;
  assign and1411 = a1411 & b1411;
  assign or1411  = a1411 | b1411;
  assign c1412 = (a1411 & b1411) | (a1411 & c1411) | (b1411 & c1411);
  wire c_sub1412;
  assign c_sub1412 = (a1411 & b_inv1411) | (a1411 & c1411) | (b_inv1411 & c1411);
  wire s1412, sub1412, and1412, or1412;
  wire b_inv1412;
  assign b_inv1412 = ~b1412;
  assign s1412  = a1412 ^ b1412 ^ c1412;
  assign sub1412 = a1412 ^ b_inv1412 ^ c1412;
  assign and1412 = a1412 & b1412;
  assign or1412  = a1412 | b1412;
  assign c1413 = (a1412 & b1412) | (a1412 & c1412) | (b1412 & c1412);
  wire c_sub1413;
  assign c_sub1413 = (a1412 & b_inv1412) | (a1412 & c1412) | (b_inv1412 & c1412);
  wire s1413, sub1413, and1413, or1413;
  wire b_inv1413;
  assign b_inv1413 = ~b1413;
  assign s1413  = a1413 ^ b1413 ^ c1413;
  assign sub1413 = a1413 ^ b_inv1413 ^ c1413;
  assign and1413 = a1413 & b1413;
  assign or1413  = a1413 | b1413;
  assign c1414 = (a1413 & b1413) | (a1413 & c1413) | (b1413 & c1413);
  wire c_sub1414;
  assign c_sub1414 = (a1413 & b_inv1413) | (a1413 & c1413) | (b_inv1413 & c1413);
  wire s1414, sub1414, and1414, or1414;
  wire b_inv1414;
  assign b_inv1414 = ~b1414;
  assign s1414  = a1414 ^ b1414 ^ c1414;
  assign sub1414 = a1414 ^ b_inv1414 ^ c1414;
  assign and1414 = a1414 & b1414;
  assign or1414  = a1414 | b1414;
  assign c1415 = (a1414 & b1414) | (a1414 & c1414) | (b1414 & c1414);
  wire c_sub1415;
  assign c_sub1415 = (a1414 & b_inv1414) | (a1414 & c1414) | (b_inv1414 & c1414);
  wire s1415, sub1415, and1415, or1415;
  wire b_inv1415;
  assign b_inv1415 = ~b1415;
  assign s1415  = a1415 ^ b1415 ^ c1415;
  assign sub1415 = a1415 ^ b_inv1415 ^ c1415;
  assign and1415 = a1415 & b1415;
  assign or1415  = a1415 | b1415;
  assign c1416 = (a1415 & b1415) | (a1415 & c1415) | (b1415 & c1415);
  wire c_sub1416;
  assign c_sub1416 = (a1415 & b_inv1415) | (a1415 & c1415) | (b_inv1415 & c1415);
  wire s1416, sub1416, and1416, or1416;
  wire b_inv1416;
  assign b_inv1416 = ~b1416;
  assign s1416  = a1416 ^ b1416 ^ c1416;
  assign sub1416 = a1416 ^ b_inv1416 ^ c1416;
  assign and1416 = a1416 & b1416;
  assign or1416  = a1416 | b1416;
  assign c1417 = (a1416 & b1416) | (a1416 & c1416) | (b1416 & c1416);
  wire c_sub1417;
  assign c_sub1417 = (a1416 & b_inv1416) | (a1416 & c1416) | (b_inv1416 & c1416);
  wire s1417, sub1417, and1417, or1417;
  wire b_inv1417;
  assign b_inv1417 = ~b1417;
  assign s1417  = a1417 ^ b1417 ^ c1417;
  assign sub1417 = a1417 ^ b_inv1417 ^ c1417;
  assign and1417 = a1417 & b1417;
  assign or1417  = a1417 | b1417;
  assign c1418 = (a1417 & b1417) | (a1417 & c1417) | (b1417 & c1417);
  wire c_sub1418;
  assign c_sub1418 = (a1417 & b_inv1417) | (a1417 & c1417) | (b_inv1417 & c1417);
  wire s1418, sub1418, and1418, or1418;
  wire b_inv1418;
  assign b_inv1418 = ~b1418;
  assign s1418  = a1418 ^ b1418 ^ c1418;
  assign sub1418 = a1418 ^ b_inv1418 ^ c1418;
  assign and1418 = a1418 & b1418;
  assign or1418  = a1418 | b1418;
  assign c1419 = (a1418 & b1418) | (a1418 & c1418) | (b1418 & c1418);
  wire c_sub1419;
  assign c_sub1419 = (a1418 & b_inv1418) | (a1418 & c1418) | (b_inv1418 & c1418);
  wire s1419, sub1419, and1419, or1419;
  wire b_inv1419;
  assign b_inv1419 = ~b1419;
  assign s1419  = a1419 ^ b1419 ^ c1419;
  assign sub1419 = a1419 ^ b_inv1419 ^ c1419;
  assign and1419 = a1419 & b1419;
  assign or1419  = a1419 | b1419;
  assign c1420 = (a1419 & b1419) | (a1419 & c1419) | (b1419 & c1419);
  wire c_sub1420;
  assign c_sub1420 = (a1419 & b_inv1419) | (a1419 & c1419) | (b_inv1419 & c1419);
  wire s1420, sub1420, and1420, or1420;
  wire b_inv1420;
  assign b_inv1420 = ~b1420;
  assign s1420  = a1420 ^ b1420 ^ c1420;
  assign sub1420 = a1420 ^ b_inv1420 ^ c1420;
  assign and1420 = a1420 & b1420;
  assign or1420  = a1420 | b1420;
  assign c1421 = (a1420 & b1420) | (a1420 & c1420) | (b1420 & c1420);
  wire c_sub1421;
  assign c_sub1421 = (a1420 & b_inv1420) | (a1420 & c1420) | (b_inv1420 & c1420);
  wire s1421, sub1421, and1421, or1421;
  wire b_inv1421;
  assign b_inv1421 = ~b1421;
  assign s1421  = a1421 ^ b1421 ^ c1421;
  assign sub1421 = a1421 ^ b_inv1421 ^ c1421;
  assign and1421 = a1421 & b1421;
  assign or1421  = a1421 | b1421;
  assign c1422 = (a1421 & b1421) | (a1421 & c1421) | (b1421 & c1421);
  wire c_sub1422;
  assign c_sub1422 = (a1421 & b_inv1421) | (a1421 & c1421) | (b_inv1421 & c1421);
  wire s1422, sub1422, and1422, or1422;
  wire b_inv1422;
  assign b_inv1422 = ~b1422;
  assign s1422  = a1422 ^ b1422 ^ c1422;
  assign sub1422 = a1422 ^ b_inv1422 ^ c1422;
  assign and1422 = a1422 & b1422;
  assign or1422  = a1422 | b1422;
  assign c1423 = (a1422 & b1422) | (a1422 & c1422) | (b1422 & c1422);
  wire c_sub1423;
  assign c_sub1423 = (a1422 & b_inv1422) | (a1422 & c1422) | (b_inv1422 & c1422);
  wire s1423, sub1423, and1423, or1423;
  wire b_inv1423;
  assign b_inv1423 = ~b1423;
  assign s1423  = a1423 ^ b1423 ^ c1423;
  assign sub1423 = a1423 ^ b_inv1423 ^ c1423;
  assign and1423 = a1423 & b1423;
  assign or1423  = a1423 | b1423;
  assign c1424 = (a1423 & b1423) | (a1423 & c1423) | (b1423 & c1423);
  wire c_sub1424;
  assign c_sub1424 = (a1423 & b_inv1423) | (a1423 & c1423) | (b_inv1423 & c1423);
  wire s1424, sub1424, and1424, or1424;
  wire b_inv1424;
  assign b_inv1424 = ~b1424;
  assign s1424  = a1424 ^ b1424 ^ c1424;
  assign sub1424 = a1424 ^ b_inv1424 ^ c1424;
  assign and1424 = a1424 & b1424;
  assign or1424  = a1424 | b1424;
  assign c1425 = (a1424 & b1424) | (a1424 & c1424) | (b1424 & c1424);
  wire c_sub1425;
  assign c_sub1425 = (a1424 & b_inv1424) | (a1424 & c1424) | (b_inv1424 & c1424);
  wire s1425, sub1425, and1425, or1425;
  wire b_inv1425;
  assign b_inv1425 = ~b1425;
  assign s1425  = a1425 ^ b1425 ^ c1425;
  assign sub1425 = a1425 ^ b_inv1425 ^ c1425;
  assign and1425 = a1425 & b1425;
  assign or1425  = a1425 | b1425;
  assign c1426 = (a1425 & b1425) | (a1425 & c1425) | (b1425 & c1425);
  wire c_sub1426;
  assign c_sub1426 = (a1425 & b_inv1425) | (a1425 & c1425) | (b_inv1425 & c1425);
  wire s1426, sub1426, and1426, or1426;
  wire b_inv1426;
  assign b_inv1426 = ~b1426;
  assign s1426  = a1426 ^ b1426 ^ c1426;
  assign sub1426 = a1426 ^ b_inv1426 ^ c1426;
  assign and1426 = a1426 & b1426;
  assign or1426  = a1426 | b1426;
  assign c1427 = (a1426 & b1426) | (a1426 & c1426) | (b1426 & c1426);
  wire c_sub1427;
  assign c_sub1427 = (a1426 & b_inv1426) | (a1426 & c1426) | (b_inv1426 & c1426);
  wire s1427, sub1427, and1427, or1427;
  wire b_inv1427;
  assign b_inv1427 = ~b1427;
  assign s1427  = a1427 ^ b1427 ^ c1427;
  assign sub1427 = a1427 ^ b_inv1427 ^ c1427;
  assign and1427 = a1427 & b1427;
  assign or1427  = a1427 | b1427;
  assign c1428 = (a1427 & b1427) | (a1427 & c1427) | (b1427 & c1427);
  wire c_sub1428;
  assign c_sub1428 = (a1427 & b_inv1427) | (a1427 & c1427) | (b_inv1427 & c1427);
  wire s1428, sub1428, and1428, or1428;
  wire b_inv1428;
  assign b_inv1428 = ~b1428;
  assign s1428  = a1428 ^ b1428 ^ c1428;
  assign sub1428 = a1428 ^ b_inv1428 ^ c1428;
  assign and1428 = a1428 & b1428;
  assign or1428  = a1428 | b1428;
  assign c1429 = (a1428 & b1428) | (a1428 & c1428) | (b1428 & c1428);
  wire c_sub1429;
  assign c_sub1429 = (a1428 & b_inv1428) | (a1428 & c1428) | (b_inv1428 & c1428);
  wire s1429, sub1429, and1429, or1429;
  wire b_inv1429;
  assign b_inv1429 = ~b1429;
  assign s1429  = a1429 ^ b1429 ^ c1429;
  assign sub1429 = a1429 ^ b_inv1429 ^ c1429;
  assign and1429 = a1429 & b1429;
  assign or1429  = a1429 | b1429;
  assign c1430 = (a1429 & b1429) | (a1429 & c1429) | (b1429 & c1429);
  wire c_sub1430;
  assign c_sub1430 = (a1429 & b_inv1429) | (a1429 & c1429) | (b_inv1429 & c1429);
  wire s1430, sub1430, and1430, or1430;
  wire b_inv1430;
  assign b_inv1430 = ~b1430;
  assign s1430  = a1430 ^ b1430 ^ c1430;
  assign sub1430 = a1430 ^ b_inv1430 ^ c1430;
  assign and1430 = a1430 & b1430;
  assign or1430  = a1430 | b1430;
  assign c1431 = (a1430 & b1430) | (a1430 & c1430) | (b1430 & c1430);
  wire c_sub1431;
  assign c_sub1431 = (a1430 & b_inv1430) | (a1430 & c1430) | (b_inv1430 & c1430);
  wire s1431, sub1431, and1431, or1431;
  wire b_inv1431;
  assign b_inv1431 = ~b1431;
  assign s1431  = a1431 ^ b1431 ^ c1431;
  assign sub1431 = a1431 ^ b_inv1431 ^ c1431;
  assign and1431 = a1431 & b1431;
  assign or1431  = a1431 | b1431;
  assign c1432 = (a1431 & b1431) | (a1431 & c1431) | (b1431 & c1431);
  wire c_sub1432;
  assign c_sub1432 = (a1431 & b_inv1431) | (a1431 & c1431) | (b_inv1431 & c1431);
  wire s1432, sub1432, and1432, or1432;
  wire b_inv1432;
  assign b_inv1432 = ~b1432;
  assign s1432  = a1432 ^ b1432 ^ c1432;
  assign sub1432 = a1432 ^ b_inv1432 ^ c1432;
  assign and1432 = a1432 & b1432;
  assign or1432  = a1432 | b1432;
  assign c1433 = (a1432 & b1432) | (a1432 & c1432) | (b1432 & c1432);
  wire c_sub1433;
  assign c_sub1433 = (a1432 & b_inv1432) | (a1432 & c1432) | (b_inv1432 & c1432);
  wire s1433, sub1433, and1433, or1433;
  wire b_inv1433;
  assign b_inv1433 = ~b1433;
  assign s1433  = a1433 ^ b1433 ^ c1433;
  assign sub1433 = a1433 ^ b_inv1433 ^ c1433;
  assign and1433 = a1433 & b1433;
  assign or1433  = a1433 | b1433;
  assign c1434 = (a1433 & b1433) | (a1433 & c1433) | (b1433 & c1433);
  wire c_sub1434;
  assign c_sub1434 = (a1433 & b_inv1433) | (a1433 & c1433) | (b_inv1433 & c1433);
  wire s1434, sub1434, and1434, or1434;
  wire b_inv1434;
  assign b_inv1434 = ~b1434;
  assign s1434  = a1434 ^ b1434 ^ c1434;
  assign sub1434 = a1434 ^ b_inv1434 ^ c1434;
  assign and1434 = a1434 & b1434;
  assign or1434  = a1434 | b1434;
  assign c1435 = (a1434 & b1434) | (a1434 & c1434) | (b1434 & c1434);
  wire c_sub1435;
  assign c_sub1435 = (a1434 & b_inv1434) | (a1434 & c1434) | (b_inv1434 & c1434);
  wire s1435, sub1435, and1435, or1435;
  wire b_inv1435;
  assign b_inv1435 = ~b1435;
  assign s1435  = a1435 ^ b1435 ^ c1435;
  assign sub1435 = a1435 ^ b_inv1435 ^ c1435;
  assign and1435 = a1435 & b1435;
  assign or1435  = a1435 | b1435;
  assign c1436 = (a1435 & b1435) | (a1435 & c1435) | (b1435 & c1435);
  wire c_sub1436;
  assign c_sub1436 = (a1435 & b_inv1435) | (a1435 & c1435) | (b_inv1435 & c1435);
  wire s1436, sub1436, and1436, or1436;
  wire b_inv1436;
  assign b_inv1436 = ~b1436;
  assign s1436  = a1436 ^ b1436 ^ c1436;
  assign sub1436 = a1436 ^ b_inv1436 ^ c1436;
  assign and1436 = a1436 & b1436;
  assign or1436  = a1436 | b1436;
  assign c1437 = (a1436 & b1436) | (a1436 & c1436) | (b1436 & c1436);
  wire c_sub1437;
  assign c_sub1437 = (a1436 & b_inv1436) | (a1436 & c1436) | (b_inv1436 & c1436);
  wire s1437, sub1437, and1437, or1437;
  wire b_inv1437;
  assign b_inv1437 = ~b1437;
  assign s1437  = a1437 ^ b1437 ^ c1437;
  assign sub1437 = a1437 ^ b_inv1437 ^ c1437;
  assign and1437 = a1437 & b1437;
  assign or1437  = a1437 | b1437;
  assign c1438 = (a1437 & b1437) | (a1437 & c1437) | (b1437 & c1437);
  wire c_sub1438;
  assign c_sub1438 = (a1437 & b_inv1437) | (a1437 & c1437) | (b_inv1437 & c1437);
  wire s1438, sub1438, and1438, or1438;
  wire b_inv1438;
  assign b_inv1438 = ~b1438;
  assign s1438  = a1438 ^ b1438 ^ c1438;
  assign sub1438 = a1438 ^ b_inv1438 ^ c1438;
  assign and1438 = a1438 & b1438;
  assign or1438  = a1438 | b1438;
  assign c1439 = (a1438 & b1438) | (a1438 & c1438) | (b1438 & c1438);
  wire c_sub1439;
  assign c_sub1439 = (a1438 & b_inv1438) | (a1438 & c1438) | (b_inv1438 & c1438);
  wire s1439, sub1439, and1439, or1439;
  wire b_inv1439;
  assign b_inv1439 = ~b1439;
  assign s1439  = a1439 ^ b1439 ^ c1439;
  assign sub1439 = a1439 ^ b_inv1439 ^ c1439;
  assign and1439 = a1439 & b1439;
  assign or1439  = a1439 | b1439;
  assign c1440 = (a1439 & b1439) | (a1439 & c1439) | (b1439 & c1439);
  wire c_sub1440;
  assign c_sub1440 = (a1439 & b_inv1439) | (a1439 & c1439) | (b_inv1439 & c1439);
  wire s1440, sub1440, and1440, or1440;
  wire b_inv1440;
  assign b_inv1440 = ~b1440;
  assign s1440  = a1440 ^ b1440 ^ c1440;
  assign sub1440 = a1440 ^ b_inv1440 ^ c1440;
  assign and1440 = a1440 & b1440;
  assign or1440  = a1440 | b1440;
  assign c1441 = (a1440 & b1440) | (a1440 & c1440) | (b1440 & c1440);
  wire c_sub1441;
  assign c_sub1441 = (a1440 & b_inv1440) | (a1440 & c1440) | (b_inv1440 & c1440);
  wire s1441, sub1441, and1441, or1441;
  wire b_inv1441;
  assign b_inv1441 = ~b1441;
  assign s1441  = a1441 ^ b1441 ^ c1441;
  assign sub1441 = a1441 ^ b_inv1441 ^ c1441;
  assign and1441 = a1441 & b1441;
  assign or1441  = a1441 | b1441;
  assign c1442 = (a1441 & b1441) | (a1441 & c1441) | (b1441 & c1441);
  wire c_sub1442;
  assign c_sub1442 = (a1441 & b_inv1441) | (a1441 & c1441) | (b_inv1441 & c1441);
  wire s1442, sub1442, and1442, or1442;
  wire b_inv1442;
  assign b_inv1442 = ~b1442;
  assign s1442  = a1442 ^ b1442 ^ c1442;
  assign sub1442 = a1442 ^ b_inv1442 ^ c1442;
  assign and1442 = a1442 & b1442;
  assign or1442  = a1442 | b1442;
  assign c1443 = (a1442 & b1442) | (a1442 & c1442) | (b1442 & c1442);
  wire c_sub1443;
  assign c_sub1443 = (a1442 & b_inv1442) | (a1442 & c1442) | (b_inv1442 & c1442);
  wire s1443, sub1443, and1443, or1443;
  wire b_inv1443;
  assign b_inv1443 = ~b1443;
  assign s1443  = a1443 ^ b1443 ^ c1443;
  assign sub1443 = a1443 ^ b_inv1443 ^ c1443;
  assign and1443 = a1443 & b1443;
  assign or1443  = a1443 | b1443;
  assign c1444 = (a1443 & b1443) | (a1443 & c1443) | (b1443 & c1443);
  wire c_sub1444;
  assign c_sub1444 = (a1443 & b_inv1443) | (a1443 & c1443) | (b_inv1443 & c1443);
  wire s1444, sub1444, and1444, or1444;
  wire b_inv1444;
  assign b_inv1444 = ~b1444;
  assign s1444  = a1444 ^ b1444 ^ c1444;
  assign sub1444 = a1444 ^ b_inv1444 ^ c1444;
  assign and1444 = a1444 & b1444;
  assign or1444  = a1444 | b1444;
  assign c1445 = (a1444 & b1444) | (a1444 & c1444) | (b1444 & c1444);
  wire c_sub1445;
  assign c_sub1445 = (a1444 & b_inv1444) | (a1444 & c1444) | (b_inv1444 & c1444);
  wire s1445, sub1445, and1445, or1445;
  wire b_inv1445;
  assign b_inv1445 = ~b1445;
  assign s1445  = a1445 ^ b1445 ^ c1445;
  assign sub1445 = a1445 ^ b_inv1445 ^ c1445;
  assign and1445 = a1445 & b1445;
  assign or1445  = a1445 | b1445;
  assign c1446 = (a1445 & b1445) | (a1445 & c1445) | (b1445 & c1445);
  wire c_sub1446;
  assign c_sub1446 = (a1445 & b_inv1445) | (a1445 & c1445) | (b_inv1445 & c1445);
  wire s1446, sub1446, and1446, or1446;
  wire b_inv1446;
  assign b_inv1446 = ~b1446;
  assign s1446  = a1446 ^ b1446 ^ c1446;
  assign sub1446 = a1446 ^ b_inv1446 ^ c1446;
  assign and1446 = a1446 & b1446;
  assign or1446  = a1446 | b1446;
  assign c1447 = (a1446 & b1446) | (a1446 & c1446) | (b1446 & c1446);
  wire c_sub1447;
  assign c_sub1447 = (a1446 & b_inv1446) | (a1446 & c1446) | (b_inv1446 & c1446);
  wire s1447, sub1447, and1447, or1447;
  wire b_inv1447;
  assign b_inv1447 = ~b1447;
  assign s1447  = a1447 ^ b1447 ^ c1447;
  assign sub1447 = a1447 ^ b_inv1447 ^ c1447;
  assign and1447 = a1447 & b1447;
  assign or1447  = a1447 | b1447;
  assign c1448 = (a1447 & b1447) | (a1447 & c1447) | (b1447 & c1447);
  wire c_sub1448;
  assign c_sub1448 = (a1447 & b_inv1447) | (a1447 & c1447) | (b_inv1447 & c1447);
  wire s1448, sub1448, and1448, or1448;
  wire b_inv1448;
  assign b_inv1448 = ~b1448;
  assign s1448  = a1448 ^ b1448 ^ c1448;
  assign sub1448 = a1448 ^ b_inv1448 ^ c1448;
  assign and1448 = a1448 & b1448;
  assign or1448  = a1448 | b1448;
  assign c1449 = (a1448 & b1448) | (a1448 & c1448) | (b1448 & c1448);
  wire c_sub1449;
  assign c_sub1449 = (a1448 & b_inv1448) | (a1448 & c1448) | (b_inv1448 & c1448);
  wire s1449, sub1449, and1449, or1449;
  wire b_inv1449;
  assign b_inv1449 = ~b1449;
  assign s1449  = a1449 ^ b1449 ^ c1449;
  assign sub1449 = a1449 ^ b_inv1449 ^ c1449;
  assign and1449 = a1449 & b1449;
  assign or1449  = a1449 | b1449;
  assign c1450 = (a1449 & b1449) | (a1449 & c1449) | (b1449 & c1449);
  wire c_sub1450;
  assign c_sub1450 = (a1449 & b_inv1449) | (a1449 & c1449) | (b_inv1449 & c1449);
  wire s1450, sub1450, and1450, or1450;
  wire b_inv1450;
  assign b_inv1450 = ~b1450;
  assign s1450  = a1450 ^ b1450 ^ c1450;
  assign sub1450 = a1450 ^ b_inv1450 ^ c1450;
  assign and1450 = a1450 & b1450;
  assign or1450  = a1450 | b1450;
  assign c1451 = (a1450 & b1450) | (a1450 & c1450) | (b1450 & c1450);
  wire c_sub1451;
  assign c_sub1451 = (a1450 & b_inv1450) | (a1450 & c1450) | (b_inv1450 & c1450);
  wire s1451, sub1451, and1451, or1451;
  wire b_inv1451;
  assign b_inv1451 = ~b1451;
  assign s1451  = a1451 ^ b1451 ^ c1451;
  assign sub1451 = a1451 ^ b_inv1451 ^ c1451;
  assign and1451 = a1451 & b1451;
  assign or1451  = a1451 | b1451;
  assign c1452 = (a1451 & b1451) | (a1451 & c1451) | (b1451 & c1451);
  wire c_sub1452;
  assign c_sub1452 = (a1451 & b_inv1451) | (a1451 & c1451) | (b_inv1451 & c1451);
  wire s1452, sub1452, and1452, or1452;
  wire b_inv1452;
  assign b_inv1452 = ~b1452;
  assign s1452  = a1452 ^ b1452 ^ c1452;
  assign sub1452 = a1452 ^ b_inv1452 ^ c1452;
  assign and1452 = a1452 & b1452;
  assign or1452  = a1452 | b1452;
  assign c1453 = (a1452 & b1452) | (a1452 & c1452) | (b1452 & c1452);
  wire c_sub1453;
  assign c_sub1453 = (a1452 & b_inv1452) | (a1452 & c1452) | (b_inv1452 & c1452);
  wire s1453, sub1453, and1453, or1453;
  wire b_inv1453;
  assign b_inv1453 = ~b1453;
  assign s1453  = a1453 ^ b1453 ^ c1453;
  assign sub1453 = a1453 ^ b_inv1453 ^ c1453;
  assign and1453 = a1453 & b1453;
  assign or1453  = a1453 | b1453;
  assign c1454 = (a1453 & b1453) | (a1453 & c1453) | (b1453 & c1453);
  wire c_sub1454;
  assign c_sub1454 = (a1453 & b_inv1453) | (a1453 & c1453) | (b_inv1453 & c1453);
  wire s1454, sub1454, and1454, or1454;
  wire b_inv1454;
  assign b_inv1454 = ~b1454;
  assign s1454  = a1454 ^ b1454 ^ c1454;
  assign sub1454 = a1454 ^ b_inv1454 ^ c1454;
  assign and1454 = a1454 & b1454;
  assign or1454  = a1454 | b1454;
  assign c1455 = (a1454 & b1454) | (a1454 & c1454) | (b1454 & c1454);
  wire c_sub1455;
  assign c_sub1455 = (a1454 & b_inv1454) | (a1454 & c1454) | (b_inv1454 & c1454);
  wire s1455, sub1455, and1455, or1455;
  wire b_inv1455;
  assign b_inv1455 = ~b1455;
  assign s1455  = a1455 ^ b1455 ^ c1455;
  assign sub1455 = a1455 ^ b_inv1455 ^ c1455;
  assign and1455 = a1455 & b1455;
  assign or1455  = a1455 | b1455;
  assign c1456 = (a1455 & b1455) | (a1455 & c1455) | (b1455 & c1455);
  wire c_sub1456;
  assign c_sub1456 = (a1455 & b_inv1455) | (a1455 & c1455) | (b_inv1455 & c1455);
  wire s1456, sub1456, and1456, or1456;
  wire b_inv1456;
  assign b_inv1456 = ~b1456;
  assign s1456  = a1456 ^ b1456 ^ c1456;
  assign sub1456 = a1456 ^ b_inv1456 ^ c1456;
  assign and1456 = a1456 & b1456;
  assign or1456  = a1456 | b1456;
  assign c1457 = (a1456 & b1456) | (a1456 & c1456) | (b1456 & c1456);
  wire c_sub1457;
  assign c_sub1457 = (a1456 & b_inv1456) | (a1456 & c1456) | (b_inv1456 & c1456);
  wire s1457, sub1457, and1457, or1457;
  wire b_inv1457;
  assign b_inv1457 = ~b1457;
  assign s1457  = a1457 ^ b1457 ^ c1457;
  assign sub1457 = a1457 ^ b_inv1457 ^ c1457;
  assign and1457 = a1457 & b1457;
  assign or1457  = a1457 | b1457;
  assign c1458 = (a1457 & b1457) | (a1457 & c1457) | (b1457 & c1457);
  wire c_sub1458;
  assign c_sub1458 = (a1457 & b_inv1457) | (a1457 & c1457) | (b_inv1457 & c1457);
  wire s1458, sub1458, and1458, or1458;
  wire b_inv1458;
  assign b_inv1458 = ~b1458;
  assign s1458  = a1458 ^ b1458 ^ c1458;
  assign sub1458 = a1458 ^ b_inv1458 ^ c1458;
  assign and1458 = a1458 & b1458;
  assign or1458  = a1458 | b1458;
  assign c1459 = (a1458 & b1458) | (a1458 & c1458) | (b1458 & c1458);
  wire c_sub1459;
  assign c_sub1459 = (a1458 & b_inv1458) | (a1458 & c1458) | (b_inv1458 & c1458);
  wire s1459, sub1459, and1459, or1459;
  wire b_inv1459;
  assign b_inv1459 = ~b1459;
  assign s1459  = a1459 ^ b1459 ^ c1459;
  assign sub1459 = a1459 ^ b_inv1459 ^ c1459;
  assign and1459 = a1459 & b1459;
  assign or1459  = a1459 | b1459;
  assign c1460 = (a1459 & b1459) | (a1459 & c1459) | (b1459 & c1459);
  wire c_sub1460;
  assign c_sub1460 = (a1459 & b_inv1459) | (a1459 & c1459) | (b_inv1459 & c1459);
  wire s1460, sub1460, and1460, or1460;
  wire b_inv1460;
  assign b_inv1460 = ~b1460;
  assign s1460  = a1460 ^ b1460 ^ c1460;
  assign sub1460 = a1460 ^ b_inv1460 ^ c1460;
  assign and1460 = a1460 & b1460;
  assign or1460  = a1460 | b1460;
  assign c1461 = (a1460 & b1460) | (a1460 & c1460) | (b1460 & c1460);
  wire c_sub1461;
  assign c_sub1461 = (a1460 & b_inv1460) | (a1460 & c1460) | (b_inv1460 & c1460);
  wire s1461, sub1461, and1461, or1461;
  wire b_inv1461;
  assign b_inv1461 = ~b1461;
  assign s1461  = a1461 ^ b1461 ^ c1461;
  assign sub1461 = a1461 ^ b_inv1461 ^ c1461;
  assign and1461 = a1461 & b1461;
  assign or1461  = a1461 | b1461;
  assign c1462 = (a1461 & b1461) | (a1461 & c1461) | (b1461 & c1461);
  wire c_sub1462;
  assign c_sub1462 = (a1461 & b_inv1461) | (a1461 & c1461) | (b_inv1461 & c1461);
  wire s1462, sub1462, and1462, or1462;
  wire b_inv1462;
  assign b_inv1462 = ~b1462;
  assign s1462  = a1462 ^ b1462 ^ c1462;
  assign sub1462 = a1462 ^ b_inv1462 ^ c1462;
  assign and1462 = a1462 & b1462;
  assign or1462  = a1462 | b1462;
  assign c1463 = (a1462 & b1462) | (a1462 & c1462) | (b1462 & c1462);
  wire c_sub1463;
  assign c_sub1463 = (a1462 & b_inv1462) | (a1462 & c1462) | (b_inv1462 & c1462);
  wire s1463, sub1463, and1463, or1463;
  wire b_inv1463;
  assign b_inv1463 = ~b1463;
  assign s1463  = a1463 ^ b1463 ^ c1463;
  assign sub1463 = a1463 ^ b_inv1463 ^ c1463;
  assign and1463 = a1463 & b1463;
  assign or1463  = a1463 | b1463;
  assign c1464 = (a1463 & b1463) | (a1463 & c1463) | (b1463 & c1463);
  wire c_sub1464;
  assign c_sub1464 = (a1463 & b_inv1463) | (a1463 & c1463) | (b_inv1463 & c1463);
  wire s1464, sub1464, and1464, or1464;
  wire b_inv1464;
  assign b_inv1464 = ~b1464;
  assign s1464  = a1464 ^ b1464 ^ c1464;
  assign sub1464 = a1464 ^ b_inv1464 ^ c1464;
  assign and1464 = a1464 & b1464;
  assign or1464  = a1464 | b1464;
  assign c1465 = (a1464 & b1464) | (a1464 & c1464) | (b1464 & c1464);
  wire c_sub1465;
  assign c_sub1465 = (a1464 & b_inv1464) | (a1464 & c1464) | (b_inv1464 & c1464);
  wire s1465, sub1465, and1465, or1465;
  wire b_inv1465;
  assign b_inv1465 = ~b1465;
  assign s1465  = a1465 ^ b1465 ^ c1465;
  assign sub1465 = a1465 ^ b_inv1465 ^ c1465;
  assign and1465 = a1465 & b1465;
  assign or1465  = a1465 | b1465;
  assign c1466 = (a1465 & b1465) | (a1465 & c1465) | (b1465 & c1465);
  wire c_sub1466;
  assign c_sub1466 = (a1465 & b_inv1465) | (a1465 & c1465) | (b_inv1465 & c1465);
  wire s1466, sub1466, and1466, or1466;
  wire b_inv1466;
  assign b_inv1466 = ~b1466;
  assign s1466  = a1466 ^ b1466 ^ c1466;
  assign sub1466 = a1466 ^ b_inv1466 ^ c1466;
  assign and1466 = a1466 & b1466;
  assign or1466  = a1466 | b1466;
  assign c1467 = (a1466 & b1466) | (a1466 & c1466) | (b1466 & c1466);
  wire c_sub1467;
  assign c_sub1467 = (a1466 & b_inv1466) | (a1466 & c1466) | (b_inv1466 & c1466);
  wire s1467, sub1467, and1467, or1467;
  wire b_inv1467;
  assign b_inv1467 = ~b1467;
  assign s1467  = a1467 ^ b1467 ^ c1467;
  assign sub1467 = a1467 ^ b_inv1467 ^ c1467;
  assign and1467 = a1467 & b1467;
  assign or1467  = a1467 | b1467;
  assign c1468 = (a1467 & b1467) | (a1467 & c1467) | (b1467 & c1467);
  wire c_sub1468;
  assign c_sub1468 = (a1467 & b_inv1467) | (a1467 & c1467) | (b_inv1467 & c1467);
  wire s1468, sub1468, and1468, or1468;
  wire b_inv1468;
  assign b_inv1468 = ~b1468;
  assign s1468  = a1468 ^ b1468 ^ c1468;
  assign sub1468 = a1468 ^ b_inv1468 ^ c1468;
  assign and1468 = a1468 & b1468;
  assign or1468  = a1468 | b1468;
  assign c1469 = (a1468 & b1468) | (a1468 & c1468) | (b1468 & c1468);
  wire c_sub1469;
  assign c_sub1469 = (a1468 & b_inv1468) | (a1468 & c1468) | (b_inv1468 & c1468);
  wire s1469, sub1469, and1469, or1469;
  wire b_inv1469;
  assign b_inv1469 = ~b1469;
  assign s1469  = a1469 ^ b1469 ^ c1469;
  assign sub1469 = a1469 ^ b_inv1469 ^ c1469;
  assign and1469 = a1469 & b1469;
  assign or1469  = a1469 | b1469;
  assign c1470 = (a1469 & b1469) | (a1469 & c1469) | (b1469 & c1469);
  wire c_sub1470;
  assign c_sub1470 = (a1469 & b_inv1469) | (a1469 & c1469) | (b_inv1469 & c1469);
  wire s1470, sub1470, and1470, or1470;
  wire b_inv1470;
  assign b_inv1470 = ~b1470;
  assign s1470  = a1470 ^ b1470 ^ c1470;
  assign sub1470 = a1470 ^ b_inv1470 ^ c1470;
  assign and1470 = a1470 & b1470;
  assign or1470  = a1470 | b1470;
  assign c1471 = (a1470 & b1470) | (a1470 & c1470) | (b1470 & c1470);
  wire c_sub1471;
  assign c_sub1471 = (a1470 & b_inv1470) | (a1470 & c1470) | (b_inv1470 & c1470);
  wire s1471, sub1471, and1471, or1471;
  wire b_inv1471;
  assign b_inv1471 = ~b1471;
  assign s1471  = a1471 ^ b1471 ^ c1471;
  assign sub1471 = a1471 ^ b_inv1471 ^ c1471;
  assign and1471 = a1471 & b1471;
  assign or1471  = a1471 | b1471;
  assign c1472 = (a1471 & b1471) | (a1471 & c1471) | (b1471 & c1471);
  wire c_sub1472;
  assign c_sub1472 = (a1471 & b_inv1471) | (a1471 & c1471) | (b_inv1471 & c1471);
  wire s1472, sub1472, and1472, or1472;
  wire b_inv1472;
  assign b_inv1472 = ~b1472;
  assign s1472  = a1472 ^ b1472 ^ c1472;
  assign sub1472 = a1472 ^ b_inv1472 ^ c1472;
  assign and1472 = a1472 & b1472;
  assign or1472  = a1472 | b1472;
  assign c1473 = (a1472 & b1472) | (a1472 & c1472) | (b1472 & c1472);
  wire c_sub1473;
  assign c_sub1473 = (a1472 & b_inv1472) | (a1472 & c1472) | (b_inv1472 & c1472);
  wire s1473, sub1473, and1473, or1473;
  wire b_inv1473;
  assign b_inv1473 = ~b1473;
  assign s1473  = a1473 ^ b1473 ^ c1473;
  assign sub1473 = a1473 ^ b_inv1473 ^ c1473;
  assign and1473 = a1473 & b1473;
  assign or1473  = a1473 | b1473;
  assign c1474 = (a1473 & b1473) | (a1473 & c1473) | (b1473 & c1473);
  wire c_sub1474;
  assign c_sub1474 = (a1473 & b_inv1473) | (a1473 & c1473) | (b_inv1473 & c1473);
  wire s1474, sub1474, and1474, or1474;
  wire b_inv1474;
  assign b_inv1474 = ~b1474;
  assign s1474  = a1474 ^ b1474 ^ c1474;
  assign sub1474 = a1474 ^ b_inv1474 ^ c1474;
  assign and1474 = a1474 & b1474;
  assign or1474  = a1474 | b1474;
  assign c1475 = (a1474 & b1474) | (a1474 & c1474) | (b1474 & c1474);
  wire c_sub1475;
  assign c_sub1475 = (a1474 & b_inv1474) | (a1474 & c1474) | (b_inv1474 & c1474);
  wire s1475, sub1475, and1475, or1475;
  wire b_inv1475;
  assign b_inv1475 = ~b1475;
  assign s1475  = a1475 ^ b1475 ^ c1475;
  assign sub1475 = a1475 ^ b_inv1475 ^ c1475;
  assign and1475 = a1475 & b1475;
  assign or1475  = a1475 | b1475;
  assign c1476 = (a1475 & b1475) | (a1475 & c1475) | (b1475 & c1475);
  wire c_sub1476;
  assign c_sub1476 = (a1475 & b_inv1475) | (a1475 & c1475) | (b_inv1475 & c1475);
  wire s1476, sub1476, and1476, or1476;
  wire b_inv1476;
  assign b_inv1476 = ~b1476;
  assign s1476  = a1476 ^ b1476 ^ c1476;
  assign sub1476 = a1476 ^ b_inv1476 ^ c1476;
  assign and1476 = a1476 & b1476;
  assign or1476  = a1476 | b1476;
  assign c1477 = (a1476 & b1476) | (a1476 & c1476) | (b1476 & c1476);
  wire c_sub1477;
  assign c_sub1477 = (a1476 & b_inv1476) | (a1476 & c1476) | (b_inv1476 & c1476);
  wire s1477, sub1477, and1477, or1477;
  wire b_inv1477;
  assign b_inv1477 = ~b1477;
  assign s1477  = a1477 ^ b1477 ^ c1477;
  assign sub1477 = a1477 ^ b_inv1477 ^ c1477;
  assign and1477 = a1477 & b1477;
  assign or1477  = a1477 | b1477;
  assign c1478 = (a1477 & b1477) | (a1477 & c1477) | (b1477 & c1477);
  wire c_sub1478;
  assign c_sub1478 = (a1477 & b_inv1477) | (a1477 & c1477) | (b_inv1477 & c1477);
  wire s1478, sub1478, and1478, or1478;
  wire b_inv1478;
  assign b_inv1478 = ~b1478;
  assign s1478  = a1478 ^ b1478 ^ c1478;
  assign sub1478 = a1478 ^ b_inv1478 ^ c1478;
  assign and1478 = a1478 & b1478;
  assign or1478  = a1478 | b1478;
  assign c1479 = (a1478 & b1478) | (a1478 & c1478) | (b1478 & c1478);
  wire c_sub1479;
  assign c_sub1479 = (a1478 & b_inv1478) | (a1478 & c1478) | (b_inv1478 & c1478);
  wire s1479, sub1479, and1479, or1479;
  wire b_inv1479;
  assign b_inv1479 = ~b1479;
  assign s1479  = a1479 ^ b1479 ^ c1479;
  assign sub1479 = a1479 ^ b_inv1479 ^ c1479;
  assign and1479 = a1479 & b1479;
  assign or1479  = a1479 | b1479;
  assign c1480 = (a1479 & b1479) | (a1479 & c1479) | (b1479 & c1479);
  wire c_sub1480;
  assign c_sub1480 = (a1479 & b_inv1479) | (a1479 & c1479) | (b_inv1479 & c1479);
  wire s1480, sub1480, and1480, or1480;
  wire b_inv1480;
  assign b_inv1480 = ~b1480;
  assign s1480  = a1480 ^ b1480 ^ c1480;
  assign sub1480 = a1480 ^ b_inv1480 ^ c1480;
  assign and1480 = a1480 & b1480;
  assign or1480  = a1480 | b1480;
  assign c1481 = (a1480 & b1480) | (a1480 & c1480) | (b1480 & c1480);
  wire c_sub1481;
  assign c_sub1481 = (a1480 & b_inv1480) | (a1480 & c1480) | (b_inv1480 & c1480);
  wire s1481, sub1481, and1481, or1481;
  wire b_inv1481;
  assign b_inv1481 = ~b1481;
  assign s1481  = a1481 ^ b1481 ^ c1481;
  assign sub1481 = a1481 ^ b_inv1481 ^ c1481;
  assign and1481 = a1481 & b1481;
  assign or1481  = a1481 | b1481;
  assign c1482 = (a1481 & b1481) | (a1481 & c1481) | (b1481 & c1481);
  wire c_sub1482;
  assign c_sub1482 = (a1481 & b_inv1481) | (a1481 & c1481) | (b_inv1481 & c1481);
  wire s1482, sub1482, and1482, or1482;
  wire b_inv1482;
  assign b_inv1482 = ~b1482;
  assign s1482  = a1482 ^ b1482 ^ c1482;
  assign sub1482 = a1482 ^ b_inv1482 ^ c1482;
  assign and1482 = a1482 & b1482;
  assign or1482  = a1482 | b1482;
  assign c1483 = (a1482 & b1482) | (a1482 & c1482) | (b1482 & c1482);
  wire c_sub1483;
  assign c_sub1483 = (a1482 & b_inv1482) | (a1482 & c1482) | (b_inv1482 & c1482);
  wire s1483, sub1483, and1483, or1483;
  wire b_inv1483;
  assign b_inv1483 = ~b1483;
  assign s1483  = a1483 ^ b1483 ^ c1483;
  assign sub1483 = a1483 ^ b_inv1483 ^ c1483;
  assign and1483 = a1483 & b1483;
  assign or1483  = a1483 | b1483;
  assign c1484 = (a1483 & b1483) | (a1483 & c1483) | (b1483 & c1483);
  wire c_sub1484;
  assign c_sub1484 = (a1483 & b_inv1483) | (a1483 & c1483) | (b_inv1483 & c1483);
  wire s1484, sub1484, and1484, or1484;
  wire b_inv1484;
  assign b_inv1484 = ~b1484;
  assign s1484  = a1484 ^ b1484 ^ c1484;
  assign sub1484 = a1484 ^ b_inv1484 ^ c1484;
  assign and1484 = a1484 & b1484;
  assign or1484  = a1484 | b1484;
  assign c1485 = (a1484 & b1484) | (a1484 & c1484) | (b1484 & c1484);
  wire c_sub1485;
  assign c_sub1485 = (a1484 & b_inv1484) | (a1484 & c1484) | (b_inv1484 & c1484);
  wire s1485, sub1485, and1485, or1485;
  wire b_inv1485;
  assign b_inv1485 = ~b1485;
  assign s1485  = a1485 ^ b1485 ^ c1485;
  assign sub1485 = a1485 ^ b_inv1485 ^ c1485;
  assign and1485 = a1485 & b1485;
  assign or1485  = a1485 | b1485;
  assign c1486 = (a1485 & b1485) | (a1485 & c1485) | (b1485 & c1485);
  wire c_sub1486;
  assign c_sub1486 = (a1485 & b_inv1485) | (a1485 & c1485) | (b_inv1485 & c1485);
  wire s1486, sub1486, and1486, or1486;
  wire b_inv1486;
  assign b_inv1486 = ~b1486;
  assign s1486  = a1486 ^ b1486 ^ c1486;
  assign sub1486 = a1486 ^ b_inv1486 ^ c1486;
  assign and1486 = a1486 & b1486;
  assign or1486  = a1486 | b1486;
  assign c1487 = (a1486 & b1486) | (a1486 & c1486) | (b1486 & c1486);
  wire c_sub1487;
  assign c_sub1487 = (a1486 & b_inv1486) | (a1486 & c1486) | (b_inv1486 & c1486);
  wire s1487, sub1487, and1487, or1487;
  wire b_inv1487;
  assign b_inv1487 = ~b1487;
  assign s1487  = a1487 ^ b1487 ^ c1487;
  assign sub1487 = a1487 ^ b_inv1487 ^ c1487;
  assign and1487 = a1487 & b1487;
  assign or1487  = a1487 | b1487;
  assign c1488 = (a1487 & b1487) | (a1487 & c1487) | (b1487 & c1487);
  wire c_sub1488;
  assign c_sub1488 = (a1487 & b_inv1487) | (a1487 & c1487) | (b_inv1487 & c1487);
  wire s1488, sub1488, and1488, or1488;
  wire b_inv1488;
  assign b_inv1488 = ~b1488;
  assign s1488  = a1488 ^ b1488 ^ c1488;
  assign sub1488 = a1488 ^ b_inv1488 ^ c1488;
  assign and1488 = a1488 & b1488;
  assign or1488  = a1488 | b1488;
  assign c1489 = (a1488 & b1488) | (a1488 & c1488) | (b1488 & c1488);
  wire c_sub1489;
  assign c_sub1489 = (a1488 & b_inv1488) | (a1488 & c1488) | (b_inv1488 & c1488);
  wire s1489, sub1489, and1489, or1489;
  wire b_inv1489;
  assign b_inv1489 = ~b1489;
  assign s1489  = a1489 ^ b1489 ^ c1489;
  assign sub1489 = a1489 ^ b_inv1489 ^ c1489;
  assign and1489 = a1489 & b1489;
  assign or1489  = a1489 | b1489;
  assign c1490 = (a1489 & b1489) | (a1489 & c1489) | (b1489 & c1489);
  wire c_sub1490;
  assign c_sub1490 = (a1489 & b_inv1489) | (a1489 & c1489) | (b_inv1489 & c1489);
  wire s1490, sub1490, and1490, or1490;
  wire b_inv1490;
  assign b_inv1490 = ~b1490;
  assign s1490  = a1490 ^ b1490 ^ c1490;
  assign sub1490 = a1490 ^ b_inv1490 ^ c1490;
  assign and1490 = a1490 & b1490;
  assign or1490  = a1490 | b1490;
  assign c1491 = (a1490 & b1490) | (a1490 & c1490) | (b1490 & c1490);
  wire c_sub1491;
  assign c_sub1491 = (a1490 & b_inv1490) | (a1490 & c1490) | (b_inv1490 & c1490);
  wire s1491, sub1491, and1491, or1491;
  wire b_inv1491;
  assign b_inv1491 = ~b1491;
  assign s1491  = a1491 ^ b1491 ^ c1491;
  assign sub1491 = a1491 ^ b_inv1491 ^ c1491;
  assign and1491 = a1491 & b1491;
  assign or1491  = a1491 | b1491;
  assign c1492 = (a1491 & b1491) | (a1491 & c1491) | (b1491 & c1491);
  wire c_sub1492;
  assign c_sub1492 = (a1491 & b_inv1491) | (a1491 & c1491) | (b_inv1491 & c1491);
  wire s1492, sub1492, and1492, or1492;
  wire b_inv1492;
  assign b_inv1492 = ~b1492;
  assign s1492  = a1492 ^ b1492 ^ c1492;
  assign sub1492 = a1492 ^ b_inv1492 ^ c1492;
  assign and1492 = a1492 & b1492;
  assign or1492  = a1492 | b1492;
  assign c1493 = (a1492 & b1492) | (a1492 & c1492) | (b1492 & c1492);
  wire c_sub1493;
  assign c_sub1493 = (a1492 & b_inv1492) | (a1492 & c1492) | (b_inv1492 & c1492);
  wire s1493, sub1493, and1493, or1493;
  wire b_inv1493;
  assign b_inv1493 = ~b1493;
  assign s1493  = a1493 ^ b1493 ^ c1493;
  assign sub1493 = a1493 ^ b_inv1493 ^ c1493;
  assign and1493 = a1493 & b1493;
  assign or1493  = a1493 | b1493;
  assign c1494 = (a1493 & b1493) | (a1493 & c1493) | (b1493 & c1493);
  wire c_sub1494;
  assign c_sub1494 = (a1493 & b_inv1493) | (a1493 & c1493) | (b_inv1493 & c1493);
  wire s1494, sub1494, and1494, or1494;
  wire b_inv1494;
  assign b_inv1494 = ~b1494;
  assign s1494  = a1494 ^ b1494 ^ c1494;
  assign sub1494 = a1494 ^ b_inv1494 ^ c1494;
  assign and1494 = a1494 & b1494;
  assign or1494  = a1494 | b1494;
  assign c1495 = (a1494 & b1494) | (a1494 & c1494) | (b1494 & c1494);
  wire c_sub1495;
  assign c_sub1495 = (a1494 & b_inv1494) | (a1494 & c1494) | (b_inv1494 & c1494);
  wire s1495, sub1495, and1495, or1495;
  wire b_inv1495;
  assign b_inv1495 = ~b1495;
  assign s1495  = a1495 ^ b1495 ^ c1495;
  assign sub1495 = a1495 ^ b_inv1495 ^ c1495;
  assign and1495 = a1495 & b1495;
  assign or1495  = a1495 | b1495;
  assign c1496 = (a1495 & b1495) | (a1495 & c1495) | (b1495 & c1495);
  wire c_sub1496;
  assign c_sub1496 = (a1495 & b_inv1495) | (a1495 & c1495) | (b_inv1495 & c1495);
  wire s1496, sub1496, and1496, or1496;
  wire b_inv1496;
  assign b_inv1496 = ~b1496;
  assign s1496  = a1496 ^ b1496 ^ c1496;
  assign sub1496 = a1496 ^ b_inv1496 ^ c1496;
  assign and1496 = a1496 & b1496;
  assign or1496  = a1496 | b1496;
  assign c1497 = (a1496 & b1496) | (a1496 & c1496) | (b1496 & c1496);
  wire c_sub1497;
  assign c_sub1497 = (a1496 & b_inv1496) | (a1496 & c1496) | (b_inv1496 & c1496);
  wire s1497, sub1497, and1497, or1497;
  wire b_inv1497;
  assign b_inv1497 = ~b1497;
  assign s1497  = a1497 ^ b1497 ^ c1497;
  assign sub1497 = a1497 ^ b_inv1497 ^ c1497;
  assign and1497 = a1497 & b1497;
  assign or1497  = a1497 | b1497;
  assign c1498 = (a1497 & b1497) | (a1497 & c1497) | (b1497 & c1497);
  wire c_sub1498;
  assign c_sub1498 = (a1497 & b_inv1497) | (a1497 & c1497) | (b_inv1497 & c1497);
  wire s1498, sub1498, and1498, or1498;
  wire b_inv1498;
  assign b_inv1498 = ~b1498;
  assign s1498  = a1498 ^ b1498 ^ c1498;
  assign sub1498 = a1498 ^ b_inv1498 ^ c1498;
  assign and1498 = a1498 & b1498;
  assign or1498  = a1498 | b1498;
  assign c1499 = (a1498 & b1498) | (a1498 & c1498) | (b1498 & c1498);
  wire c_sub1499;
  assign c_sub1499 = (a1498 & b_inv1498) | (a1498 & c1498) | (b_inv1498 & c1498);
  wire s1499, sub1499, and1499, or1499;
  wire b_inv1499;
  assign b_inv1499 = ~b1499;
  assign s1499  = a1499 ^ b1499 ^ c1499;
  assign sub1499 = a1499 ^ b_inv1499 ^ c1499;
  assign and1499 = a1499 & b1499;
  assign or1499  = a1499 | b1499;
  assign c1500 = (a1499 & b1499) | (a1499 & c1499) | (b1499 & c1499);
  wire c_sub1500;
  assign c_sub1500 = (a1499 & b_inv1499) | (a1499 & c1499) | (b_inv1499 & c1499);
  wire s1500, sub1500, and1500, or1500;
  wire b_inv1500;
  assign b_inv1500 = ~b1500;
  assign s1500  = a1500 ^ b1500 ^ c1500;
  assign sub1500 = a1500 ^ b_inv1500 ^ c1500;
  assign and1500 = a1500 & b1500;
  assign or1500  = a1500 | b1500;
  assign c1501 = (a1500 & b1500) | (a1500 & c1500) | (b1500 & c1500);
  wire c_sub1501;
  assign c_sub1501 = (a1500 & b_inv1500) | (a1500 & c1500) | (b_inv1500 & c1500);
  wire s1501, sub1501, and1501, or1501;
  wire b_inv1501;
  assign b_inv1501 = ~b1501;
  assign s1501  = a1501 ^ b1501 ^ c1501;
  assign sub1501 = a1501 ^ b_inv1501 ^ c1501;
  assign and1501 = a1501 & b1501;
  assign or1501  = a1501 | b1501;
  assign c1502 = (a1501 & b1501) | (a1501 & c1501) | (b1501 & c1501);
  wire c_sub1502;
  assign c_sub1502 = (a1501 & b_inv1501) | (a1501 & c1501) | (b_inv1501 & c1501);
  wire s1502, sub1502, and1502, or1502;
  wire b_inv1502;
  assign b_inv1502 = ~b1502;
  assign s1502  = a1502 ^ b1502 ^ c1502;
  assign sub1502 = a1502 ^ b_inv1502 ^ c1502;
  assign and1502 = a1502 & b1502;
  assign or1502  = a1502 | b1502;
  assign c1503 = (a1502 & b1502) | (a1502 & c1502) | (b1502 & c1502);
  wire c_sub1503;
  assign c_sub1503 = (a1502 & b_inv1502) | (a1502 & c1502) | (b_inv1502 & c1502);
  wire s1503, sub1503, and1503, or1503;
  wire b_inv1503;
  assign b_inv1503 = ~b1503;
  assign s1503  = a1503 ^ b1503 ^ c1503;
  assign sub1503 = a1503 ^ b_inv1503 ^ c1503;
  assign and1503 = a1503 & b1503;
  assign or1503  = a1503 | b1503;
  assign c1504 = (a1503 & b1503) | (a1503 & c1503) | (b1503 & c1503);
  wire c_sub1504;
  assign c_sub1504 = (a1503 & b_inv1503) | (a1503 & c1503) | (b_inv1503 & c1503);
  wire s1504, sub1504, and1504, or1504;
  wire b_inv1504;
  assign b_inv1504 = ~b1504;
  assign s1504  = a1504 ^ b1504 ^ c1504;
  assign sub1504 = a1504 ^ b_inv1504 ^ c1504;
  assign and1504 = a1504 & b1504;
  assign or1504  = a1504 | b1504;
  assign c1505 = (a1504 & b1504) | (a1504 & c1504) | (b1504 & c1504);
  wire c_sub1505;
  assign c_sub1505 = (a1504 & b_inv1504) | (a1504 & c1504) | (b_inv1504 & c1504);
  wire s1505, sub1505, and1505, or1505;
  wire b_inv1505;
  assign b_inv1505 = ~b1505;
  assign s1505  = a1505 ^ b1505 ^ c1505;
  assign sub1505 = a1505 ^ b_inv1505 ^ c1505;
  assign and1505 = a1505 & b1505;
  assign or1505  = a1505 | b1505;
  assign c1506 = (a1505 & b1505) | (a1505 & c1505) | (b1505 & c1505);
  wire c_sub1506;
  assign c_sub1506 = (a1505 & b_inv1505) | (a1505 & c1505) | (b_inv1505 & c1505);
  wire s1506, sub1506, and1506, or1506;
  wire b_inv1506;
  assign b_inv1506 = ~b1506;
  assign s1506  = a1506 ^ b1506 ^ c1506;
  assign sub1506 = a1506 ^ b_inv1506 ^ c1506;
  assign and1506 = a1506 & b1506;
  assign or1506  = a1506 | b1506;
  assign c1507 = (a1506 & b1506) | (a1506 & c1506) | (b1506 & c1506);
  wire c_sub1507;
  assign c_sub1507 = (a1506 & b_inv1506) | (a1506 & c1506) | (b_inv1506 & c1506);
  wire s1507, sub1507, and1507, or1507;
  wire b_inv1507;
  assign b_inv1507 = ~b1507;
  assign s1507  = a1507 ^ b1507 ^ c1507;
  assign sub1507 = a1507 ^ b_inv1507 ^ c1507;
  assign and1507 = a1507 & b1507;
  assign or1507  = a1507 | b1507;
  assign c1508 = (a1507 & b1507) | (a1507 & c1507) | (b1507 & c1507);
  wire c_sub1508;
  assign c_sub1508 = (a1507 & b_inv1507) | (a1507 & c1507) | (b_inv1507 & c1507);
  wire s1508, sub1508, and1508, or1508;
  wire b_inv1508;
  assign b_inv1508 = ~b1508;
  assign s1508  = a1508 ^ b1508 ^ c1508;
  assign sub1508 = a1508 ^ b_inv1508 ^ c1508;
  assign and1508 = a1508 & b1508;
  assign or1508  = a1508 | b1508;
  assign c1509 = (a1508 & b1508) | (a1508 & c1508) | (b1508 & c1508);
  wire c_sub1509;
  assign c_sub1509 = (a1508 & b_inv1508) | (a1508 & c1508) | (b_inv1508 & c1508);
  wire s1509, sub1509, and1509, or1509;
  wire b_inv1509;
  assign b_inv1509 = ~b1509;
  assign s1509  = a1509 ^ b1509 ^ c1509;
  assign sub1509 = a1509 ^ b_inv1509 ^ c1509;
  assign and1509 = a1509 & b1509;
  assign or1509  = a1509 | b1509;
  assign c1510 = (a1509 & b1509) | (a1509 & c1509) | (b1509 & c1509);
  wire c_sub1510;
  assign c_sub1510 = (a1509 & b_inv1509) | (a1509 & c1509) | (b_inv1509 & c1509);
  wire s1510, sub1510, and1510, or1510;
  wire b_inv1510;
  assign b_inv1510 = ~b1510;
  assign s1510  = a1510 ^ b1510 ^ c1510;
  assign sub1510 = a1510 ^ b_inv1510 ^ c1510;
  assign and1510 = a1510 & b1510;
  assign or1510  = a1510 | b1510;
  assign c1511 = (a1510 & b1510) | (a1510 & c1510) | (b1510 & c1510);
  wire c_sub1511;
  assign c_sub1511 = (a1510 & b_inv1510) | (a1510 & c1510) | (b_inv1510 & c1510);
  wire s1511, sub1511, and1511, or1511;
  wire b_inv1511;
  assign b_inv1511 = ~b1511;
  assign s1511  = a1511 ^ b1511 ^ c1511;
  assign sub1511 = a1511 ^ b_inv1511 ^ c1511;
  assign and1511 = a1511 & b1511;
  assign or1511  = a1511 | b1511;
  assign c1512 = (a1511 & b1511) | (a1511 & c1511) | (b1511 & c1511);
  wire c_sub1512;
  assign c_sub1512 = (a1511 & b_inv1511) | (a1511 & c1511) | (b_inv1511 & c1511);
  wire s1512, sub1512, and1512, or1512;
  wire b_inv1512;
  assign b_inv1512 = ~b1512;
  assign s1512  = a1512 ^ b1512 ^ c1512;
  assign sub1512 = a1512 ^ b_inv1512 ^ c1512;
  assign and1512 = a1512 & b1512;
  assign or1512  = a1512 | b1512;
  assign c1513 = (a1512 & b1512) | (a1512 & c1512) | (b1512 & c1512);
  wire c_sub1513;
  assign c_sub1513 = (a1512 & b_inv1512) | (a1512 & c1512) | (b_inv1512 & c1512);
  wire s1513, sub1513, and1513, or1513;
  wire b_inv1513;
  assign b_inv1513 = ~b1513;
  assign s1513  = a1513 ^ b1513 ^ c1513;
  assign sub1513 = a1513 ^ b_inv1513 ^ c1513;
  assign and1513 = a1513 & b1513;
  assign or1513  = a1513 | b1513;
  assign c1514 = (a1513 & b1513) | (a1513 & c1513) | (b1513 & c1513);
  wire c_sub1514;
  assign c_sub1514 = (a1513 & b_inv1513) | (a1513 & c1513) | (b_inv1513 & c1513);
  wire s1514, sub1514, and1514, or1514;
  wire b_inv1514;
  assign b_inv1514 = ~b1514;
  assign s1514  = a1514 ^ b1514 ^ c1514;
  assign sub1514 = a1514 ^ b_inv1514 ^ c1514;
  assign and1514 = a1514 & b1514;
  assign or1514  = a1514 | b1514;
  assign c1515 = (a1514 & b1514) | (a1514 & c1514) | (b1514 & c1514);
  wire c_sub1515;
  assign c_sub1515 = (a1514 & b_inv1514) | (a1514 & c1514) | (b_inv1514 & c1514);
  wire s1515, sub1515, and1515, or1515;
  wire b_inv1515;
  assign b_inv1515 = ~b1515;
  assign s1515  = a1515 ^ b1515 ^ c1515;
  assign sub1515 = a1515 ^ b_inv1515 ^ c1515;
  assign and1515 = a1515 & b1515;
  assign or1515  = a1515 | b1515;
  assign c1516 = (a1515 & b1515) | (a1515 & c1515) | (b1515 & c1515);
  wire c_sub1516;
  assign c_sub1516 = (a1515 & b_inv1515) | (a1515 & c1515) | (b_inv1515 & c1515);
  wire s1516, sub1516, and1516, or1516;
  wire b_inv1516;
  assign b_inv1516 = ~b1516;
  assign s1516  = a1516 ^ b1516 ^ c1516;
  assign sub1516 = a1516 ^ b_inv1516 ^ c1516;
  assign and1516 = a1516 & b1516;
  assign or1516  = a1516 | b1516;
  assign c1517 = (a1516 & b1516) | (a1516 & c1516) | (b1516 & c1516);
  wire c_sub1517;
  assign c_sub1517 = (a1516 & b_inv1516) | (a1516 & c1516) | (b_inv1516 & c1516);
  wire s1517, sub1517, and1517, or1517;
  wire b_inv1517;
  assign b_inv1517 = ~b1517;
  assign s1517  = a1517 ^ b1517 ^ c1517;
  assign sub1517 = a1517 ^ b_inv1517 ^ c1517;
  assign and1517 = a1517 & b1517;
  assign or1517  = a1517 | b1517;
  assign c1518 = (a1517 & b1517) | (a1517 & c1517) | (b1517 & c1517);
  wire c_sub1518;
  assign c_sub1518 = (a1517 & b_inv1517) | (a1517 & c1517) | (b_inv1517 & c1517);
  wire s1518, sub1518, and1518, or1518;
  wire b_inv1518;
  assign b_inv1518 = ~b1518;
  assign s1518  = a1518 ^ b1518 ^ c1518;
  assign sub1518 = a1518 ^ b_inv1518 ^ c1518;
  assign and1518 = a1518 & b1518;
  assign or1518  = a1518 | b1518;
  assign c1519 = (a1518 & b1518) | (a1518 & c1518) | (b1518 & c1518);
  wire c_sub1519;
  assign c_sub1519 = (a1518 & b_inv1518) | (a1518 & c1518) | (b_inv1518 & c1518);
  wire s1519, sub1519, and1519, or1519;
  wire b_inv1519;
  assign b_inv1519 = ~b1519;
  assign s1519  = a1519 ^ b1519 ^ c1519;
  assign sub1519 = a1519 ^ b_inv1519 ^ c1519;
  assign and1519 = a1519 & b1519;
  assign or1519  = a1519 | b1519;
  assign c1520 = (a1519 & b1519) | (a1519 & c1519) | (b1519 & c1519);
  wire c_sub1520;
  assign c_sub1520 = (a1519 & b_inv1519) | (a1519 & c1519) | (b_inv1519 & c1519);
  wire s1520, sub1520, and1520, or1520;
  wire b_inv1520;
  assign b_inv1520 = ~b1520;
  assign s1520  = a1520 ^ b1520 ^ c1520;
  assign sub1520 = a1520 ^ b_inv1520 ^ c1520;
  assign and1520 = a1520 & b1520;
  assign or1520  = a1520 | b1520;
  assign c1521 = (a1520 & b1520) | (a1520 & c1520) | (b1520 & c1520);
  wire c_sub1521;
  assign c_sub1521 = (a1520 & b_inv1520) | (a1520 & c1520) | (b_inv1520 & c1520);
  wire s1521, sub1521, and1521, or1521;
  wire b_inv1521;
  assign b_inv1521 = ~b1521;
  assign s1521  = a1521 ^ b1521 ^ c1521;
  assign sub1521 = a1521 ^ b_inv1521 ^ c1521;
  assign and1521 = a1521 & b1521;
  assign or1521  = a1521 | b1521;
  assign c1522 = (a1521 & b1521) | (a1521 & c1521) | (b1521 & c1521);
  wire c_sub1522;
  assign c_sub1522 = (a1521 & b_inv1521) | (a1521 & c1521) | (b_inv1521 & c1521);
  wire s1522, sub1522, and1522, or1522;
  wire b_inv1522;
  assign b_inv1522 = ~b1522;
  assign s1522  = a1522 ^ b1522 ^ c1522;
  assign sub1522 = a1522 ^ b_inv1522 ^ c1522;
  assign and1522 = a1522 & b1522;
  assign or1522  = a1522 | b1522;
  assign c1523 = (a1522 & b1522) | (a1522 & c1522) | (b1522 & c1522);
  wire c_sub1523;
  assign c_sub1523 = (a1522 & b_inv1522) | (a1522 & c1522) | (b_inv1522 & c1522);
  wire s1523, sub1523, and1523, or1523;
  wire b_inv1523;
  assign b_inv1523 = ~b1523;
  assign s1523  = a1523 ^ b1523 ^ c1523;
  assign sub1523 = a1523 ^ b_inv1523 ^ c1523;
  assign and1523 = a1523 & b1523;
  assign or1523  = a1523 | b1523;
  assign c1524 = (a1523 & b1523) | (a1523 & c1523) | (b1523 & c1523);
  wire c_sub1524;
  assign c_sub1524 = (a1523 & b_inv1523) | (a1523 & c1523) | (b_inv1523 & c1523);
  wire s1524, sub1524, and1524, or1524;
  wire b_inv1524;
  assign b_inv1524 = ~b1524;
  assign s1524  = a1524 ^ b1524 ^ c1524;
  assign sub1524 = a1524 ^ b_inv1524 ^ c1524;
  assign and1524 = a1524 & b1524;
  assign or1524  = a1524 | b1524;
  assign c1525 = (a1524 & b1524) | (a1524 & c1524) | (b1524 & c1524);
  wire c_sub1525;
  assign c_sub1525 = (a1524 & b_inv1524) | (a1524 & c1524) | (b_inv1524 & c1524);
  wire s1525, sub1525, and1525, or1525;
  wire b_inv1525;
  assign b_inv1525 = ~b1525;
  assign s1525  = a1525 ^ b1525 ^ c1525;
  assign sub1525 = a1525 ^ b_inv1525 ^ c1525;
  assign and1525 = a1525 & b1525;
  assign or1525  = a1525 | b1525;
  assign c1526 = (a1525 & b1525) | (a1525 & c1525) | (b1525 & c1525);
  wire c_sub1526;
  assign c_sub1526 = (a1525 & b_inv1525) | (a1525 & c1525) | (b_inv1525 & c1525);
  wire s1526, sub1526, and1526, or1526;
  wire b_inv1526;
  assign b_inv1526 = ~b1526;
  assign s1526  = a1526 ^ b1526 ^ c1526;
  assign sub1526 = a1526 ^ b_inv1526 ^ c1526;
  assign and1526 = a1526 & b1526;
  assign or1526  = a1526 | b1526;
  assign c1527 = (a1526 & b1526) | (a1526 & c1526) | (b1526 & c1526);
  wire c_sub1527;
  assign c_sub1527 = (a1526 & b_inv1526) | (a1526 & c1526) | (b_inv1526 & c1526);
  wire s1527, sub1527, and1527, or1527;
  wire b_inv1527;
  assign b_inv1527 = ~b1527;
  assign s1527  = a1527 ^ b1527 ^ c1527;
  assign sub1527 = a1527 ^ b_inv1527 ^ c1527;
  assign and1527 = a1527 & b1527;
  assign or1527  = a1527 | b1527;
  assign c1528 = (a1527 & b1527) | (a1527 & c1527) | (b1527 & c1527);
  wire c_sub1528;
  assign c_sub1528 = (a1527 & b_inv1527) | (a1527 & c1527) | (b_inv1527 & c1527);
  wire s1528, sub1528, and1528, or1528;
  wire b_inv1528;
  assign b_inv1528 = ~b1528;
  assign s1528  = a1528 ^ b1528 ^ c1528;
  assign sub1528 = a1528 ^ b_inv1528 ^ c1528;
  assign and1528 = a1528 & b1528;
  assign or1528  = a1528 | b1528;
  assign c1529 = (a1528 & b1528) | (a1528 & c1528) | (b1528 & c1528);
  wire c_sub1529;
  assign c_sub1529 = (a1528 & b_inv1528) | (a1528 & c1528) | (b_inv1528 & c1528);
  wire s1529, sub1529, and1529, or1529;
  wire b_inv1529;
  assign b_inv1529 = ~b1529;
  assign s1529  = a1529 ^ b1529 ^ c1529;
  assign sub1529 = a1529 ^ b_inv1529 ^ c1529;
  assign and1529 = a1529 & b1529;
  assign or1529  = a1529 | b1529;
  assign c1530 = (a1529 & b1529) | (a1529 & c1529) | (b1529 & c1529);
  wire c_sub1530;
  assign c_sub1530 = (a1529 & b_inv1529) | (a1529 & c1529) | (b_inv1529 & c1529);
  wire s1530, sub1530, and1530, or1530;
  wire b_inv1530;
  assign b_inv1530 = ~b1530;
  assign s1530  = a1530 ^ b1530 ^ c1530;
  assign sub1530 = a1530 ^ b_inv1530 ^ c1530;
  assign and1530 = a1530 & b1530;
  assign or1530  = a1530 | b1530;
  assign c1531 = (a1530 & b1530) | (a1530 & c1530) | (b1530 & c1530);
  wire c_sub1531;
  assign c_sub1531 = (a1530 & b_inv1530) | (a1530 & c1530) | (b_inv1530 & c1530);
  wire s1531, sub1531, and1531, or1531;
  wire b_inv1531;
  assign b_inv1531 = ~b1531;
  assign s1531  = a1531 ^ b1531 ^ c1531;
  assign sub1531 = a1531 ^ b_inv1531 ^ c1531;
  assign and1531 = a1531 & b1531;
  assign or1531  = a1531 | b1531;
  assign c1532 = (a1531 & b1531) | (a1531 & c1531) | (b1531 & c1531);
  wire c_sub1532;
  assign c_sub1532 = (a1531 & b_inv1531) | (a1531 & c1531) | (b_inv1531 & c1531);
  wire s1532, sub1532, and1532, or1532;
  wire b_inv1532;
  assign b_inv1532 = ~b1532;
  assign s1532  = a1532 ^ b1532 ^ c1532;
  assign sub1532 = a1532 ^ b_inv1532 ^ c1532;
  assign and1532 = a1532 & b1532;
  assign or1532  = a1532 | b1532;
  assign c1533 = (a1532 & b1532) | (a1532 & c1532) | (b1532 & c1532);
  wire c_sub1533;
  assign c_sub1533 = (a1532 & b_inv1532) | (a1532 & c1532) | (b_inv1532 & c1532);
  wire s1533, sub1533, and1533, or1533;
  wire b_inv1533;
  assign b_inv1533 = ~b1533;
  assign s1533  = a1533 ^ b1533 ^ c1533;
  assign sub1533 = a1533 ^ b_inv1533 ^ c1533;
  assign and1533 = a1533 & b1533;
  assign or1533  = a1533 | b1533;
  assign c1534 = (a1533 & b1533) | (a1533 & c1533) | (b1533 & c1533);
  wire c_sub1534;
  assign c_sub1534 = (a1533 & b_inv1533) | (a1533 & c1533) | (b_inv1533 & c1533);
  wire s1534, sub1534, and1534, or1534;
  wire b_inv1534;
  assign b_inv1534 = ~b1534;
  assign s1534  = a1534 ^ b1534 ^ c1534;
  assign sub1534 = a1534 ^ b_inv1534 ^ c1534;
  assign and1534 = a1534 & b1534;
  assign or1534  = a1534 | b1534;
  assign c1535 = (a1534 & b1534) | (a1534 & c1534) | (b1534 & c1534);
  wire c_sub1535;
  assign c_sub1535 = (a1534 & b_inv1534) | (a1534 & c1534) | (b_inv1534 & c1534);
  wire s1535, sub1535, and1535, or1535;
  wire b_inv1535;
  assign b_inv1535 = ~b1535;
  assign s1535  = a1535 ^ b1535 ^ c1535;
  assign sub1535 = a1535 ^ b_inv1535 ^ c1535;
  assign and1535 = a1535 & b1535;
  assign or1535  = a1535 | b1535;
  assign c1536 = (a1535 & b1535) | (a1535 & c1535) | (b1535 & c1535);
  wire c_sub1536;
  assign c_sub1536 = (a1535 & b_inv1535) | (a1535 & c1535) | (b_inv1535 & c1535);
  wire s1536, sub1536, and1536, or1536;
  wire b_inv1536;
  assign b_inv1536 = ~b1536;
  assign s1536  = a1536 ^ b1536 ^ c1536;
  assign sub1536 = a1536 ^ b_inv1536 ^ c1536;
  assign and1536 = a1536 & b1536;
  assign or1536  = a1536 | b1536;
  assign c1537 = (a1536 & b1536) | (a1536 & c1536) | (b1536 & c1536);
  wire c_sub1537;
  assign c_sub1537 = (a1536 & b_inv1536) | (a1536 & c1536) | (b_inv1536 & c1536);
  wire s1537, sub1537, and1537, or1537;
  wire b_inv1537;
  assign b_inv1537 = ~b1537;
  assign s1537  = a1537 ^ b1537 ^ c1537;
  assign sub1537 = a1537 ^ b_inv1537 ^ c1537;
  assign and1537 = a1537 & b1537;
  assign or1537  = a1537 | b1537;
  assign c1538 = (a1537 & b1537) | (a1537 & c1537) | (b1537 & c1537);
  wire c_sub1538;
  assign c_sub1538 = (a1537 & b_inv1537) | (a1537 & c1537) | (b_inv1537 & c1537);
  wire s1538, sub1538, and1538, or1538;
  wire b_inv1538;
  assign b_inv1538 = ~b1538;
  assign s1538  = a1538 ^ b1538 ^ c1538;
  assign sub1538 = a1538 ^ b_inv1538 ^ c1538;
  assign and1538 = a1538 & b1538;
  assign or1538  = a1538 | b1538;
  assign c1539 = (a1538 & b1538) | (a1538 & c1538) | (b1538 & c1538);
  wire c_sub1539;
  assign c_sub1539 = (a1538 & b_inv1538) | (a1538 & c1538) | (b_inv1538 & c1538);
  wire s1539, sub1539, and1539, or1539;
  wire b_inv1539;
  assign b_inv1539 = ~b1539;
  assign s1539  = a1539 ^ b1539 ^ c1539;
  assign sub1539 = a1539 ^ b_inv1539 ^ c1539;
  assign and1539 = a1539 & b1539;
  assign or1539  = a1539 | b1539;
  assign c1540 = (a1539 & b1539) | (a1539 & c1539) | (b1539 & c1539);
  wire c_sub1540;
  assign c_sub1540 = (a1539 & b_inv1539) | (a1539 & c1539) | (b_inv1539 & c1539);
  wire s1540, sub1540, and1540, or1540;
  wire b_inv1540;
  assign b_inv1540 = ~b1540;
  assign s1540  = a1540 ^ b1540 ^ c1540;
  assign sub1540 = a1540 ^ b_inv1540 ^ c1540;
  assign and1540 = a1540 & b1540;
  assign or1540  = a1540 | b1540;
  assign c1541 = (a1540 & b1540) | (a1540 & c1540) | (b1540 & c1540);
  wire c_sub1541;
  assign c_sub1541 = (a1540 & b_inv1540) | (a1540 & c1540) | (b_inv1540 & c1540);
  wire s1541, sub1541, and1541, or1541;
  wire b_inv1541;
  assign b_inv1541 = ~b1541;
  assign s1541  = a1541 ^ b1541 ^ c1541;
  assign sub1541 = a1541 ^ b_inv1541 ^ c1541;
  assign and1541 = a1541 & b1541;
  assign or1541  = a1541 | b1541;
  assign c1542 = (a1541 & b1541) | (a1541 & c1541) | (b1541 & c1541);
  wire c_sub1542;
  assign c_sub1542 = (a1541 & b_inv1541) | (a1541 & c1541) | (b_inv1541 & c1541);
  wire s1542, sub1542, and1542, or1542;
  wire b_inv1542;
  assign b_inv1542 = ~b1542;
  assign s1542  = a1542 ^ b1542 ^ c1542;
  assign sub1542 = a1542 ^ b_inv1542 ^ c1542;
  assign and1542 = a1542 & b1542;
  assign or1542  = a1542 | b1542;
  assign c1543 = (a1542 & b1542) | (a1542 & c1542) | (b1542 & c1542);
  wire c_sub1543;
  assign c_sub1543 = (a1542 & b_inv1542) | (a1542 & c1542) | (b_inv1542 & c1542);
  wire s1543, sub1543, and1543, or1543;
  wire b_inv1543;
  assign b_inv1543 = ~b1543;
  assign s1543  = a1543 ^ b1543 ^ c1543;
  assign sub1543 = a1543 ^ b_inv1543 ^ c1543;
  assign and1543 = a1543 & b1543;
  assign or1543  = a1543 | b1543;
  assign c1544 = (a1543 & b1543) | (a1543 & c1543) | (b1543 & c1543);
  wire c_sub1544;
  assign c_sub1544 = (a1543 & b_inv1543) | (a1543 & c1543) | (b_inv1543 & c1543);
  wire s1544, sub1544, and1544, or1544;
  wire b_inv1544;
  assign b_inv1544 = ~b1544;
  assign s1544  = a1544 ^ b1544 ^ c1544;
  assign sub1544 = a1544 ^ b_inv1544 ^ c1544;
  assign and1544 = a1544 & b1544;
  assign or1544  = a1544 | b1544;
  assign c1545 = (a1544 & b1544) | (a1544 & c1544) | (b1544 & c1544);
  wire c_sub1545;
  assign c_sub1545 = (a1544 & b_inv1544) | (a1544 & c1544) | (b_inv1544 & c1544);
  wire s1545, sub1545, and1545, or1545;
  wire b_inv1545;
  assign b_inv1545 = ~b1545;
  assign s1545  = a1545 ^ b1545 ^ c1545;
  assign sub1545 = a1545 ^ b_inv1545 ^ c1545;
  assign and1545 = a1545 & b1545;
  assign or1545  = a1545 | b1545;
  assign c1546 = (a1545 & b1545) | (a1545 & c1545) | (b1545 & c1545);
  wire c_sub1546;
  assign c_sub1546 = (a1545 & b_inv1545) | (a1545 & c1545) | (b_inv1545 & c1545);
  wire s1546, sub1546, and1546, or1546;
  wire b_inv1546;
  assign b_inv1546 = ~b1546;
  assign s1546  = a1546 ^ b1546 ^ c1546;
  assign sub1546 = a1546 ^ b_inv1546 ^ c1546;
  assign and1546 = a1546 & b1546;
  assign or1546  = a1546 | b1546;
  assign c1547 = (a1546 & b1546) | (a1546 & c1546) | (b1546 & c1546);
  wire c_sub1547;
  assign c_sub1547 = (a1546 & b_inv1546) | (a1546 & c1546) | (b_inv1546 & c1546);
  wire s1547, sub1547, and1547, or1547;
  wire b_inv1547;
  assign b_inv1547 = ~b1547;
  assign s1547  = a1547 ^ b1547 ^ c1547;
  assign sub1547 = a1547 ^ b_inv1547 ^ c1547;
  assign and1547 = a1547 & b1547;
  assign or1547  = a1547 | b1547;
  assign c1548 = (a1547 & b1547) | (a1547 & c1547) | (b1547 & c1547);
  wire c_sub1548;
  assign c_sub1548 = (a1547 & b_inv1547) | (a1547 & c1547) | (b_inv1547 & c1547);
  wire s1548, sub1548, and1548, or1548;
  wire b_inv1548;
  assign b_inv1548 = ~b1548;
  assign s1548  = a1548 ^ b1548 ^ c1548;
  assign sub1548 = a1548 ^ b_inv1548 ^ c1548;
  assign and1548 = a1548 & b1548;
  assign or1548  = a1548 | b1548;
  assign c1549 = (a1548 & b1548) | (a1548 & c1548) | (b1548 & c1548);
  wire c_sub1549;
  assign c_sub1549 = (a1548 & b_inv1548) | (a1548 & c1548) | (b_inv1548 & c1548);
  wire s1549, sub1549, and1549, or1549;
  wire b_inv1549;
  assign b_inv1549 = ~b1549;
  assign s1549  = a1549 ^ b1549 ^ c1549;
  assign sub1549 = a1549 ^ b_inv1549 ^ c1549;
  assign and1549 = a1549 & b1549;
  assign or1549  = a1549 | b1549;
  assign c1550 = (a1549 & b1549) | (a1549 & c1549) | (b1549 & c1549);
  wire c_sub1550;
  assign c_sub1550 = (a1549 & b_inv1549) | (a1549 & c1549) | (b_inv1549 & c1549);
  wire s1550, sub1550, and1550, or1550;
  wire b_inv1550;
  assign b_inv1550 = ~b1550;
  assign s1550  = a1550 ^ b1550 ^ c1550;
  assign sub1550 = a1550 ^ b_inv1550 ^ c1550;
  assign and1550 = a1550 & b1550;
  assign or1550  = a1550 | b1550;
  assign c1551 = (a1550 & b1550) | (a1550 & c1550) | (b1550 & c1550);
  wire c_sub1551;
  assign c_sub1551 = (a1550 & b_inv1550) | (a1550 & c1550) | (b_inv1550 & c1550);
  wire s1551, sub1551, and1551, or1551;
  wire b_inv1551;
  assign b_inv1551 = ~b1551;
  assign s1551  = a1551 ^ b1551 ^ c1551;
  assign sub1551 = a1551 ^ b_inv1551 ^ c1551;
  assign and1551 = a1551 & b1551;
  assign or1551  = a1551 | b1551;
  assign c1552 = (a1551 & b1551) | (a1551 & c1551) | (b1551 & c1551);
  wire c_sub1552;
  assign c_sub1552 = (a1551 & b_inv1551) | (a1551 & c1551) | (b_inv1551 & c1551);
  wire s1552, sub1552, and1552, or1552;
  wire b_inv1552;
  assign b_inv1552 = ~b1552;
  assign s1552  = a1552 ^ b1552 ^ c1552;
  assign sub1552 = a1552 ^ b_inv1552 ^ c1552;
  assign and1552 = a1552 & b1552;
  assign or1552  = a1552 | b1552;
  assign c1553 = (a1552 & b1552) | (a1552 & c1552) | (b1552 & c1552);
  wire c_sub1553;
  assign c_sub1553 = (a1552 & b_inv1552) | (a1552 & c1552) | (b_inv1552 & c1552);
  wire s1553, sub1553, and1553, or1553;
  wire b_inv1553;
  assign b_inv1553 = ~b1553;
  assign s1553  = a1553 ^ b1553 ^ c1553;
  assign sub1553 = a1553 ^ b_inv1553 ^ c1553;
  assign and1553 = a1553 & b1553;
  assign or1553  = a1553 | b1553;
  assign c1554 = (a1553 & b1553) | (a1553 & c1553) | (b1553 & c1553);
  wire c_sub1554;
  assign c_sub1554 = (a1553 & b_inv1553) | (a1553 & c1553) | (b_inv1553 & c1553);
  wire s1554, sub1554, and1554, or1554;
  wire b_inv1554;
  assign b_inv1554 = ~b1554;
  assign s1554  = a1554 ^ b1554 ^ c1554;
  assign sub1554 = a1554 ^ b_inv1554 ^ c1554;
  assign and1554 = a1554 & b1554;
  assign or1554  = a1554 | b1554;
  assign c1555 = (a1554 & b1554) | (a1554 & c1554) | (b1554 & c1554);
  wire c_sub1555;
  assign c_sub1555 = (a1554 & b_inv1554) | (a1554 & c1554) | (b_inv1554 & c1554);
  wire s1555, sub1555, and1555, or1555;
  wire b_inv1555;
  assign b_inv1555 = ~b1555;
  assign s1555  = a1555 ^ b1555 ^ c1555;
  assign sub1555 = a1555 ^ b_inv1555 ^ c1555;
  assign and1555 = a1555 & b1555;
  assign or1555  = a1555 | b1555;
  assign c1556 = (a1555 & b1555) | (a1555 & c1555) | (b1555 & c1555);
  wire c_sub1556;
  assign c_sub1556 = (a1555 & b_inv1555) | (a1555 & c1555) | (b_inv1555 & c1555);
  wire s1556, sub1556, and1556, or1556;
  wire b_inv1556;
  assign b_inv1556 = ~b1556;
  assign s1556  = a1556 ^ b1556 ^ c1556;
  assign sub1556 = a1556 ^ b_inv1556 ^ c1556;
  assign and1556 = a1556 & b1556;
  assign or1556  = a1556 | b1556;
  assign c1557 = (a1556 & b1556) | (a1556 & c1556) | (b1556 & c1556);
  wire c_sub1557;
  assign c_sub1557 = (a1556 & b_inv1556) | (a1556 & c1556) | (b_inv1556 & c1556);
  wire s1557, sub1557, and1557, or1557;
  wire b_inv1557;
  assign b_inv1557 = ~b1557;
  assign s1557  = a1557 ^ b1557 ^ c1557;
  assign sub1557 = a1557 ^ b_inv1557 ^ c1557;
  assign and1557 = a1557 & b1557;
  assign or1557  = a1557 | b1557;
  assign c1558 = (a1557 & b1557) | (a1557 & c1557) | (b1557 & c1557);
  wire c_sub1558;
  assign c_sub1558 = (a1557 & b_inv1557) | (a1557 & c1557) | (b_inv1557 & c1557);
  wire s1558, sub1558, and1558, or1558;
  wire b_inv1558;
  assign b_inv1558 = ~b1558;
  assign s1558  = a1558 ^ b1558 ^ c1558;
  assign sub1558 = a1558 ^ b_inv1558 ^ c1558;
  assign and1558 = a1558 & b1558;
  assign or1558  = a1558 | b1558;
  assign c1559 = (a1558 & b1558) | (a1558 & c1558) | (b1558 & c1558);
  wire c_sub1559;
  assign c_sub1559 = (a1558 & b_inv1558) | (a1558 & c1558) | (b_inv1558 & c1558);
  wire s1559, sub1559, and1559, or1559;
  wire b_inv1559;
  assign b_inv1559 = ~b1559;
  assign s1559  = a1559 ^ b1559 ^ c1559;
  assign sub1559 = a1559 ^ b_inv1559 ^ c1559;
  assign and1559 = a1559 & b1559;
  assign or1559  = a1559 | b1559;
  assign c1560 = (a1559 & b1559) | (a1559 & c1559) | (b1559 & c1559);
  wire c_sub1560;
  assign c_sub1560 = (a1559 & b_inv1559) | (a1559 & c1559) | (b_inv1559 & c1559);
  wire s1560, sub1560, and1560, or1560;
  wire b_inv1560;
  assign b_inv1560 = ~b1560;
  assign s1560  = a1560 ^ b1560 ^ c1560;
  assign sub1560 = a1560 ^ b_inv1560 ^ c1560;
  assign and1560 = a1560 & b1560;
  assign or1560  = a1560 | b1560;
  assign c1561 = (a1560 & b1560) | (a1560 & c1560) | (b1560 & c1560);
  wire c_sub1561;
  assign c_sub1561 = (a1560 & b_inv1560) | (a1560 & c1560) | (b_inv1560 & c1560);
  wire s1561, sub1561, and1561, or1561;
  wire b_inv1561;
  assign b_inv1561 = ~b1561;
  assign s1561  = a1561 ^ b1561 ^ c1561;
  assign sub1561 = a1561 ^ b_inv1561 ^ c1561;
  assign and1561 = a1561 & b1561;
  assign or1561  = a1561 | b1561;
  assign c1562 = (a1561 & b1561) | (a1561 & c1561) | (b1561 & c1561);
  wire c_sub1562;
  assign c_sub1562 = (a1561 & b_inv1561) | (a1561 & c1561) | (b_inv1561 & c1561);
  wire s1562, sub1562, and1562, or1562;
  wire b_inv1562;
  assign b_inv1562 = ~b1562;
  assign s1562  = a1562 ^ b1562 ^ c1562;
  assign sub1562 = a1562 ^ b_inv1562 ^ c1562;
  assign and1562 = a1562 & b1562;
  assign or1562  = a1562 | b1562;
  assign c1563 = (a1562 & b1562) | (a1562 & c1562) | (b1562 & c1562);
  wire c_sub1563;
  assign c_sub1563 = (a1562 & b_inv1562) | (a1562 & c1562) | (b_inv1562 & c1562);
  wire s1563, sub1563, and1563, or1563;
  wire b_inv1563;
  assign b_inv1563 = ~b1563;
  assign s1563  = a1563 ^ b1563 ^ c1563;
  assign sub1563 = a1563 ^ b_inv1563 ^ c1563;
  assign and1563 = a1563 & b1563;
  assign or1563  = a1563 | b1563;
  assign c1564 = (a1563 & b1563) | (a1563 & c1563) | (b1563 & c1563);
  wire c_sub1564;
  assign c_sub1564 = (a1563 & b_inv1563) | (a1563 & c1563) | (b_inv1563 & c1563);
  wire s1564, sub1564, and1564, or1564;
  wire b_inv1564;
  assign b_inv1564 = ~b1564;
  assign s1564  = a1564 ^ b1564 ^ c1564;
  assign sub1564 = a1564 ^ b_inv1564 ^ c1564;
  assign and1564 = a1564 & b1564;
  assign or1564  = a1564 | b1564;
  assign c1565 = (a1564 & b1564) | (a1564 & c1564) | (b1564 & c1564);
  wire c_sub1565;
  assign c_sub1565 = (a1564 & b_inv1564) | (a1564 & c1564) | (b_inv1564 & c1564);
  wire s1565, sub1565, and1565, or1565;
  wire b_inv1565;
  assign b_inv1565 = ~b1565;
  assign s1565  = a1565 ^ b1565 ^ c1565;
  assign sub1565 = a1565 ^ b_inv1565 ^ c1565;
  assign and1565 = a1565 & b1565;
  assign or1565  = a1565 | b1565;
  assign c1566 = (a1565 & b1565) | (a1565 & c1565) | (b1565 & c1565);
  wire c_sub1566;
  assign c_sub1566 = (a1565 & b_inv1565) | (a1565 & c1565) | (b_inv1565 & c1565);
  wire s1566, sub1566, and1566, or1566;
  wire b_inv1566;
  assign b_inv1566 = ~b1566;
  assign s1566  = a1566 ^ b1566 ^ c1566;
  assign sub1566 = a1566 ^ b_inv1566 ^ c1566;
  assign and1566 = a1566 & b1566;
  assign or1566  = a1566 | b1566;
  assign c1567 = (a1566 & b1566) | (a1566 & c1566) | (b1566 & c1566);
  wire c_sub1567;
  assign c_sub1567 = (a1566 & b_inv1566) | (a1566 & c1566) | (b_inv1566 & c1566);
  wire s1567, sub1567, and1567, or1567;
  wire b_inv1567;
  assign b_inv1567 = ~b1567;
  assign s1567  = a1567 ^ b1567 ^ c1567;
  assign sub1567 = a1567 ^ b_inv1567 ^ c1567;
  assign and1567 = a1567 & b1567;
  assign or1567  = a1567 | b1567;
  assign c1568 = (a1567 & b1567) | (a1567 & c1567) | (b1567 & c1567);
  wire c_sub1568;
  assign c_sub1568 = (a1567 & b_inv1567) | (a1567 & c1567) | (b_inv1567 & c1567);
  wire s1568, sub1568, and1568, or1568;
  wire b_inv1568;
  assign b_inv1568 = ~b1568;
  assign s1568  = a1568 ^ b1568 ^ c1568;
  assign sub1568 = a1568 ^ b_inv1568 ^ c1568;
  assign and1568 = a1568 & b1568;
  assign or1568  = a1568 | b1568;
  assign c1569 = (a1568 & b1568) | (a1568 & c1568) | (b1568 & c1568);
  wire c_sub1569;
  assign c_sub1569 = (a1568 & b_inv1568) | (a1568 & c1568) | (b_inv1568 & c1568);
  wire s1569, sub1569, and1569, or1569;
  wire b_inv1569;
  assign b_inv1569 = ~b1569;
  assign s1569  = a1569 ^ b1569 ^ c1569;
  assign sub1569 = a1569 ^ b_inv1569 ^ c1569;
  assign and1569 = a1569 & b1569;
  assign or1569  = a1569 | b1569;
  assign c1570 = (a1569 & b1569) | (a1569 & c1569) | (b1569 & c1569);
  wire c_sub1570;
  assign c_sub1570 = (a1569 & b_inv1569) | (a1569 & c1569) | (b_inv1569 & c1569);
  wire s1570, sub1570, and1570, or1570;
  wire b_inv1570;
  assign b_inv1570 = ~b1570;
  assign s1570  = a1570 ^ b1570 ^ c1570;
  assign sub1570 = a1570 ^ b_inv1570 ^ c1570;
  assign and1570 = a1570 & b1570;
  assign or1570  = a1570 | b1570;
  assign c1571 = (a1570 & b1570) | (a1570 & c1570) | (b1570 & c1570);
  wire c_sub1571;
  assign c_sub1571 = (a1570 & b_inv1570) | (a1570 & c1570) | (b_inv1570 & c1570);
  wire s1571, sub1571, and1571, or1571;
  wire b_inv1571;
  assign b_inv1571 = ~b1571;
  assign s1571  = a1571 ^ b1571 ^ c1571;
  assign sub1571 = a1571 ^ b_inv1571 ^ c1571;
  assign and1571 = a1571 & b1571;
  assign or1571  = a1571 | b1571;
  assign c1572 = (a1571 & b1571) | (a1571 & c1571) | (b1571 & c1571);
  wire c_sub1572;
  assign c_sub1572 = (a1571 & b_inv1571) | (a1571 & c1571) | (b_inv1571 & c1571);
  wire s1572, sub1572, and1572, or1572;
  wire b_inv1572;
  assign b_inv1572 = ~b1572;
  assign s1572  = a1572 ^ b1572 ^ c1572;
  assign sub1572 = a1572 ^ b_inv1572 ^ c1572;
  assign and1572 = a1572 & b1572;
  assign or1572  = a1572 | b1572;
  assign c1573 = (a1572 & b1572) | (a1572 & c1572) | (b1572 & c1572);
  wire c_sub1573;
  assign c_sub1573 = (a1572 & b_inv1572) | (a1572 & c1572) | (b_inv1572 & c1572);
  wire s1573, sub1573, and1573, or1573;
  wire b_inv1573;
  assign b_inv1573 = ~b1573;
  assign s1573  = a1573 ^ b1573 ^ c1573;
  assign sub1573 = a1573 ^ b_inv1573 ^ c1573;
  assign and1573 = a1573 & b1573;
  assign or1573  = a1573 | b1573;
  assign c1574 = (a1573 & b1573) | (a1573 & c1573) | (b1573 & c1573);
  wire c_sub1574;
  assign c_sub1574 = (a1573 & b_inv1573) | (a1573 & c1573) | (b_inv1573 & c1573);
  wire s1574, sub1574, and1574, or1574;
  wire b_inv1574;
  assign b_inv1574 = ~b1574;
  assign s1574  = a1574 ^ b1574 ^ c1574;
  assign sub1574 = a1574 ^ b_inv1574 ^ c1574;
  assign and1574 = a1574 & b1574;
  assign or1574  = a1574 | b1574;
  assign c1575 = (a1574 & b1574) | (a1574 & c1574) | (b1574 & c1574);
  wire c_sub1575;
  assign c_sub1575 = (a1574 & b_inv1574) | (a1574 & c1574) | (b_inv1574 & c1574);
  wire s1575, sub1575, and1575, or1575;
  wire b_inv1575;
  assign b_inv1575 = ~b1575;
  assign s1575  = a1575 ^ b1575 ^ c1575;
  assign sub1575 = a1575 ^ b_inv1575 ^ c1575;
  assign and1575 = a1575 & b1575;
  assign or1575  = a1575 | b1575;
  assign c1576 = (a1575 & b1575) | (a1575 & c1575) | (b1575 & c1575);
  wire c_sub1576;
  assign c_sub1576 = (a1575 & b_inv1575) | (a1575 & c1575) | (b_inv1575 & c1575);
  wire s1576, sub1576, and1576, or1576;
  wire b_inv1576;
  assign b_inv1576 = ~b1576;
  assign s1576  = a1576 ^ b1576 ^ c1576;
  assign sub1576 = a1576 ^ b_inv1576 ^ c1576;
  assign and1576 = a1576 & b1576;
  assign or1576  = a1576 | b1576;
  assign c1577 = (a1576 & b1576) | (a1576 & c1576) | (b1576 & c1576);
  wire c_sub1577;
  assign c_sub1577 = (a1576 & b_inv1576) | (a1576 & c1576) | (b_inv1576 & c1576);
  wire s1577, sub1577, and1577, or1577;
  wire b_inv1577;
  assign b_inv1577 = ~b1577;
  assign s1577  = a1577 ^ b1577 ^ c1577;
  assign sub1577 = a1577 ^ b_inv1577 ^ c1577;
  assign and1577 = a1577 & b1577;
  assign or1577  = a1577 | b1577;
  assign c1578 = (a1577 & b1577) | (a1577 & c1577) | (b1577 & c1577);
  wire c_sub1578;
  assign c_sub1578 = (a1577 & b_inv1577) | (a1577 & c1577) | (b_inv1577 & c1577);
  wire s1578, sub1578, and1578, or1578;
  wire b_inv1578;
  assign b_inv1578 = ~b1578;
  assign s1578  = a1578 ^ b1578 ^ c1578;
  assign sub1578 = a1578 ^ b_inv1578 ^ c1578;
  assign and1578 = a1578 & b1578;
  assign or1578  = a1578 | b1578;
  assign c1579 = (a1578 & b1578) | (a1578 & c1578) | (b1578 & c1578);
  wire c_sub1579;
  assign c_sub1579 = (a1578 & b_inv1578) | (a1578 & c1578) | (b_inv1578 & c1578);
  wire s1579, sub1579, and1579, or1579;
  wire b_inv1579;
  assign b_inv1579 = ~b1579;
  assign s1579  = a1579 ^ b1579 ^ c1579;
  assign sub1579 = a1579 ^ b_inv1579 ^ c1579;
  assign and1579 = a1579 & b1579;
  assign or1579  = a1579 | b1579;
  assign c1580 = (a1579 & b1579) | (a1579 & c1579) | (b1579 & c1579);
  wire c_sub1580;
  assign c_sub1580 = (a1579 & b_inv1579) | (a1579 & c1579) | (b_inv1579 & c1579);
  wire s1580, sub1580, and1580, or1580;
  wire b_inv1580;
  assign b_inv1580 = ~b1580;
  assign s1580  = a1580 ^ b1580 ^ c1580;
  assign sub1580 = a1580 ^ b_inv1580 ^ c1580;
  assign and1580 = a1580 & b1580;
  assign or1580  = a1580 | b1580;
  assign c1581 = (a1580 & b1580) | (a1580 & c1580) | (b1580 & c1580);
  wire c_sub1581;
  assign c_sub1581 = (a1580 & b_inv1580) | (a1580 & c1580) | (b_inv1580 & c1580);
  wire s1581, sub1581, and1581, or1581;
  wire b_inv1581;
  assign b_inv1581 = ~b1581;
  assign s1581  = a1581 ^ b1581 ^ c1581;
  assign sub1581 = a1581 ^ b_inv1581 ^ c1581;
  assign and1581 = a1581 & b1581;
  assign or1581  = a1581 | b1581;
  assign c1582 = (a1581 & b1581) | (a1581 & c1581) | (b1581 & c1581);
  wire c_sub1582;
  assign c_sub1582 = (a1581 & b_inv1581) | (a1581 & c1581) | (b_inv1581 & c1581);
  wire s1582, sub1582, and1582, or1582;
  wire b_inv1582;
  assign b_inv1582 = ~b1582;
  assign s1582  = a1582 ^ b1582 ^ c1582;
  assign sub1582 = a1582 ^ b_inv1582 ^ c1582;
  assign and1582 = a1582 & b1582;
  assign or1582  = a1582 | b1582;
  assign c1583 = (a1582 & b1582) | (a1582 & c1582) | (b1582 & c1582);
  wire c_sub1583;
  assign c_sub1583 = (a1582 & b_inv1582) | (a1582 & c1582) | (b_inv1582 & c1582);
  wire s1583, sub1583, and1583, or1583;
  wire b_inv1583;
  assign b_inv1583 = ~b1583;
  assign s1583  = a1583 ^ b1583 ^ c1583;
  assign sub1583 = a1583 ^ b_inv1583 ^ c1583;
  assign and1583 = a1583 & b1583;
  assign or1583  = a1583 | b1583;
  assign c1584 = (a1583 & b1583) | (a1583 & c1583) | (b1583 & c1583);
  wire c_sub1584;
  assign c_sub1584 = (a1583 & b_inv1583) | (a1583 & c1583) | (b_inv1583 & c1583);
  wire s1584, sub1584, and1584, or1584;
  wire b_inv1584;
  assign b_inv1584 = ~b1584;
  assign s1584  = a1584 ^ b1584 ^ c1584;
  assign sub1584 = a1584 ^ b_inv1584 ^ c1584;
  assign and1584 = a1584 & b1584;
  assign or1584  = a1584 | b1584;
  assign c1585 = (a1584 & b1584) | (a1584 & c1584) | (b1584 & c1584);
  wire c_sub1585;
  assign c_sub1585 = (a1584 & b_inv1584) | (a1584 & c1584) | (b_inv1584 & c1584);
  wire s1585, sub1585, and1585, or1585;
  wire b_inv1585;
  assign b_inv1585 = ~b1585;
  assign s1585  = a1585 ^ b1585 ^ c1585;
  assign sub1585 = a1585 ^ b_inv1585 ^ c1585;
  assign and1585 = a1585 & b1585;
  assign or1585  = a1585 | b1585;
  assign c1586 = (a1585 & b1585) | (a1585 & c1585) | (b1585 & c1585);
  wire c_sub1586;
  assign c_sub1586 = (a1585 & b_inv1585) | (a1585 & c1585) | (b_inv1585 & c1585);
  wire s1586, sub1586, and1586, or1586;
  wire b_inv1586;
  assign b_inv1586 = ~b1586;
  assign s1586  = a1586 ^ b1586 ^ c1586;
  assign sub1586 = a1586 ^ b_inv1586 ^ c1586;
  assign and1586 = a1586 & b1586;
  assign or1586  = a1586 | b1586;
  assign c1587 = (a1586 & b1586) | (a1586 & c1586) | (b1586 & c1586);
  wire c_sub1587;
  assign c_sub1587 = (a1586 & b_inv1586) | (a1586 & c1586) | (b_inv1586 & c1586);
  wire s1587, sub1587, and1587, or1587;
  wire b_inv1587;
  assign b_inv1587 = ~b1587;
  assign s1587  = a1587 ^ b1587 ^ c1587;
  assign sub1587 = a1587 ^ b_inv1587 ^ c1587;
  assign and1587 = a1587 & b1587;
  assign or1587  = a1587 | b1587;
  assign c1588 = (a1587 & b1587) | (a1587 & c1587) | (b1587 & c1587);
  wire c_sub1588;
  assign c_sub1588 = (a1587 & b_inv1587) | (a1587 & c1587) | (b_inv1587 & c1587);
  wire s1588, sub1588, and1588, or1588;
  wire b_inv1588;
  assign b_inv1588 = ~b1588;
  assign s1588  = a1588 ^ b1588 ^ c1588;
  assign sub1588 = a1588 ^ b_inv1588 ^ c1588;
  assign and1588 = a1588 & b1588;
  assign or1588  = a1588 | b1588;
  assign c1589 = (a1588 & b1588) | (a1588 & c1588) | (b1588 & c1588);
  wire c_sub1589;
  assign c_sub1589 = (a1588 & b_inv1588) | (a1588 & c1588) | (b_inv1588 & c1588);
  wire s1589, sub1589, and1589, or1589;
  wire b_inv1589;
  assign b_inv1589 = ~b1589;
  assign s1589  = a1589 ^ b1589 ^ c1589;
  assign sub1589 = a1589 ^ b_inv1589 ^ c1589;
  assign and1589 = a1589 & b1589;
  assign or1589  = a1589 | b1589;
  assign c1590 = (a1589 & b1589) | (a1589 & c1589) | (b1589 & c1589);
  wire c_sub1590;
  assign c_sub1590 = (a1589 & b_inv1589) | (a1589 & c1589) | (b_inv1589 & c1589);
  wire s1590, sub1590, and1590, or1590;
  wire b_inv1590;
  assign b_inv1590 = ~b1590;
  assign s1590  = a1590 ^ b1590 ^ c1590;
  assign sub1590 = a1590 ^ b_inv1590 ^ c1590;
  assign and1590 = a1590 & b1590;
  assign or1590  = a1590 | b1590;
  assign c1591 = (a1590 & b1590) | (a1590 & c1590) | (b1590 & c1590);
  wire c_sub1591;
  assign c_sub1591 = (a1590 & b_inv1590) | (a1590 & c1590) | (b_inv1590 & c1590);
  wire s1591, sub1591, and1591, or1591;
  wire b_inv1591;
  assign b_inv1591 = ~b1591;
  assign s1591  = a1591 ^ b1591 ^ c1591;
  assign sub1591 = a1591 ^ b_inv1591 ^ c1591;
  assign and1591 = a1591 & b1591;
  assign or1591  = a1591 | b1591;
  assign c1592 = (a1591 & b1591) | (a1591 & c1591) | (b1591 & c1591);
  wire c_sub1592;
  assign c_sub1592 = (a1591 & b_inv1591) | (a1591 & c1591) | (b_inv1591 & c1591);
  wire s1592, sub1592, and1592, or1592;
  wire b_inv1592;
  assign b_inv1592 = ~b1592;
  assign s1592  = a1592 ^ b1592 ^ c1592;
  assign sub1592 = a1592 ^ b_inv1592 ^ c1592;
  assign and1592 = a1592 & b1592;
  assign or1592  = a1592 | b1592;
  assign c1593 = (a1592 & b1592) | (a1592 & c1592) | (b1592 & c1592);
  wire c_sub1593;
  assign c_sub1593 = (a1592 & b_inv1592) | (a1592 & c1592) | (b_inv1592 & c1592);
  wire s1593, sub1593, and1593, or1593;
  wire b_inv1593;
  assign b_inv1593 = ~b1593;
  assign s1593  = a1593 ^ b1593 ^ c1593;
  assign sub1593 = a1593 ^ b_inv1593 ^ c1593;
  assign and1593 = a1593 & b1593;
  assign or1593  = a1593 | b1593;
  assign c1594 = (a1593 & b1593) | (a1593 & c1593) | (b1593 & c1593);
  wire c_sub1594;
  assign c_sub1594 = (a1593 & b_inv1593) | (a1593 & c1593) | (b_inv1593 & c1593);
  wire s1594, sub1594, and1594, or1594;
  wire b_inv1594;
  assign b_inv1594 = ~b1594;
  assign s1594  = a1594 ^ b1594 ^ c1594;
  assign sub1594 = a1594 ^ b_inv1594 ^ c1594;
  assign and1594 = a1594 & b1594;
  assign or1594  = a1594 | b1594;
  assign c1595 = (a1594 & b1594) | (a1594 & c1594) | (b1594 & c1594);
  wire c_sub1595;
  assign c_sub1595 = (a1594 & b_inv1594) | (a1594 & c1594) | (b_inv1594 & c1594);
  wire s1595, sub1595, and1595, or1595;
  wire b_inv1595;
  assign b_inv1595 = ~b1595;
  assign s1595  = a1595 ^ b1595 ^ c1595;
  assign sub1595 = a1595 ^ b_inv1595 ^ c1595;
  assign and1595 = a1595 & b1595;
  assign or1595  = a1595 | b1595;
  assign c1596 = (a1595 & b1595) | (a1595 & c1595) | (b1595 & c1595);
  wire c_sub1596;
  assign c_sub1596 = (a1595 & b_inv1595) | (a1595 & c1595) | (b_inv1595 & c1595);
  wire s1596, sub1596, and1596, or1596;
  wire b_inv1596;
  assign b_inv1596 = ~b1596;
  assign s1596  = a1596 ^ b1596 ^ c1596;
  assign sub1596 = a1596 ^ b_inv1596 ^ c1596;
  assign and1596 = a1596 & b1596;
  assign or1596  = a1596 | b1596;
  assign c1597 = (a1596 & b1596) | (a1596 & c1596) | (b1596 & c1596);
  wire c_sub1597;
  assign c_sub1597 = (a1596 & b_inv1596) | (a1596 & c1596) | (b_inv1596 & c1596);
  wire s1597, sub1597, and1597, or1597;
  wire b_inv1597;
  assign b_inv1597 = ~b1597;
  assign s1597  = a1597 ^ b1597 ^ c1597;
  assign sub1597 = a1597 ^ b_inv1597 ^ c1597;
  assign and1597 = a1597 & b1597;
  assign or1597  = a1597 | b1597;
  assign c1598 = (a1597 & b1597) | (a1597 & c1597) | (b1597 & c1597);
  wire c_sub1598;
  assign c_sub1598 = (a1597 & b_inv1597) | (a1597 & c1597) | (b_inv1597 & c1597);
  wire s1598, sub1598, and1598, or1598;
  wire b_inv1598;
  assign b_inv1598 = ~b1598;
  assign s1598  = a1598 ^ b1598 ^ c1598;
  assign sub1598 = a1598 ^ b_inv1598 ^ c1598;
  assign and1598 = a1598 & b1598;
  assign or1598  = a1598 | b1598;
  assign c1599 = (a1598 & b1598) | (a1598 & c1598) | (b1598 & c1598);
  wire c_sub1599;
  assign c_sub1599 = (a1598 & b_inv1598) | (a1598 & c1598) | (b_inv1598 & c1598);
  wire s1599, sub1599, and1599, or1599;
  wire b_inv1599;
  assign b_inv1599 = ~b1599;
  assign s1599  = a1599 ^ b1599 ^ c1599;
  assign sub1599 = a1599 ^ b_inv1599 ^ c1599;
  assign and1599 = a1599 & b1599;
  assign or1599  = a1599 | b1599;
  assign c1600 = (a1599 & b1599) | (a1599 & c1599) | (b1599 & c1599);
  wire c_sub1600;
  assign c_sub1600 = (a1599 & b_inv1599) | (a1599 & c1599) | (b_inv1599 & c1599);
  wire s1600, sub1600, and1600, or1600;
  wire b_inv1600;
  assign b_inv1600 = ~b1600;
  assign s1600  = a1600 ^ b1600 ^ c1600;
  assign sub1600 = a1600 ^ b_inv1600 ^ c1600;
  assign and1600 = a1600 & b1600;
  assign or1600  = a1600 | b1600;
  assign c1601 = (a1600 & b1600) | (a1600 & c1600) | (b1600 & c1600);
  wire c_sub1601;
  assign c_sub1601 = (a1600 & b_inv1600) | (a1600 & c1600) | (b_inv1600 & c1600);
  wire s1601, sub1601, and1601, or1601;
  wire b_inv1601;
  assign b_inv1601 = ~b1601;
  assign s1601  = a1601 ^ b1601 ^ c1601;
  assign sub1601 = a1601 ^ b_inv1601 ^ c1601;
  assign and1601 = a1601 & b1601;
  assign or1601  = a1601 | b1601;
  assign c1602 = (a1601 & b1601) | (a1601 & c1601) | (b1601 & c1601);
  wire c_sub1602;
  assign c_sub1602 = (a1601 & b_inv1601) | (a1601 & c1601) | (b_inv1601 & c1601);
  wire s1602, sub1602, and1602, or1602;
  wire b_inv1602;
  assign b_inv1602 = ~b1602;
  assign s1602  = a1602 ^ b1602 ^ c1602;
  assign sub1602 = a1602 ^ b_inv1602 ^ c1602;
  assign and1602 = a1602 & b1602;
  assign or1602  = a1602 | b1602;
  assign c1603 = (a1602 & b1602) | (a1602 & c1602) | (b1602 & c1602);
  wire c_sub1603;
  assign c_sub1603 = (a1602 & b_inv1602) | (a1602 & c1602) | (b_inv1602 & c1602);
  wire s1603, sub1603, and1603, or1603;
  wire b_inv1603;
  assign b_inv1603 = ~b1603;
  assign s1603  = a1603 ^ b1603 ^ c1603;
  assign sub1603 = a1603 ^ b_inv1603 ^ c1603;
  assign and1603 = a1603 & b1603;
  assign or1603  = a1603 | b1603;
  assign c1604 = (a1603 & b1603) | (a1603 & c1603) | (b1603 & c1603);
  wire c_sub1604;
  assign c_sub1604 = (a1603 & b_inv1603) | (a1603 & c1603) | (b_inv1603 & c1603);
  wire s1604, sub1604, and1604, or1604;
  wire b_inv1604;
  assign b_inv1604 = ~b1604;
  assign s1604  = a1604 ^ b1604 ^ c1604;
  assign sub1604 = a1604 ^ b_inv1604 ^ c1604;
  assign and1604 = a1604 & b1604;
  assign or1604  = a1604 | b1604;
  assign c1605 = (a1604 & b1604) | (a1604 & c1604) | (b1604 & c1604);
  wire c_sub1605;
  assign c_sub1605 = (a1604 & b_inv1604) | (a1604 & c1604) | (b_inv1604 & c1604);
  wire s1605, sub1605, and1605, or1605;
  wire b_inv1605;
  assign b_inv1605 = ~b1605;
  assign s1605  = a1605 ^ b1605 ^ c1605;
  assign sub1605 = a1605 ^ b_inv1605 ^ c1605;
  assign and1605 = a1605 & b1605;
  assign or1605  = a1605 | b1605;
  assign c1606 = (a1605 & b1605) | (a1605 & c1605) | (b1605 & c1605);
  wire c_sub1606;
  assign c_sub1606 = (a1605 & b_inv1605) | (a1605 & c1605) | (b_inv1605 & c1605);
  wire s1606, sub1606, and1606, or1606;
  wire b_inv1606;
  assign b_inv1606 = ~b1606;
  assign s1606  = a1606 ^ b1606 ^ c1606;
  assign sub1606 = a1606 ^ b_inv1606 ^ c1606;
  assign and1606 = a1606 & b1606;
  assign or1606  = a1606 | b1606;
  assign c1607 = (a1606 & b1606) | (a1606 & c1606) | (b1606 & c1606);
  wire c_sub1607;
  assign c_sub1607 = (a1606 & b_inv1606) | (a1606 & c1606) | (b_inv1606 & c1606);
  wire s1607, sub1607, and1607, or1607;
  wire b_inv1607;
  assign b_inv1607 = ~b1607;
  assign s1607  = a1607 ^ b1607 ^ c1607;
  assign sub1607 = a1607 ^ b_inv1607 ^ c1607;
  assign and1607 = a1607 & b1607;
  assign or1607  = a1607 | b1607;
  assign c1608 = (a1607 & b1607) | (a1607 & c1607) | (b1607 & c1607);
  wire c_sub1608;
  assign c_sub1608 = (a1607 & b_inv1607) | (a1607 & c1607) | (b_inv1607 & c1607);
  wire s1608, sub1608, and1608, or1608;
  wire b_inv1608;
  assign b_inv1608 = ~b1608;
  assign s1608  = a1608 ^ b1608 ^ c1608;
  assign sub1608 = a1608 ^ b_inv1608 ^ c1608;
  assign and1608 = a1608 & b1608;
  assign or1608  = a1608 | b1608;
  assign c1609 = (a1608 & b1608) | (a1608 & c1608) | (b1608 & c1608);
  wire c_sub1609;
  assign c_sub1609 = (a1608 & b_inv1608) | (a1608 & c1608) | (b_inv1608 & c1608);
  wire s1609, sub1609, and1609, or1609;
  wire b_inv1609;
  assign b_inv1609 = ~b1609;
  assign s1609  = a1609 ^ b1609 ^ c1609;
  assign sub1609 = a1609 ^ b_inv1609 ^ c1609;
  assign and1609 = a1609 & b1609;
  assign or1609  = a1609 | b1609;
  assign c1610 = (a1609 & b1609) | (a1609 & c1609) | (b1609 & c1609);
  wire c_sub1610;
  assign c_sub1610 = (a1609 & b_inv1609) | (a1609 & c1609) | (b_inv1609 & c1609);
  wire s1610, sub1610, and1610, or1610;
  wire b_inv1610;
  assign b_inv1610 = ~b1610;
  assign s1610  = a1610 ^ b1610 ^ c1610;
  assign sub1610 = a1610 ^ b_inv1610 ^ c1610;
  assign and1610 = a1610 & b1610;
  assign or1610  = a1610 | b1610;
  assign c1611 = (a1610 & b1610) | (a1610 & c1610) | (b1610 & c1610);
  wire c_sub1611;
  assign c_sub1611 = (a1610 & b_inv1610) | (a1610 & c1610) | (b_inv1610 & c1610);
  wire s1611, sub1611, and1611, or1611;
  wire b_inv1611;
  assign b_inv1611 = ~b1611;
  assign s1611  = a1611 ^ b1611 ^ c1611;
  assign sub1611 = a1611 ^ b_inv1611 ^ c1611;
  assign and1611 = a1611 & b1611;
  assign or1611  = a1611 | b1611;
  assign c1612 = (a1611 & b1611) | (a1611 & c1611) | (b1611 & c1611);
  wire c_sub1612;
  assign c_sub1612 = (a1611 & b_inv1611) | (a1611 & c1611) | (b_inv1611 & c1611);
  wire s1612, sub1612, and1612, or1612;
  wire b_inv1612;
  assign b_inv1612 = ~b1612;
  assign s1612  = a1612 ^ b1612 ^ c1612;
  assign sub1612 = a1612 ^ b_inv1612 ^ c1612;
  assign and1612 = a1612 & b1612;
  assign or1612  = a1612 | b1612;
  assign c1613 = (a1612 & b1612) | (a1612 & c1612) | (b1612 & c1612);
  wire c_sub1613;
  assign c_sub1613 = (a1612 & b_inv1612) | (a1612 & c1612) | (b_inv1612 & c1612);
  wire s1613, sub1613, and1613, or1613;
  wire b_inv1613;
  assign b_inv1613 = ~b1613;
  assign s1613  = a1613 ^ b1613 ^ c1613;
  assign sub1613 = a1613 ^ b_inv1613 ^ c1613;
  assign and1613 = a1613 & b1613;
  assign or1613  = a1613 | b1613;
  assign c1614 = (a1613 & b1613) | (a1613 & c1613) | (b1613 & c1613);
  wire c_sub1614;
  assign c_sub1614 = (a1613 & b_inv1613) | (a1613 & c1613) | (b_inv1613 & c1613);
  wire s1614, sub1614, and1614, or1614;
  wire b_inv1614;
  assign b_inv1614 = ~b1614;
  assign s1614  = a1614 ^ b1614 ^ c1614;
  assign sub1614 = a1614 ^ b_inv1614 ^ c1614;
  assign and1614 = a1614 & b1614;
  assign or1614  = a1614 | b1614;
  assign c1615 = (a1614 & b1614) | (a1614 & c1614) | (b1614 & c1614);
  wire c_sub1615;
  assign c_sub1615 = (a1614 & b_inv1614) | (a1614 & c1614) | (b_inv1614 & c1614);
  wire s1615, sub1615, and1615, or1615;
  wire b_inv1615;
  assign b_inv1615 = ~b1615;
  assign s1615  = a1615 ^ b1615 ^ c1615;
  assign sub1615 = a1615 ^ b_inv1615 ^ c1615;
  assign and1615 = a1615 & b1615;
  assign or1615  = a1615 | b1615;
  assign c1616 = (a1615 & b1615) | (a1615 & c1615) | (b1615 & c1615);
  wire c_sub1616;
  assign c_sub1616 = (a1615 & b_inv1615) | (a1615 & c1615) | (b_inv1615 & c1615);
  wire s1616, sub1616, and1616, or1616;
  wire b_inv1616;
  assign b_inv1616 = ~b1616;
  assign s1616  = a1616 ^ b1616 ^ c1616;
  assign sub1616 = a1616 ^ b_inv1616 ^ c1616;
  assign and1616 = a1616 & b1616;
  assign or1616  = a1616 | b1616;
  assign c1617 = (a1616 & b1616) | (a1616 & c1616) | (b1616 & c1616);
  wire c_sub1617;
  assign c_sub1617 = (a1616 & b_inv1616) | (a1616 & c1616) | (b_inv1616 & c1616);
  wire s1617, sub1617, and1617, or1617;
  wire b_inv1617;
  assign b_inv1617 = ~b1617;
  assign s1617  = a1617 ^ b1617 ^ c1617;
  assign sub1617 = a1617 ^ b_inv1617 ^ c1617;
  assign and1617 = a1617 & b1617;
  assign or1617  = a1617 | b1617;
  assign c1618 = (a1617 & b1617) | (a1617 & c1617) | (b1617 & c1617);
  wire c_sub1618;
  assign c_sub1618 = (a1617 & b_inv1617) | (a1617 & c1617) | (b_inv1617 & c1617);
  wire s1618, sub1618, and1618, or1618;
  wire b_inv1618;
  assign b_inv1618 = ~b1618;
  assign s1618  = a1618 ^ b1618 ^ c1618;
  assign sub1618 = a1618 ^ b_inv1618 ^ c1618;
  assign and1618 = a1618 & b1618;
  assign or1618  = a1618 | b1618;
  assign c1619 = (a1618 & b1618) | (a1618 & c1618) | (b1618 & c1618);
  wire c_sub1619;
  assign c_sub1619 = (a1618 & b_inv1618) | (a1618 & c1618) | (b_inv1618 & c1618);
  wire s1619, sub1619, and1619, or1619;
  wire b_inv1619;
  assign b_inv1619 = ~b1619;
  assign s1619  = a1619 ^ b1619 ^ c1619;
  assign sub1619 = a1619 ^ b_inv1619 ^ c1619;
  assign and1619 = a1619 & b1619;
  assign or1619  = a1619 | b1619;
  assign c1620 = (a1619 & b1619) | (a1619 & c1619) | (b1619 & c1619);
  wire c_sub1620;
  assign c_sub1620 = (a1619 & b_inv1619) | (a1619 & c1619) | (b_inv1619 & c1619);
  wire s1620, sub1620, and1620, or1620;
  wire b_inv1620;
  assign b_inv1620 = ~b1620;
  assign s1620  = a1620 ^ b1620 ^ c1620;
  assign sub1620 = a1620 ^ b_inv1620 ^ c1620;
  assign and1620 = a1620 & b1620;
  assign or1620  = a1620 | b1620;
  assign c1621 = (a1620 & b1620) | (a1620 & c1620) | (b1620 & c1620);
  wire c_sub1621;
  assign c_sub1621 = (a1620 & b_inv1620) | (a1620 & c1620) | (b_inv1620 & c1620);
  wire s1621, sub1621, and1621, or1621;
  wire b_inv1621;
  assign b_inv1621 = ~b1621;
  assign s1621  = a1621 ^ b1621 ^ c1621;
  assign sub1621 = a1621 ^ b_inv1621 ^ c1621;
  assign and1621 = a1621 & b1621;
  assign or1621  = a1621 | b1621;
  assign c1622 = (a1621 & b1621) | (a1621 & c1621) | (b1621 & c1621);
  wire c_sub1622;
  assign c_sub1622 = (a1621 & b_inv1621) | (a1621 & c1621) | (b_inv1621 & c1621);
  wire s1622, sub1622, and1622, or1622;
  wire b_inv1622;
  assign b_inv1622 = ~b1622;
  assign s1622  = a1622 ^ b1622 ^ c1622;
  assign sub1622 = a1622 ^ b_inv1622 ^ c1622;
  assign and1622 = a1622 & b1622;
  assign or1622  = a1622 | b1622;
  assign c1623 = (a1622 & b1622) | (a1622 & c1622) | (b1622 & c1622);
  wire c_sub1623;
  assign c_sub1623 = (a1622 & b_inv1622) | (a1622 & c1622) | (b_inv1622 & c1622);
  wire s1623, sub1623, and1623, or1623;
  wire b_inv1623;
  assign b_inv1623 = ~b1623;
  assign s1623  = a1623 ^ b1623 ^ c1623;
  assign sub1623 = a1623 ^ b_inv1623 ^ c1623;
  assign and1623 = a1623 & b1623;
  assign or1623  = a1623 | b1623;
  assign c1624 = (a1623 & b1623) | (a1623 & c1623) | (b1623 & c1623);
  wire c_sub1624;
  assign c_sub1624 = (a1623 & b_inv1623) | (a1623 & c1623) | (b_inv1623 & c1623);
  wire s1624, sub1624, and1624, or1624;
  wire b_inv1624;
  assign b_inv1624 = ~b1624;
  assign s1624  = a1624 ^ b1624 ^ c1624;
  assign sub1624 = a1624 ^ b_inv1624 ^ c1624;
  assign and1624 = a1624 & b1624;
  assign or1624  = a1624 | b1624;
  assign c1625 = (a1624 & b1624) | (a1624 & c1624) | (b1624 & c1624);
  wire c_sub1625;
  assign c_sub1625 = (a1624 & b_inv1624) | (a1624 & c1624) | (b_inv1624 & c1624);
  wire s1625, sub1625, and1625, or1625;
  wire b_inv1625;
  assign b_inv1625 = ~b1625;
  assign s1625  = a1625 ^ b1625 ^ c1625;
  assign sub1625 = a1625 ^ b_inv1625 ^ c1625;
  assign and1625 = a1625 & b1625;
  assign or1625  = a1625 | b1625;
  assign c1626 = (a1625 & b1625) | (a1625 & c1625) | (b1625 & c1625);
  wire c_sub1626;
  assign c_sub1626 = (a1625 & b_inv1625) | (a1625 & c1625) | (b_inv1625 & c1625);
  wire s1626, sub1626, and1626, or1626;
  wire b_inv1626;
  assign b_inv1626 = ~b1626;
  assign s1626  = a1626 ^ b1626 ^ c1626;
  assign sub1626 = a1626 ^ b_inv1626 ^ c1626;
  assign and1626 = a1626 & b1626;
  assign or1626  = a1626 | b1626;
  assign c1627 = (a1626 & b1626) | (a1626 & c1626) | (b1626 & c1626);
  wire c_sub1627;
  assign c_sub1627 = (a1626 & b_inv1626) | (a1626 & c1626) | (b_inv1626 & c1626);
  wire s1627, sub1627, and1627, or1627;
  wire b_inv1627;
  assign b_inv1627 = ~b1627;
  assign s1627  = a1627 ^ b1627 ^ c1627;
  assign sub1627 = a1627 ^ b_inv1627 ^ c1627;
  assign and1627 = a1627 & b1627;
  assign or1627  = a1627 | b1627;
  assign c1628 = (a1627 & b1627) | (a1627 & c1627) | (b1627 & c1627);
  wire c_sub1628;
  assign c_sub1628 = (a1627 & b_inv1627) | (a1627 & c1627) | (b_inv1627 & c1627);
  wire s1628, sub1628, and1628, or1628;
  wire b_inv1628;
  assign b_inv1628 = ~b1628;
  assign s1628  = a1628 ^ b1628 ^ c1628;
  assign sub1628 = a1628 ^ b_inv1628 ^ c1628;
  assign and1628 = a1628 & b1628;
  assign or1628  = a1628 | b1628;
  assign c1629 = (a1628 & b1628) | (a1628 & c1628) | (b1628 & c1628);
  wire c_sub1629;
  assign c_sub1629 = (a1628 & b_inv1628) | (a1628 & c1628) | (b_inv1628 & c1628);
  wire s1629, sub1629, and1629, or1629;
  wire b_inv1629;
  assign b_inv1629 = ~b1629;
  assign s1629  = a1629 ^ b1629 ^ c1629;
  assign sub1629 = a1629 ^ b_inv1629 ^ c1629;
  assign and1629 = a1629 & b1629;
  assign or1629  = a1629 | b1629;
  assign c1630 = (a1629 & b1629) | (a1629 & c1629) | (b1629 & c1629);
  wire c_sub1630;
  assign c_sub1630 = (a1629 & b_inv1629) | (a1629 & c1629) | (b_inv1629 & c1629);
  wire s1630, sub1630, and1630, or1630;
  wire b_inv1630;
  assign b_inv1630 = ~b1630;
  assign s1630  = a1630 ^ b1630 ^ c1630;
  assign sub1630 = a1630 ^ b_inv1630 ^ c1630;
  assign and1630 = a1630 & b1630;
  assign or1630  = a1630 | b1630;
  assign c1631 = (a1630 & b1630) | (a1630 & c1630) | (b1630 & c1630);
  wire c_sub1631;
  assign c_sub1631 = (a1630 & b_inv1630) | (a1630 & c1630) | (b_inv1630 & c1630);
  wire s1631, sub1631, and1631, or1631;
  wire b_inv1631;
  assign b_inv1631 = ~b1631;
  assign s1631  = a1631 ^ b1631 ^ c1631;
  assign sub1631 = a1631 ^ b_inv1631 ^ c1631;
  assign and1631 = a1631 & b1631;
  assign or1631  = a1631 | b1631;
  assign c1632 = (a1631 & b1631) | (a1631 & c1631) | (b1631 & c1631);
  wire c_sub1632;
  assign c_sub1632 = (a1631 & b_inv1631) | (a1631 & c1631) | (b_inv1631 & c1631);
  wire s1632, sub1632, and1632, or1632;
  wire b_inv1632;
  assign b_inv1632 = ~b1632;
  assign s1632  = a1632 ^ b1632 ^ c1632;
  assign sub1632 = a1632 ^ b_inv1632 ^ c1632;
  assign and1632 = a1632 & b1632;
  assign or1632  = a1632 | b1632;
  assign c1633 = (a1632 & b1632) | (a1632 & c1632) | (b1632 & c1632);
  wire c_sub1633;
  assign c_sub1633 = (a1632 & b_inv1632) | (a1632 & c1632) | (b_inv1632 & c1632);
  wire s1633, sub1633, and1633, or1633;
  wire b_inv1633;
  assign b_inv1633 = ~b1633;
  assign s1633  = a1633 ^ b1633 ^ c1633;
  assign sub1633 = a1633 ^ b_inv1633 ^ c1633;
  assign and1633 = a1633 & b1633;
  assign or1633  = a1633 | b1633;
  assign c1634 = (a1633 & b1633) | (a1633 & c1633) | (b1633 & c1633);
  wire c_sub1634;
  assign c_sub1634 = (a1633 & b_inv1633) | (a1633 & c1633) | (b_inv1633 & c1633);
  wire s1634, sub1634, and1634, or1634;
  wire b_inv1634;
  assign b_inv1634 = ~b1634;
  assign s1634  = a1634 ^ b1634 ^ c1634;
  assign sub1634 = a1634 ^ b_inv1634 ^ c1634;
  assign and1634 = a1634 & b1634;
  assign or1634  = a1634 | b1634;
  assign c1635 = (a1634 & b1634) | (a1634 & c1634) | (b1634 & c1634);
  wire c_sub1635;
  assign c_sub1635 = (a1634 & b_inv1634) | (a1634 & c1634) | (b_inv1634 & c1634);
  wire s1635, sub1635, and1635, or1635;
  wire b_inv1635;
  assign b_inv1635 = ~b1635;
  assign s1635  = a1635 ^ b1635 ^ c1635;
  assign sub1635 = a1635 ^ b_inv1635 ^ c1635;
  assign and1635 = a1635 & b1635;
  assign or1635  = a1635 | b1635;
  assign c1636 = (a1635 & b1635) | (a1635 & c1635) | (b1635 & c1635);
  wire c_sub1636;
  assign c_sub1636 = (a1635 & b_inv1635) | (a1635 & c1635) | (b_inv1635 & c1635);
  wire s1636, sub1636, and1636, or1636;
  wire b_inv1636;
  assign b_inv1636 = ~b1636;
  assign s1636  = a1636 ^ b1636 ^ c1636;
  assign sub1636 = a1636 ^ b_inv1636 ^ c1636;
  assign and1636 = a1636 & b1636;
  assign or1636  = a1636 | b1636;
  assign c1637 = (a1636 & b1636) | (a1636 & c1636) | (b1636 & c1636);
  wire c_sub1637;
  assign c_sub1637 = (a1636 & b_inv1636) | (a1636 & c1636) | (b_inv1636 & c1636);
  wire s1637, sub1637, and1637, or1637;
  wire b_inv1637;
  assign b_inv1637 = ~b1637;
  assign s1637  = a1637 ^ b1637 ^ c1637;
  assign sub1637 = a1637 ^ b_inv1637 ^ c1637;
  assign and1637 = a1637 & b1637;
  assign or1637  = a1637 | b1637;
  assign c1638 = (a1637 & b1637) | (a1637 & c1637) | (b1637 & c1637);
  wire c_sub1638;
  assign c_sub1638 = (a1637 & b_inv1637) | (a1637 & c1637) | (b_inv1637 & c1637);
  wire s1638, sub1638, and1638, or1638;
  wire b_inv1638;
  assign b_inv1638 = ~b1638;
  assign s1638  = a1638 ^ b1638 ^ c1638;
  assign sub1638 = a1638 ^ b_inv1638 ^ c1638;
  assign and1638 = a1638 & b1638;
  assign or1638  = a1638 | b1638;
  assign c1639 = (a1638 & b1638) | (a1638 & c1638) | (b1638 & c1638);
  wire c_sub1639;
  assign c_sub1639 = (a1638 & b_inv1638) | (a1638 & c1638) | (b_inv1638 & c1638);
  wire s1639, sub1639, and1639, or1639;
  wire b_inv1639;
  assign b_inv1639 = ~b1639;
  assign s1639  = a1639 ^ b1639 ^ c1639;
  assign sub1639 = a1639 ^ b_inv1639 ^ c1639;
  assign and1639 = a1639 & b1639;
  assign or1639  = a1639 | b1639;
  assign c1640 = (a1639 & b1639) | (a1639 & c1639) | (b1639 & c1639);
  wire c_sub1640;
  assign c_sub1640 = (a1639 & b_inv1639) | (a1639 & c1639) | (b_inv1639 & c1639);
  wire s1640, sub1640, and1640, or1640;
  wire b_inv1640;
  assign b_inv1640 = ~b1640;
  assign s1640  = a1640 ^ b1640 ^ c1640;
  assign sub1640 = a1640 ^ b_inv1640 ^ c1640;
  assign and1640 = a1640 & b1640;
  assign or1640  = a1640 | b1640;
  assign c1641 = (a1640 & b1640) | (a1640 & c1640) | (b1640 & c1640);
  wire c_sub1641;
  assign c_sub1641 = (a1640 & b_inv1640) | (a1640 & c1640) | (b_inv1640 & c1640);
  wire s1641, sub1641, and1641, or1641;
  wire b_inv1641;
  assign b_inv1641 = ~b1641;
  assign s1641  = a1641 ^ b1641 ^ c1641;
  assign sub1641 = a1641 ^ b_inv1641 ^ c1641;
  assign and1641 = a1641 & b1641;
  assign or1641  = a1641 | b1641;
  assign c1642 = (a1641 & b1641) | (a1641 & c1641) | (b1641 & c1641);
  wire c_sub1642;
  assign c_sub1642 = (a1641 & b_inv1641) | (a1641 & c1641) | (b_inv1641 & c1641);
  wire s1642, sub1642, and1642, or1642;
  wire b_inv1642;
  assign b_inv1642 = ~b1642;
  assign s1642  = a1642 ^ b1642 ^ c1642;
  assign sub1642 = a1642 ^ b_inv1642 ^ c1642;
  assign and1642 = a1642 & b1642;
  assign or1642  = a1642 | b1642;
  assign c1643 = (a1642 & b1642) | (a1642 & c1642) | (b1642 & c1642);
  wire c_sub1643;
  assign c_sub1643 = (a1642 & b_inv1642) | (a1642 & c1642) | (b_inv1642 & c1642);
  wire s1643, sub1643, and1643, or1643;
  wire b_inv1643;
  assign b_inv1643 = ~b1643;
  assign s1643  = a1643 ^ b1643 ^ c1643;
  assign sub1643 = a1643 ^ b_inv1643 ^ c1643;
  assign and1643 = a1643 & b1643;
  assign or1643  = a1643 | b1643;
  assign c1644 = (a1643 & b1643) | (a1643 & c1643) | (b1643 & c1643);
  wire c_sub1644;
  assign c_sub1644 = (a1643 & b_inv1643) | (a1643 & c1643) | (b_inv1643 & c1643);
  wire s1644, sub1644, and1644, or1644;
  wire b_inv1644;
  assign b_inv1644 = ~b1644;
  assign s1644  = a1644 ^ b1644 ^ c1644;
  assign sub1644 = a1644 ^ b_inv1644 ^ c1644;
  assign and1644 = a1644 & b1644;
  assign or1644  = a1644 | b1644;
  assign c1645 = (a1644 & b1644) | (a1644 & c1644) | (b1644 & c1644);
  wire c_sub1645;
  assign c_sub1645 = (a1644 & b_inv1644) | (a1644 & c1644) | (b_inv1644 & c1644);
  wire s1645, sub1645, and1645, or1645;
  wire b_inv1645;
  assign b_inv1645 = ~b1645;
  assign s1645  = a1645 ^ b1645 ^ c1645;
  assign sub1645 = a1645 ^ b_inv1645 ^ c1645;
  assign and1645 = a1645 & b1645;
  assign or1645  = a1645 | b1645;
  assign c1646 = (a1645 & b1645) | (a1645 & c1645) | (b1645 & c1645);
  wire c_sub1646;
  assign c_sub1646 = (a1645 & b_inv1645) | (a1645 & c1645) | (b_inv1645 & c1645);
  wire s1646, sub1646, and1646, or1646;
  wire b_inv1646;
  assign b_inv1646 = ~b1646;
  assign s1646  = a1646 ^ b1646 ^ c1646;
  assign sub1646 = a1646 ^ b_inv1646 ^ c1646;
  assign and1646 = a1646 & b1646;
  assign or1646  = a1646 | b1646;
  assign c1647 = (a1646 & b1646) | (a1646 & c1646) | (b1646 & c1646);
  wire c_sub1647;
  assign c_sub1647 = (a1646 & b_inv1646) | (a1646 & c1646) | (b_inv1646 & c1646);
  wire s1647, sub1647, and1647, or1647;
  wire b_inv1647;
  assign b_inv1647 = ~b1647;
  assign s1647  = a1647 ^ b1647 ^ c1647;
  assign sub1647 = a1647 ^ b_inv1647 ^ c1647;
  assign and1647 = a1647 & b1647;
  assign or1647  = a1647 | b1647;
  assign c1648 = (a1647 & b1647) | (a1647 & c1647) | (b1647 & c1647);
  wire c_sub1648;
  assign c_sub1648 = (a1647 & b_inv1647) | (a1647 & c1647) | (b_inv1647 & c1647);
  wire s1648, sub1648, and1648, or1648;
  wire b_inv1648;
  assign b_inv1648 = ~b1648;
  assign s1648  = a1648 ^ b1648 ^ c1648;
  assign sub1648 = a1648 ^ b_inv1648 ^ c1648;
  assign and1648 = a1648 & b1648;
  assign or1648  = a1648 | b1648;
  assign c1649 = (a1648 & b1648) | (a1648 & c1648) | (b1648 & c1648);
  wire c_sub1649;
  assign c_sub1649 = (a1648 & b_inv1648) | (a1648 & c1648) | (b_inv1648 & c1648);
  wire s1649, sub1649, and1649, or1649;
  wire b_inv1649;
  assign b_inv1649 = ~b1649;
  assign s1649  = a1649 ^ b1649 ^ c1649;
  assign sub1649 = a1649 ^ b_inv1649 ^ c1649;
  assign and1649 = a1649 & b1649;
  assign or1649  = a1649 | b1649;
  assign c1650 = (a1649 & b1649) | (a1649 & c1649) | (b1649 & c1649);
  wire c_sub1650;
  assign c_sub1650 = (a1649 & b_inv1649) | (a1649 & c1649) | (b_inv1649 & c1649);
  wire s1650, sub1650, and1650, or1650;
  wire b_inv1650;
  assign b_inv1650 = ~b1650;
  assign s1650  = a1650 ^ b1650 ^ c1650;
  assign sub1650 = a1650 ^ b_inv1650 ^ c1650;
  assign and1650 = a1650 & b1650;
  assign or1650  = a1650 | b1650;
  assign c1651 = (a1650 & b1650) | (a1650 & c1650) | (b1650 & c1650);
  wire c_sub1651;
  assign c_sub1651 = (a1650 & b_inv1650) | (a1650 & c1650) | (b_inv1650 & c1650);
  wire s1651, sub1651, and1651, or1651;
  wire b_inv1651;
  assign b_inv1651 = ~b1651;
  assign s1651  = a1651 ^ b1651 ^ c1651;
  assign sub1651 = a1651 ^ b_inv1651 ^ c1651;
  assign and1651 = a1651 & b1651;
  assign or1651  = a1651 | b1651;
  assign c1652 = (a1651 & b1651) | (a1651 & c1651) | (b1651 & c1651);
  wire c_sub1652;
  assign c_sub1652 = (a1651 & b_inv1651) | (a1651 & c1651) | (b_inv1651 & c1651);
  wire s1652, sub1652, and1652, or1652;
  wire b_inv1652;
  assign b_inv1652 = ~b1652;
  assign s1652  = a1652 ^ b1652 ^ c1652;
  assign sub1652 = a1652 ^ b_inv1652 ^ c1652;
  assign and1652 = a1652 & b1652;
  assign or1652  = a1652 | b1652;
  assign c1653 = (a1652 & b1652) | (a1652 & c1652) | (b1652 & c1652);
  wire c_sub1653;
  assign c_sub1653 = (a1652 & b_inv1652) | (a1652 & c1652) | (b_inv1652 & c1652);
  wire s1653, sub1653, and1653, or1653;
  wire b_inv1653;
  assign b_inv1653 = ~b1653;
  assign s1653  = a1653 ^ b1653 ^ c1653;
  assign sub1653 = a1653 ^ b_inv1653 ^ c1653;
  assign and1653 = a1653 & b1653;
  assign or1653  = a1653 | b1653;
  assign c1654 = (a1653 & b1653) | (a1653 & c1653) | (b1653 & c1653);
  wire c_sub1654;
  assign c_sub1654 = (a1653 & b_inv1653) | (a1653 & c1653) | (b_inv1653 & c1653);
  wire s1654, sub1654, and1654, or1654;
  wire b_inv1654;
  assign b_inv1654 = ~b1654;
  assign s1654  = a1654 ^ b1654 ^ c1654;
  assign sub1654 = a1654 ^ b_inv1654 ^ c1654;
  assign and1654 = a1654 & b1654;
  assign or1654  = a1654 | b1654;
  assign c1655 = (a1654 & b1654) | (a1654 & c1654) | (b1654 & c1654);
  wire c_sub1655;
  assign c_sub1655 = (a1654 & b_inv1654) | (a1654 & c1654) | (b_inv1654 & c1654);
  wire s1655, sub1655, and1655, or1655;
  wire b_inv1655;
  assign b_inv1655 = ~b1655;
  assign s1655  = a1655 ^ b1655 ^ c1655;
  assign sub1655 = a1655 ^ b_inv1655 ^ c1655;
  assign and1655 = a1655 & b1655;
  assign or1655  = a1655 | b1655;
  assign c1656 = (a1655 & b1655) | (a1655 & c1655) | (b1655 & c1655);
  wire c_sub1656;
  assign c_sub1656 = (a1655 & b_inv1655) | (a1655 & c1655) | (b_inv1655 & c1655);
  wire s1656, sub1656, and1656, or1656;
  wire b_inv1656;
  assign b_inv1656 = ~b1656;
  assign s1656  = a1656 ^ b1656 ^ c1656;
  assign sub1656 = a1656 ^ b_inv1656 ^ c1656;
  assign and1656 = a1656 & b1656;
  assign or1656  = a1656 | b1656;
  assign c1657 = (a1656 & b1656) | (a1656 & c1656) | (b1656 & c1656);
  wire c_sub1657;
  assign c_sub1657 = (a1656 & b_inv1656) | (a1656 & c1656) | (b_inv1656 & c1656);
  wire s1657, sub1657, and1657, or1657;
  wire b_inv1657;
  assign b_inv1657 = ~b1657;
  assign s1657  = a1657 ^ b1657 ^ c1657;
  assign sub1657 = a1657 ^ b_inv1657 ^ c1657;
  assign and1657 = a1657 & b1657;
  assign or1657  = a1657 | b1657;
  assign c1658 = (a1657 & b1657) | (a1657 & c1657) | (b1657 & c1657);
  wire c_sub1658;
  assign c_sub1658 = (a1657 & b_inv1657) | (a1657 & c1657) | (b_inv1657 & c1657);
  wire s1658, sub1658, and1658, or1658;
  wire b_inv1658;
  assign b_inv1658 = ~b1658;
  assign s1658  = a1658 ^ b1658 ^ c1658;
  assign sub1658 = a1658 ^ b_inv1658 ^ c1658;
  assign and1658 = a1658 & b1658;
  assign or1658  = a1658 | b1658;
  assign c1659 = (a1658 & b1658) | (a1658 & c1658) | (b1658 & c1658);
  wire c_sub1659;
  assign c_sub1659 = (a1658 & b_inv1658) | (a1658 & c1658) | (b_inv1658 & c1658);
  wire s1659, sub1659, and1659, or1659;
  wire b_inv1659;
  assign b_inv1659 = ~b1659;
  assign s1659  = a1659 ^ b1659 ^ c1659;
  assign sub1659 = a1659 ^ b_inv1659 ^ c1659;
  assign and1659 = a1659 & b1659;
  assign or1659  = a1659 | b1659;
  assign c1660 = (a1659 & b1659) | (a1659 & c1659) | (b1659 & c1659);
  wire c_sub1660;
  assign c_sub1660 = (a1659 & b_inv1659) | (a1659 & c1659) | (b_inv1659 & c1659);
  wire s1660, sub1660, and1660, or1660;
  wire b_inv1660;
  assign b_inv1660 = ~b1660;
  assign s1660  = a1660 ^ b1660 ^ c1660;
  assign sub1660 = a1660 ^ b_inv1660 ^ c1660;
  assign and1660 = a1660 & b1660;
  assign or1660  = a1660 | b1660;
  assign c1661 = (a1660 & b1660) | (a1660 & c1660) | (b1660 & c1660);
  wire c_sub1661;
  assign c_sub1661 = (a1660 & b_inv1660) | (a1660 & c1660) | (b_inv1660 & c1660);
  wire s1661, sub1661, and1661, or1661;
  wire b_inv1661;
  assign b_inv1661 = ~b1661;
  assign s1661  = a1661 ^ b1661 ^ c1661;
  assign sub1661 = a1661 ^ b_inv1661 ^ c1661;
  assign and1661 = a1661 & b1661;
  assign or1661  = a1661 | b1661;
  assign c1662 = (a1661 & b1661) | (a1661 & c1661) | (b1661 & c1661);
  wire c_sub1662;
  assign c_sub1662 = (a1661 & b_inv1661) | (a1661 & c1661) | (b_inv1661 & c1661);
  wire s1662, sub1662, and1662, or1662;
  wire b_inv1662;
  assign b_inv1662 = ~b1662;
  assign s1662  = a1662 ^ b1662 ^ c1662;
  assign sub1662 = a1662 ^ b_inv1662 ^ c1662;
  assign and1662 = a1662 & b1662;
  assign or1662  = a1662 | b1662;
  assign c1663 = (a1662 & b1662) | (a1662 & c1662) | (b1662 & c1662);
  wire c_sub1663;
  assign c_sub1663 = (a1662 & b_inv1662) | (a1662 & c1662) | (b_inv1662 & c1662);
  wire s1663, sub1663, and1663, or1663;
  wire b_inv1663;
  assign b_inv1663 = ~b1663;
  assign s1663  = a1663 ^ b1663 ^ c1663;
  assign sub1663 = a1663 ^ b_inv1663 ^ c1663;
  assign and1663 = a1663 & b1663;
  assign or1663  = a1663 | b1663;
  assign c1664 = (a1663 & b1663) | (a1663 & c1663) | (b1663 & c1663);
  wire c_sub1664;
  assign c_sub1664 = (a1663 & b_inv1663) | (a1663 & c1663) | (b_inv1663 & c1663);
  wire s1664, sub1664, and1664, or1664;
  wire b_inv1664;
  assign b_inv1664 = ~b1664;
  assign s1664  = a1664 ^ b1664 ^ c1664;
  assign sub1664 = a1664 ^ b_inv1664 ^ c1664;
  assign and1664 = a1664 & b1664;
  assign or1664  = a1664 | b1664;
  assign c1665 = (a1664 & b1664) | (a1664 & c1664) | (b1664 & c1664);
  wire c_sub1665;
  assign c_sub1665 = (a1664 & b_inv1664) | (a1664 & c1664) | (b_inv1664 & c1664);
  wire s1665, sub1665, and1665, or1665;
  wire b_inv1665;
  assign b_inv1665 = ~b1665;
  assign s1665  = a1665 ^ b1665 ^ c1665;
  assign sub1665 = a1665 ^ b_inv1665 ^ c1665;
  assign and1665 = a1665 & b1665;
  assign or1665  = a1665 | b1665;
  assign c1666 = (a1665 & b1665) | (a1665 & c1665) | (b1665 & c1665);
  wire c_sub1666;
  assign c_sub1666 = (a1665 & b_inv1665) | (a1665 & c1665) | (b_inv1665 & c1665);
  wire s1666, sub1666, and1666, or1666;
  wire b_inv1666;
  assign b_inv1666 = ~b1666;
  assign s1666  = a1666 ^ b1666 ^ c1666;
  assign sub1666 = a1666 ^ b_inv1666 ^ c1666;
  assign and1666 = a1666 & b1666;
  assign or1666  = a1666 | b1666;
  assign c1667 = (a1666 & b1666) | (a1666 & c1666) | (b1666 & c1666);
  wire c_sub1667;
  assign c_sub1667 = (a1666 & b_inv1666) | (a1666 & c1666) | (b_inv1666 & c1666);
  wire s1667, sub1667, and1667, or1667;
  wire b_inv1667;
  assign b_inv1667 = ~b1667;
  assign s1667  = a1667 ^ b1667 ^ c1667;
  assign sub1667 = a1667 ^ b_inv1667 ^ c1667;
  assign and1667 = a1667 & b1667;
  assign or1667  = a1667 | b1667;
  assign c1668 = (a1667 & b1667) | (a1667 & c1667) | (b1667 & c1667);
  wire c_sub1668;
  assign c_sub1668 = (a1667 & b_inv1667) | (a1667 & c1667) | (b_inv1667 & c1667);
  wire s1668, sub1668, and1668, or1668;
  wire b_inv1668;
  assign b_inv1668 = ~b1668;
  assign s1668  = a1668 ^ b1668 ^ c1668;
  assign sub1668 = a1668 ^ b_inv1668 ^ c1668;
  assign and1668 = a1668 & b1668;
  assign or1668  = a1668 | b1668;
  assign c1669 = (a1668 & b1668) | (a1668 & c1668) | (b1668 & c1668);
  wire c_sub1669;
  assign c_sub1669 = (a1668 & b_inv1668) | (a1668 & c1668) | (b_inv1668 & c1668);
  wire s1669, sub1669, and1669, or1669;
  wire b_inv1669;
  assign b_inv1669 = ~b1669;
  assign s1669  = a1669 ^ b1669 ^ c1669;
  assign sub1669 = a1669 ^ b_inv1669 ^ c1669;
  assign and1669 = a1669 & b1669;
  assign or1669  = a1669 | b1669;
  assign c1670 = (a1669 & b1669) | (a1669 & c1669) | (b1669 & c1669);
  wire c_sub1670;
  assign c_sub1670 = (a1669 & b_inv1669) | (a1669 & c1669) | (b_inv1669 & c1669);
  wire s1670, sub1670, and1670, or1670;
  wire b_inv1670;
  assign b_inv1670 = ~b1670;
  assign s1670  = a1670 ^ b1670 ^ c1670;
  assign sub1670 = a1670 ^ b_inv1670 ^ c1670;
  assign and1670 = a1670 & b1670;
  assign or1670  = a1670 | b1670;
  assign c1671 = (a1670 & b1670) | (a1670 & c1670) | (b1670 & c1670);
  wire c_sub1671;
  assign c_sub1671 = (a1670 & b_inv1670) | (a1670 & c1670) | (b_inv1670 & c1670);
  wire s1671, sub1671, and1671, or1671;
  wire b_inv1671;
  assign b_inv1671 = ~b1671;
  assign s1671  = a1671 ^ b1671 ^ c1671;
  assign sub1671 = a1671 ^ b_inv1671 ^ c1671;
  assign and1671 = a1671 & b1671;
  assign or1671  = a1671 | b1671;
  assign c1672 = (a1671 & b1671) | (a1671 & c1671) | (b1671 & c1671);
  wire c_sub1672;
  assign c_sub1672 = (a1671 & b_inv1671) | (a1671 & c1671) | (b_inv1671 & c1671);
  wire s1672, sub1672, and1672, or1672;
  wire b_inv1672;
  assign b_inv1672 = ~b1672;
  assign s1672  = a1672 ^ b1672 ^ c1672;
  assign sub1672 = a1672 ^ b_inv1672 ^ c1672;
  assign and1672 = a1672 & b1672;
  assign or1672  = a1672 | b1672;
  assign c1673 = (a1672 & b1672) | (a1672 & c1672) | (b1672 & c1672);
  wire c_sub1673;
  assign c_sub1673 = (a1672 & b_inv1672) | (a1672 & c1672) | (b_inv1672 & c1672);
  wire s1673, sub1673, and1673, or1673;
  wire b_inv1673;
  assign b_inv1673 = ~b1673;
  assign s1673  = a1673 ^ b1673 ^ c1673;
  assign sub1673 = a1673 ^ b_inv1673 ^ c1673;
  assign and1673 = a1673 & b1673;
  assign or1673  = a1673 | b1673;
  assign c1674 = (a1673 & b1673) | (a1673 & c1673) | (b1673 & c1673);
  wire c_sub1674;
  assign c_sub1674 = (a1673 & b_inv1673) | (a1673 & c1673) | (b_inv1673 & c1673);
  wire s1674, sub1674, and1674, or1674;
  wire b_inv1674;
  assign b_inv1674 = ~b1674;
  assign s1674  = a1674 ^ b1674 ^ c1674;
  assign sub1674 = a1674 ^ b_inv1674 ^ c1674;
  assign and1674 = a1674 & b1674;
  assign or1674  = a1674 | b1674;
  assign c1675 = (a1674 & b1674) | (a1674 & c1674) | (b1674 & c1674);
  wire c_sub1675;
  assign c_sub1675 = (a1674 & b_inv1674) | (a1674 & c1674) | (b_inv1674 & c1674);
  wire s1675, sub1675, and1675, or1675;
  wire b_inv1675;
  assign b_inv1675 = ~b1675;
  assign s1675  = a1675 ^ b1675 ^ c1675;
  assign sub1675 = a1675 ^ b_inv1675 ^ c1675;
  assign and1675 = a1675 & b1675;
  assign or1675  = a1675 | b1675;
  assign c1676 = (a1675 & b1675) | (a1675 & c1675) | (b1675 & c1675);
  wire c_sub1676;
  assign c_sub1676 = (a1675 & b_inv1675) | (a1675 & c1675) | (b_inv1675 & c1675);
  wire s1676, sub1676, and1676, or1676;
  wire b_inv1676;
  assign b_inv1676 = ~b1676;
  assign s1676  = a1676 ^ b1676 ^ c1676;
  assign sub1676 = a1676 ^ b_inv1676 ^ c1676;
  assign and1676 = a1676 & b1676;
  assign or1676  = a1676 | b1676;
  assign c1677 = (a1676 & b1676) | (a1676 & c1676) | (b1676 & c1676);
  wire c_sub1677;
  assign c_sub1677 = (a1676 & b_inv1676) | (a1676 & c1676) | (b_inv1676 & c1676);
  wire s1677, sub1677, and1677, or1677;
  wire b_inv1677;
  assign b_inv1677 = ~b1677;
  assign s1677  = a1677 ^ b1677 ^ c1677;
  assign sub1677 = a1677 ^ b_inv1677 ^ c1677;
  assign and1677 = a1677 & b1677;
  assign or1677  = a1677 | b1677;
  assign c1678 = (a1677 & b1677) | (a1677 & c1677) | (b1677 & c1677);
  wire c_sub1678;
  assign c_sub1678 = (a1677 & b_inv1677) | (a1677 & c1677) | (b_inv1677 & c1677);
  wire s1678, sub1678, and1678, or1678;
  wire b_inv1678;
  assign b_inv1678 = ~b1678;
  assign s1678  = a1678 ^ b1678 ^ c1678;
  assign sub1678 = a1678 ^ b_inv1678 ^ c1678;
  assign and1678 = a1678 & b1678;
  assign or1678  = a1678 | b1678;
  assign c1679 = (a1678 & b1678) | (a1678 & c1678) | (b1678 & c1678);
  wire c_sub1679;
  assign c_sub1679 = (a1678 & b_inv1678) | (a1678 & c1678) | (b_inv1678 & c1678);
  wire s1679, sub1679, and1679, or1679;
  wire b_inv1679;
  assign b_inv1679 = ~b1679;
  assign s1679  = a1679 ^ b1679 ^ c1679;
  assign sub1679 = a1679 ^ b_inv1679 ^ c1679;
  assign and1679 = a1679 & b1679;
  assign or1679  = a1679 | b1679;
  assign c1680 = (a1679 & b1679) | (a1679 & c1679) | (b1679 & c1679);
  wire c_sub1680;
  assign c_sub1680 = (a1679 & b_inv1679) | (a1679 & c1679) | (b_inv1679 & c1679);
  wire s1680, sub1680, and1680, or1680;
  wire b_inv1680;
  assign b_inv1680 = ~b1680;
  assign s1680  = a1680 ^ b1680 ^ c1680;
  assign sub1680 = a1680 ^ b_inv1680 ^ c1680;
  assign and1680 = a1680 & b1680;
  assign or1680  = a1680 | b1680;
  assign c1681 = (a1680 & b1680) | (a1680 & c1680) | (b1680 & c1680);
  wire c_sub1681;
  assign c_sub1681 = (a1680 & b_inv1680) | (a1680 & c1680) | (b_inv1680 & c1680);
  wire s1681, sub1681, and1681, or1681;
  wire b_inv1681;
  assign b_inv1681 = ~b1681;
  assign s1681  = a1681 ^ b1681 ^ c1681;
  assign sub1681 = a1681 ^ b_inv1681 ^ c1681;
  assign and1681 = a1681 & b1681;
  assign or1681  = a1681 | b1681;
  assign c1682 = (a1681 & b1681) | (a1681 & c1681) | (b1681 & c1681);
  wire c_sub1682;
  assign c_sub1682 = (a1681 & b_inv1681) | (a1681 & c1681) | (b_inv1681 & c1681);
  wire s1682, sub1682, and1682, or1682;
  wire b_inv1682;
  assign b_inv1682 = ~b1682;
  assign s1682  = a1682 ^ b1682 ^ c1682;
  assign sub1682 = a1682 ^ b_inv1682 ^ c1682;
  assign and1682 = a1682 & b1682;
  assign or1682  = a1682 | b1682;
  assign c1683 = (a1682 & b1682) | (a1682 & c1682) | (b1682 & c1682);
  wire c_sub1683;
  assign c_sub1683 = (a1682 & b_inv1682) | (a1682 & c1682) | (b_inv1682 & c1682);
  wire s1683, sub1683, and1683, or1683;
  wire b_inv1683;
  assign b_inv1683 = ~b1683;
  assign s1683  = a1683 ^ b1683 ^ c1683;
  assign sub1683 = a1683 ^ b_inv1683 ^ c1683;
  assign and1683 = a1683 & b1683;
  assign or1683  = a1683 | b1683;
  assign c1684 = (a1683 & b1683) | (a1683 & c1683) | (b1683 & c1683);
  wire c_sub1684;
  assign c_sub1684 = (a1683 & b_inv1683) | (a1683 & c1683) | (b_inv1683 & c1683);
  wire s1684, sub1684, and1684, or1684;
  wire b_inv1684;
  assign b_inv1684 = ~b1684;
  assign s1684  = a1684 ^ b1684 ^ c1684;
  assign sub1684 = a1684 ^ b_inv1684 ^ c1684;
  assign and1684 = a1684 & b1684;
  assign or1684  = a1684 | b1684;
  assign c1685 = (a1684 & b1684) | (a1684 & c1684) | (b1684 & c1684);
  wire c_sub1685;
  assign c_sub1685 = (a1684 & b_inv1684) | (a1684 & c1684) | (b_inv1684 & c1684);
  wire s1685, sub1685, and1685, or1685;
  wire b_inv1685;
  assign b_inv1685 = ~b1685;
  assign s1685  = a1685 ^ b1685 ^ c1685;
  assign sub1685 = a1685 ^ b_inv1685 ^ c1685;
  assign and1685 = a1685 & b1685;
  assign or1685  = a1685 | b1685;
  assign c1686 = (a1685 & b1685) | (a1685 & c1685) | (b1685 & c1685);
  wire c_sub1686;
  assign c_sub1686 = (a1685 & b_inv1685) | (a1685 & c1685) | (b_inv1685 & c1685);
  wire s1686, sub1686, and1686, or1686;
  wire b_inv1686;
  assign b_inv1686 = ~b1686;
  assign s1686  = a1686 ^ b1686 ^ c1686;
  assign sub1686 = a1686 ^ b_inv1686 ^ c1686;
  assign and1686 = a1686 & b1686;
  assign or1686  = a1686 | b1686;
  assign c1687 = (a1686 & b1686) | (a1686 & c1686) | (b1686 & c1686);
  wire c_sub1687;
  assign c_sub1687 = (a1686 & b_inv1686) | (a1686 & c1686) | (b_inv1686 & c1686);
  wire s1687, sub1687, and1687, or1687;
  wire b_inv1687;
  assign b_inv1687 = ~b1687;
  assign s1687  = a1687 ^ b1687 ^ c1687;
  assign sub1687 = a1687 ^ b_inv1687 ^ c1687;
  assign and1687 = a1687 & b1687;
  assign or1687  = a1687 | b1687;
  assign c1688 = (a1687 & b1687) | (a1687 & c1687) | (b1687 & c1687);
  wire c_sub1688;
  assign c_sub1688 = (a1687 & b_inv1687) | (a1687 & c1687) | (b_inv1687 & c1687);
  wire s1688, sub1688, and1688, or1688;
  wire b_inv1688;
  assign b_inv1688 = ~b1688;
  assign s1688  = a1688 ^ b1688 ^ c1688;
  assign sub1688 = a1688 ^ b_inv1688 ^ c1688;
  assign and1688 = a1688 & b1688;
  assign or1688  = a1688 | b1688;
  assign c1689 = (a1688 & b1688) | (a1688 & c1688) | (b1688 & c1688);
  wire c_sub1689;
  assign c_sub1689 = (a1688 & b_inv1688) | (a1688 & c1688) | (b_inv1688 & c1688);
  wire s1689, sub1689, and1689, or1689;
  wire b_inv1689;
  assign b_inv1689 = ~b1689;
  assign s1689  = a1689 ^ b1689 ^ c1689;
  assign sub1689 = a1689 ^ b_inv1689 ^ c1689;
  assign and1689 = a1689 & b1689;
  assign or1689  = a1689 | b1689;
  assign c1690 = (a1689 & b1689) | (a1689 & c1689) | (b1689 & c1689);
  wire c_sub1690;
  assign c_sub1690 = (a1689 & b_inv1689) | (a1689 & c1689) | (b_inv1689 & c1689);
  wire s1690, sub1690, and1690, or1690;
  wire b_inv1690;
  assign b_inv1690 = ~b1690;
  assign s1690  = a1690 ^ b1690 ^ c1690;
  assign sub1690 = a1690 ^ b_inv1690 ^ c1690;
  assign and1690 = a1690 & b1690;
  assign or1690  = a1690 | b1690;
  assign c1691 = (a1690 & b1690) | (a1690 & c1690) | (b1690 & c1690);
  wire c_sub1691;
  assign c_sub1691 = (a1690 & b_inv1690) | (a1690 & c1690) | (b_inv1690 & c1690);
  wire s1691, sub1691, and1691, or1691;
  wire b_inv1691;
  assign b_inv1691 = ~b1691;
  assign s1691  = a1691 ^ b1691 ^ c1691;
  assign sub1691 = a1691 ^ b_inv1691 ^ c1691;
  assign and1691 = a1691 & b1691;
  assign or1691  = a1691 | b1691;
  assign c1692 = (a1691 & b1691) | (a1691 & c1691) | (b1691 & c1691);
  wire c_sub1692;
  assign c_sub1692 = (a1691 & b_inv1691) | (a1691 & c1691) | (b_inv1691 & c1691);
  wire s1692, sub1692, and1692, or1692;
  wire b_inv1692;
  assign b_inv1692 = ~b1692;
  assign s1692  = a1692 ^ b1692 ^ c1692;
  assign sub1692 = a1692 ^ b_inv1692 ^ c1692;
  assign and1692 = a1692 & b1692;
  assign or1692  = a1692 | b1692;
  assign c1693 = (a1692 & b1692) | (a1692 & c1692) | (b1692 & c1692);
  wire c_sub1693;
  assign c_sub1693 = (a1692 & b_inv1692) | (a1692 & c1692) | (b_inv1692 & c1692);
  wire s1693, sub1693, and1693, or1693;
  wire b_inv1693;
  assign b_inv1693 = ~b1693;
  assign s1693  = a1693 ^ b1693 ^ c1693;
  assign sub1693 = a1693 ^ b_inv1693 ^ c1693;
  assign and1693 = a1693 & b1693;
  assign or1693  = a1693 | b1693;
  assign c1694 = (a1693 & b1693) | (a1693 & c1693) | (b1693 & c1693);
  wire c_sub1694;
  assign c_sub1694 = (a1693 & b_inv1693) | (a1693 & c1693) | (b_inv1693 & c1693);
  wire s1694, sub1694, and1694, or1694;
  wire b_inv1694;
  assign b_inv1694 = ~b1694;
  assign s1694  = a1694 ^ b1694 ^ c1694;
  assign sub1694 = a1694 ^ b_inv1694 ^ c1694;
  assign and1694 = a1694 & b1694;
  assign or1694  = a1694 | b1694;
  assign c1695 = (a1694 & b1694) | (a1694 & c1694) | (b1694 & c1694);
  wire c_sub1695;
  assign c_sub1695 = (a1694 & b_inv1694) | (a1694 & c1694) | (b_inv1694 & c1694);
  wire s1695, sub1695, and1695, or1695;
  wire b_inv1695;
  assign b_inv1695 = ~b1695;
  assign s1695  = a1695 ^ b1695 ^ c1695;
  assign sub1695 = a1695 ^ b_inv1695 ^ c1695;
  assign and1695 = a1695 & b1695;
  assign or1695  = a1695 | b1695;
  assign c1696 = (a1695 & b1695) | (a1695 & c1695) | (b1695 & c1695);
  wire c_sub1696;
  assign c_sub1696 = (a1695 & b_inv1695) | (a1695 & c1695) | (b_inv1695 & c1695);
  wire s1696, sub1696, and1696, or1696;
  wire b_inv1696;
  assign b_inv1696 = ~b1696;
  assign s1696  = a1696 ^ b1696 ^ c1696;
  assign sub1696 = a1696 ^ b_inv1696 ^ c1696;
  assign and1696 = a1696 & b1696;
  assign or1696  = a1696 | b1696;
  assign c1697 = (a1696 & b1696) | (a1696 & c1696) | (b1696 & c1696);
  wire c_sub1697;
  assign c_sub1697 = (a1696 & b_inv1696) | (a1696 & c1696) | (b_inv1696 & c1696);
  wire s1697, sub1697, and1697, or1697;
  wire b_inv1697;
  assign b_inv1697 = ~b1697;
  assign s1697  = a1697 ^ b1697 ^ c1697;
  assign sub1697 = a1697 ^ b_inv1697 ^ c1697;
  assign and1697 = a1697 & b1697;
  assign or1697  = a1697 | b1697;
  assign c1698 = (a1697 & b1697) | (a1697 & c1697) | (b1697 & c1697);
  wire c_sub1698;
  assign c_sub1698 = (a1697 & b_inv1697) | (a1697 & c1697) | (b_inv1697 & c1697);
  wire s1698, sub1698, and1698, or1698;
  wire b_inv1698;
  assign b_inv1698 = ~b1698;
  assign s1698  = a1698 ^ b1698 ^ c1698;
  assign sub1698 = a1698 ^ b_inv1698 ^ c1698;
  assign and1698 = a1698 & b1698;
  assign or1698  = a1698 | b1698;
  assign c1699 = (a1698 & b1698) | (a1698 & c1698) | (b1698 & c1698);
  wire c_sub1699;
  assign c_sub1699 = (a1698 & b_inv1698) | (a1698 & c1698) | (b_inv1698 & c1698);
  wire s1699, sub1699, and1699, or1699;
  wire b_inv1699;
  assign b_inv1699 = ~b1699;
  assign s1699  = a1699 ^ b1699 ^ c1699;
  assign sub1699 = a1699 ^ b_inv1699 ^ c1699;
  assign and1699 = a1699 & b1699;
  assign or1699  = a1699 | b1699;
  assign c1700 = (a1699 & b1699) | (a1699 & c1699) | (b1699 & c1699);
  wire c_sub1700;
  assign c_sub1700 = (a1699 & b_inv1699) | (a1699 & c1699) | (b_inv1699 & c1699);
  wire s1700, sub1700, and1700, or1700;
  wire b_inv1700;
  assign b_inv1700 = ~b1700;
  assign s1700  = a1700 ^ b1700 ^ c1700;
  assign sub1700 = a1700 ^ b_inv1700 ^ c1700;
  assign and1700 = a1700 & b1700;
  assign or1700  = a1700 | b1700;
  assign c1701 = (a1700 & b1700) | (a1700 & c1700) | (b1700 & c1700);
  wire c_sub1701;
  assign c_sub1701 = (a1700 & b_inv1700) | (a1700 & c1700) | (b_inv1700 & c1700);
  wire s1701, sub1701, and1701, or1701;
  wire b_inv1701;
  assign b_inv1701 = ~b1701;
  assign s1701  = a1701 ^ b1701 ^ c1701;
  assign sub1701 = a1701 ^ b_inv1701 ^ c1701;
  assign and1701 = a1701 & b1701;
  assign or1701  = a1701 | b1701;
  assign c1702 = (a1701 & b1701) | (a1701 & c1701) | (b1701 & c1701);
  wire c_sub1702;
  assign c_sub1702 = (a1701 & b_inv1701) | (a1701 & c1701) | (b_inv1701 & c1701);
  wire s1702, sub1702, and1702, or1702;
  wire b_inv1702;
  assign b_inv1702 = ~b1702;
  assign s1702  = a1702 ^ b1702 ^ c1702;
  assign sub1702 = a1702 ^ b_inv1702 ^ c1702;
  assign and1702 = a1702 & b1702;
  assign or1702  = a1702 | b1702;
  assign c1703 = (a1702 & b1702) | (a1702 & c1702) | (b1702 & c1702);
  wire c_sub1703;
  assign c_sub1703 = (a1702 & b_inv1702) | (a1702 & c1702) | (b_inv1702 & c1702);
  wire s1703, sub1703, and1703, or1703;
  wire b_inv1703;
  assign b_inv1703 = ~b1703;
  assign s1703  = a1703 ^ b1703 ^ c1703;
  assign sub1703 = a1703 ^ b_inv1703 ^ c1703;
  assign and1703 = a1703 & b1703;
  assign or1703  = a1703 | b1703;
  assign c1704 = (a1703 & b1703) | (a1703 & c1703) | (b1703 & c1703);
  wire c_sub1704;
  assign c_sub1704 = (a1703 & b_inv1703) | (a1703 & c1703) | (b_inv1703 & c1703);
  wire s1704, sub1704, and1704, or1704;
  wire b_inv1704;
  assign b_inv1704 = ~b1704;
  assign s1704  = a1704 ^ b1704 ^ c1704;
  assign sub1704 = a1704 ^ b_inv1704 ^ c1704;
  assign and1704 = a1704 & b1704;
  assign or1704  = a1704 | b1704;
  assign c1705 = (a1704 & b1704) | (a1704 & c1704) | (b1704 & c1704);
  wire c_sub1705;
  assign c_sub1705 = (a1704 & b_inv1704) | (a1704 & c1704) | (b_inv1704 & c1704);
  wire s1705, sub1705, and1705, or1705;
  wire b_inv1705;
  assign b_inv1705 = ~b1705;
  assign s1705  = a1705 ^ b1705 ^ c1705;
  assign sub1705 = a1705 ^ b_inv1705 ^ c1705;
  assign and1705 = a1705 & b1705;
  assign or1705  = a1705 | b1705;
  assign c1706 = (a1705 & b1705) | (a1705 & c1705) | (b1705 & c1705);
  wire c_sub1706;
  assign c_sub1706 = (a1705 & b_inv1705) | (a1705 & c1705) | (b_inv1705 & c1705);
  wire s1706, sub1706, and1706, or1706;
  wire b_inv1706;
  assign b_inv1706 = ~b1706;
  assign s1706  = a1706 ^ b1706 ^ c1706;
  assign sub1706 = a1706 ^ b_inv1706 ^ c1706;
  assign and1706 = a1706 & b1706;
  assign or1706  = a1706 | b1706;
  assign c1707 = (a1706 & b1706) | (a1706 & c1706) | (b1706 & c1706);
  wire c_sub1707;
  assign c_sub1707 = (a1706 & b_inv1706) | (a1706 & c1706) | (b_inv1706 & c1706);
  wire s1707, sub1707, and1707, or1707;
  wire b_inv1707;
  assign b_inv1707 = ~b1707;
  assign s1707  = a1707 ^ b1707 ^ c1707;
  assign sub1707 = a1707 ^ b_inv1707 ^ c1707;
  assign and1707 = a1707 & b1707;
  assign or1707  = a1707 | b1707;
  assign c1708 = (a1707 & b1707) | (a1707 & c1707) | (b1707 & c1707);
  wire c_sub1708;
  assign c_sub1708 = (a1707 & b_inv1707) | (a1707 & c1707) | (b_inv1707 & c1707);
  wire s1708, sub1708, and1708, or1708;
  wire b_inv1708;
  assign b_inv1708 = ~b1708;
  assign s1708  = a1708 ^ b1708 ^ c1708;
  assign sub1708 = a1708 ^ b_inv1708 ^ c1708;
  assign and1708 = a1708 & b1708;
  assign or1708  = a1708 | b1708;
  assign c1709 = (a1708 & b1708) | (a1708 & c1708) | (b1708 & c1708);
  wire c_sub1709;
  assign c_sub1709 = (a1708 & b_inv1708) | (a1708 & c1708) | (b_inv1708 & c1708);
  wire s1709, sub1709, and1709, or1709;
  wire b_inv1709;
  assign b_inv1709 = ~b1709;
  assign s1709  = a1709 ^ b1709 ^ c1709;
  assign sub1709 = a1709 ^ b_inv1709 ^ c1709;
  assign and1709 = a1709 & b1709;
  assign or1709  = a1709 | b1709;
  assign c1710 = (a1709 & b1709) | (a1709 & c1709) | (b1709 & c1709);
  wire c_sub1710;
  assign c_sub1710 = (a1709 & b_inv1709) | (a1709 & c1709) | (b_inv1709 & c1709);
  wire s1710, sub1710, and1710, or1710;
  wire b_inv1710;
  assign b_inv1710 = ~b1710;
  assign s1710  = a1710 ^ b1710 ^ c1710;
  assign sub1710 = a1710 ^ b_inv1710 ^ c1710;
  assign and1710 = a1710 & b1710;
  assign or1710  = a1710 | b1710;
  assign c1711 = (a1710 & b1710) | (a1710 & c1710) | (b1710 & c1710);
  wire c_sub1711;
  assign c_sub1711 = (a1710 & b_inv1710) | (a1710 & c1710) | (b_inv1710 & c1710);
  wire s1711, sub1711, and1711, or1711;
  wire b_inv1711;
  assign b_inv1711 = ~b1711;
  assign s1711  = a1711 ^ b1711 ^ c1711;
  assign sub1711 = a1711 ^ b_inv1711 ^ c1711;
  assign and1711 = a1711 & b1711;
  assign or1711  = a1711 | b1711;
  assign c1712 = (a1711 & b1711) | (a1711 & c1711) | (b1711 & c1711);
  wire c_sub1712;
  assign c_sub1712 = (a1711 & b_inv1711) | (a1711 & c1711) | (b_inv1711 & c1711);
  wire s1712, sub1712, and1712, or1712;
  wire b_inv1712;
  assign b_inv1712 = ~b1712;
  assign s1712  = a1712 ^ b1712 ^ c1712;
  assign sub1712 = a1712 ^ b_inv1712 ^ c1712;
  assign and1712 = a1712 & b1712;
  assign or1712  = a1712 | b1712;
  assign c1713 = (a1712 & b1712) | (a1712 & c1712) | (b1712 & c1712);
  wire c_sub1713;
  assign c_sub1713 = (a1712 & b_inv1712) | (a1712 & c1712) | (b_inv1712 & c1712);
  wire s1713, sub1713, and1713, or1713;
  wire b_inv1713;
  assign b_inv1713 = ~b1713;
  assign s1713  = a1713 ^ b1713 ^ c1713;
  assign sub1713 = a1713 ^ b_inv1713 ^ c1713;
  assign and1713 = a1713 & b1713;
  assign or1713  = a1713 | b1713;
  assign c1714 = (a1713 & b1713) | (a1713 & c1713) | (b1713 & c1713);
  wire c_sub1714;
  assign c_sub1714 = (a1713 & b_inv1713) | (a1713 & c1713) | (b_inv1713 & c1713);
  wire s1714, sub1714, and1714, or1714;
  wire b_inv1714;
  assign b_inv1714 = ~b1714;
  assign s1714  = a1714 ^ b1714 ^ c1714;
  assign sub1714 = a1714 ^ b_inv1714 ^ c1714;
  assign and1714 = a1714 & b1714;
  assign or1714  = a1714 | b1714;
  assign c1715 = (a1714 & b1714) | (a1714 & c1714) | (b1714 & c1714);
  wire c_sub1715;
  assign c_sub1715 = (a1714 & b_inv1714) | (a1714 & c1714) | (b_inv1714 & c1714);
  wire s1715, sub1715, and1715, or1715;
  wire b_inv1715;
  assign b_inv1715 = ~b1715;
  assign s1715  = a1715 ^ b1715 ^ c1715;
  assign sub1715 = a1715 ^ b_inv1715 ^ c1715;
  assign and1715 = a1715 & b1715;
  assign or1715  = a1715 | b1715;
  assign c1716 = (a1715 & b1715) | (a1715 & c1715) | (b1715 & c1715);
  wire c_sub1716;
  assign c_sub1716 = (a1715 & b_inv1715) | (a1715 & c1715) | (b_inv1715 & c1715);
  wire s1716, sub1716, and1716, or1716;
  wire b_inv1716;
  assign b_inv1716 = ~b1716;
  assign s1716  = a1716 ^ b1716 ^ c1716;
  assign sub1716 = a1716 ^ b_inv1716 ^ c1716;
  assign and1716 = a1716 & b1716;
  assign or1716  = a1716 | b1716;
  assign c1717 = (a1716 & b1716) | (a1716 & c1716) | (b1716 & c1716);
  wire c_sub1717;
  assign c_sub1717 = (a1716 & b_inv1716) | (a1716 & c1716) | (b_inv1716 & c1716);
  wire s1717, sub1717, and1717, or1717;
  wire b_inv1717;
  assign b_inv1717 = ~b1717;
  assign s1717  = a1717 ^ b1717 ^ c1717;
  assign sub1717 = a1717 ^ b_inv1717 ^ c1717;
  assign and1717 = a1717 & b1717;
  assign or1717  = a1717 | b1717;
  assign c1718 = (a1717 & b1717) | (a1717 & c1717) | (b1717 & c1717);
  wire c_sub1718;
  assign c_sub1718 = (a1717 & b_inv1717) | (a1717 & c1717) | (b_inv1717 & c1717);
  wire s1718, sub1718, and1718, or1718;
  wire b_inv1718;
  assign b_inv1718 = ~b1718;
  assign s1718  = a1718 ^ b1718 ^ c1718;
  assign sub1718 = a1718 ^ b_inv1718 ^ c1718;
  assign and1718 = a1718 & b1718;
  assign or1718  = a1718 | b1718;
  assign c1719 = (a1718 & b1718) | (a1718 & c1718) | (b1718 & c1718);
  wire c_sub1719;
  assign c_sub1719 = (a1718 & b_inv1718) | (a1718 & c1718) | (b_inv1718 & c1718);
  wire s1719, sub1719, and1719, or1719;
  wire b_inv1719;
  assign b_inv1719 = ~b1719;
  assign s1719  = a1719 ^ b1719 ^ c1719;
  assign sub1719 = a1719 ^ b_inv1719 ^ c1719;
  assign and1719 = a1719 & b1719;
  assign or1719  = a1719 | b1719;
  assign c1720 = (a1719 & b1719) | (a1719 & c1719) | (b1719 & c1719);
  wire c_sub1720;
  assign c_sub1720 = (a1719 & b_inv1719) | (a1719 & c1719) | (b_inv1719 & c1719);
  wire s1720, sub1720, and1720, or1720;
  wire b_inv1720;
  assign b_inv1720 = ~b1720;
  assign s1720  = a1720 ^ b1720 ^ c1720;
  assign sub1720 = a1720 ^ b_inv1720 ^ c1720;
  assign and1720 = a1720 & b1720;
  assign or1720  = a1720 | b1720;
  assign c1721 = (a1720 & b1720) | (a1720 & c1720) | (b1720 & c1720);
  wire c_sub1721;
  assign c_sub1721 = (a1720 & b_inv1720) | (a1720 & c1720) | (b_inv1720 & c1720);
  wire s1721, sub1721, and1721, or1721;
  wire b_inv1721;
  assign b_inv1721 = ~b1721;
  assign s1721  = a1721 ^ b1721 ^ c1721;
  assign sub1721 = a1721 ^ b_inv1721 ^ c1721;
  assign and1721 = a1721 & b1721;
  assign or1721  = a1721 | b1721;
  assign c1722 = (a1721 & b1721) | (a1721 & c1721) | (b1721 & c1721);
  wire c_sub1722;
  assign c_sub1722 = (a1721 & b_inv1721) | (a1721 & c1721) | (b_inv1721 & c1721);
  wire s1722, sub1722, and1722, or1722;
  wire b_inv1722;
  assign b_inv1722 = ~b1722;
  assign s1722  = a1722 ^ b1722 ^ c1722;
  assign sub1722 = a1722 ^ b_inv1722 ^ c1722;
  assign and1722 = a1722 & b1722;
  assign or1722  = a1722 | b1722;
  assign c1723 = (a1722 & b1722) | (a1722 & c1722) | (b1722 & c1722);
  wire c_sub1723;
  assign c_sub1723 = (a1722 & b_inv1722) | (a1722 & c1722) | (b_inv1722 & c1722);
  wire s1723, sub1723, and1723, or1723;
  wire b_inv1723;
  assign b_inv1723 = ~b1723;
  assign s1723  = a1723 ^ b1723 ^ c1723;
  assign sub1723 = a1723 ^ b_inv1723 ^ c1723;
  assign and1723 = a1723 & b1723;
  assign or1723  = a1723 | b1723;
  assign c1724 = (a1723 & b1723) | (a1723 & c1723) | (b1723 & c1723);
  wire c_sub1724;
  assign c_sub1724 = (a1723 & b_inv1723) | (a1723 & c1723) | (b_inv1723 & c1723);
  wire s1724, sub1724, and1724, or1724;
  wire b_inv1724;
  assign b_inv1724 = ~b1724;
  assign s1724  = a1724 ^ b1724 ^ c1724;
  assign sub1724 = a1724 ^ b_inv1724 ^ c1724;
  assign and1724 = a1724 & b1724;
  assign or1724  = a1724 | b1724;
  assign c1725 = (a1724 & b1724) | (a1724 & c1724) | (b1724 & c1724);
  wire c_sub1725;
  assign c_sub1725 = (a1724 & b_inv1724) | (a1724 & c1724) | (b_inv1724 & c1724);
  wire s1725, sub1725, and1725, or1725;
  wire b_inv1725;
  assign b_inv1725 = ~b1725;
  assign s1725  = a1725 ^ b1725 ^ c1725;
  assign sub1725 = a1725 ^ b_inv1725 ^ c1725;
  assign and1725 = a1725 & b1725;
  assign or1725  = a1725 | b1725;
  assign c1726 = (a1725 & b1725) | (a1725 & c1725) | (b1725 & c1725);
  wire c_sub1726;
  assign c_sub1726 = (a1725 & b_inv1725) | (a1725 & c1725) | (b_inv1725 & c1725);
  wire s1726, sub1726, and1726, or1726;
  wire b_inv1726;
  assign b_inv1726 = ~b1726;
  assign s1726  = a1726 ^ b1726 ^ c1726;
  assign sub1726 = a1726 ^ b_inv1726 ^ c1726;
  assign and1726 = a1726 & b1726;
  assign or1726  = a1726 | b1726;
  assign c1727 = (a1726 & b1726) | (a1726 & c1726) | (b1726 & c1726);
  wire c_sub1727;
  assign c_sub1727 = (a1726 & b_inv1726) | (a1726 & c1726) | (b_inv1726 & c1726);
  wire s1727, sub1727, and1727, or1727;
  wire b_inv1727;
  assign b_inv1727 = ~b1727;
  assign s1727  = a1727 ^ b1727 ^ c1727;
  assign sub1727 = a1727 ^ b_inv1727 ^ c1727;
  assign and1727 = a1727 & b1727;
  assign or1727  = a1727 | b1727;
  assign c1728 = (a1727 & b1727) | (a1727 & c1727) | (b1727 & c1727);
  wire c_sub1728;
  assign c_sub1728 = (a1727 & b_inv1727) | (a1727 & c1727) | (b_inv1727 & c1727);
  wire s1728, sub1728, and1728, or1728;
  wire b_inv1728;
  assign b_inv1728 = ~b1728;
  assign s1728  = a1728 ^ b1728 ^ c1728;
  assign sub1728 = a1728 ^ b_inv1728 ^ c1728;
  assign and1728 = a1728 & b1728;
  assign or1728  = a1728 | b1728;
  assign c1729 = (a1728 & b1728) | (a1728 & c1728) | (b1728 & c1728);
  wire c_sub1729;
  assign c_sub1729 = (a1728 & b_inv1728) | (a1728 & c1728) | (b_inv1728 & c1728);
  wire s1729, sub1729, and1729, or1729;
  wire b_inv1729;
  assign b_inv1729 = ~b1729;
  assign s1729  = a1729 ^ b1729 ^ c1729;
  assign sub1729 = a1729 ^ b_inv1729 ^ c1729;
  assign and1729 = a1729 & b1729;
  assign or1729  = a1729 | b1729;
  assign c1730 = (a1729 & b1729) | (a1729 & c1729) | (b1729 & c1729);
  wire c_sub1730;
  assign c_sub1730 = (a1729 & b_inv1729) | (a1729 & c1729) | (b_inv1729 & c1729);
  wire s1730, sub1730, and1730, or1730;
  wire b_inv1730;
  assign b_inv1730 = ~b1730;
  assign s1730  = a1730 ^ b1730 ^ c1730;
  assign sub1730 = a1730 ^ b_inv1730 ^ c1730;
  assign and1730 = a1730 & b1730;
  assign or1730  = a1730 | b1730;
  assign c1731 = (a1730 & b1730) | (a1730 & c1730) | (b1730 & c1730);
  wire c_sub1731;
  assign c_sub1731 = (a1730 & b_inv1730) | (a1730 & c1730) | (b_inv1730 & c1730);
  wire s1731, sub1731, and1731, or1731;
  wire b_inv1731;
  assign b_inv1731 = ~b1731;
  assign s1731  = a1731 ^ b1731 ^ c1731;
  assign sub1731 = a1731 ^ b_inv1731 ^ c1731;
  assign and1731 = a1731 & b1731;
  assign or1731  = a1731 | b1731;
  assign c1732 = (a1731 & b1731) | (a1731 & c1731) | (b1731 & c1731);
  wire c_sub1732;
  assign c_sub1732 = (a1731 & b_inv1731) | (a1731 & c1731) | (b_inv1731 & c1731);
  wire s1732, sub1732, and1732, or1732;
  wire b_inv1732;
  assign b_inv1732 = ~b1732;
  assign s1732  = a1732 ^ b1732 ^ c1732;
  assign sub1732 = a1732 ^ b_inv1732 ^ c1732;
  assign and1732 = a1732 & b1732;
  assign or1732  = a1732 | b1732;
  assign c1733 = (a1732 & b1732) | (a1732 & c1732) | (b1732 & c1732);
  wire c_sub1733;
  assign c_sub1733 = (a1732 & b_inv1732) | (a1732 & c1732) | (b_inv1732 & c1732);
  wire s1733, sub1733, and1733, or1733;
  wire b_inv1733;
  assign b_inv1733 = ~b1733;
  assign s1733  = a1733 ^ b1733 ^ c1733;
  assign sub1733 = a1733 ^ b_inv1733 ^ c1733;
  assign and1733 = a1733 & b1733;
  assign or1733  = a1733 | b1733;
  assign c1734 = (a1733 & b1733) | (a1733 & c1733) | (b1733 & c1733);
  wire c_sub1734;
  assign c_sub1734 = (a1733 & b_inv1733) | (a1733 & c1733) | (b_inv1733 & c1733);
  wire s1734, sub1734, and1734, or1734;
  wire b_inv1734;
  assign b_inv1734 = ~b1734;
  assign s1734  = a1734 ^ b1734 ^ c1734;
  assign sub1734 = a1734 ^ b_inv1734 ^ c1734;
  assign and1734 = a1734 & b1734;
  assign or1734  = a1734 | b1734;
  assign c1735 = (a1734 & b1734) | (a1734 & c1734) | (b1734 & c1734);
  wire c_sub1735;
  assign c_sub1735 = (a1734 & b_inv1734) | (a1734 & c1734) | (b_inv1734 & c1734);
  wire s1735, sub1735, and1735, or1735;
  wire b_inv1735;
  assign b_inv1735 = ~b1735;
  assign s1735  = a1735 ^ b1735 ^ c1735;
  assign sub1735 = a1735 ^ b_inv1735 ^ c1735;
  assign and1735 = a1735 & b1735;
  assign or1735  = a1735 | b1735;
  assign c1736 = (a1735 & b1735) | (a1735 & c1735) | (b1735 & c1735);
  wire c_sub1736;
  assign c_sub1736 = (a1735 & b_inv1735) | (a1735 & c1735) | (b_inv1735 & c1735);
  wire s1736, sub1736, and1736, or1736;
  wire b_inv1736;
  assign b_inv1736 = ~b1736;
  assign s1736  = a1736 ^ b1736 ^ c1736;
  assign sub1736 = a1736 ^ b_inv1736 ^ c1736;
  assign and1736 = a1736 & b1736;
  assign or1736  = a1736 | b1736;
  assign c1737 = (a1736 & b1736) | (a1736 & c1736) | (b1736 & c1736);
  wire c_sub1737;
  assign c_sub1737 = (a1736 & b_inv1736) | (a1736 & c1736) | (b_inv1736 & c1736);
  wire s1737, sub1737, and1737, or1737;
  wire b_inv1737;
  assign b_inv1737 = ~b1737;
  assign s1737  = a1737 ^ b1737 ^ c1737;
  assign sub1737 = a1737 ^ b_inv1737 ^ c1737;
  assign and1737 = a1737 & b1737;
  assign or1737  = a1737 | b1737;
  assign c1738 = (a1737 & b1737) | (a1737 & c1737) | (b1737 & c1737);
  wire c_sub1738;
  assign c_sub1738 = (a1737 & b_inv1737) | (a1737 & c1737) | (b_inv1737 & c1737);
  wire s1738, sub1738, and1738, or1738;
  wire b_inv1738;
  assign b_inv1738 = ~b1738;
  assign s1738  = a1738 ^ b1738 ^ c1738;
  assign sub1738 = a1738 ^ b_inv1738 ^ c1738;
  assign and1738 = a1738 & b1738;
  assign or1738  = a1738 | b1738;
  assign c1739 = (a1738 & b1738) | (a1738 & c1738) | (b1738 & c1738);
  wire c_sub1739;
  assign c_sub1739 = (a1738 & b_inv1738) | (a1738 & c1738) | (b_inv1738 & c1738);
  wire s1739, sub1739, and1739, or1739;
  wire b_inv1739;
  assign b_inv1739 = ~b1739;
  assign s1739  = a1739 ^ b1739 ^ c1739;
  assign sub1739 = a1739 ^ b_inv1739 ^ c1739;
  assign and1739 = a1739 & b1739;
  assign or1739  = a1739 | b1739;
  assign c1740 = (a1739 & b1739) | (a1739 & c1739) | (b1739 & c1739);
  wire c_sub1740;
  assign c_sub1740 = (a1739 & b_inv1739) | (a1739 & c1739) | (b_inv1739 & c1739);
  wire s1740, sub1740, and1740, or1740;
  wire b_inv1740;
  assign b_inv1740 = ~b1740;
  assign s1740  = a1740 ^ b1740 ^ c1740;
  assign sub1740 = a1740 ^ b_inv1740 ^ c1740;
  assign and1740 = a1740 & b1740;
  assign or1740  = a1740 | b1740;
  assign c1741 = (a1740 & b1740) | (a1740 & c1740) | (b1740 & c1740);
  wire c_sub1741;
  assign c_sub1741 = (a1740 & b_inv1740) | (a1740 & c1740) | (b_inv1740 & c1740);
  wire s1741, sub1741, and1741, or1741;
  wire b_inv1741;
  assign b_inv1741 = ~b1741;
  assign s1741  = a1741 ^ b1741 ^ c1741;
  assign sub1741 = a1741 ^ b_inv1741 ^ c1741;
  assign and1741 = a1741 & b1741;
  assign or1741  = a1741 | b1741;
  assign c1742 = (a1741 & b1741) | (a1741 & c1741) | (b1741 & c1741);
  wire c_sub1742;
  assign c_sub1742 = (a1741 & b_inv1741) | (a1741 & c1741) | (b_inv1741 & c1741);
  wire s1742, sub1742, and1742, or1742;
  wire b_inv1742;
  assign b_inv1742 = ~b1742;
  assign s1742  = a1742 ^ b1742 ^ c1742;
  assign sub1742 = a1742 ^ b_inv1742 ^ c1742;
  assign and1742 = a1742 & b1742;
  assign or1742  = a1742 | b1742;
  assign c1743 = (a1742 & b1742) | (a1742 & c1742) | (b1742 & c1742);
  wire c_sub1743;
  assign c_sub1743 = (a1742 & b_inv1742) | (a1742 & c1742) | (b_inv1742 & c1742);
  wire s1743, sub1743, and1743, or1743;
  wire b_inv1743;
  assign b_inv1743 = ~b1743;
  assign s1743  = a1743 ^ b1743 ^ c1743;
  assign sub1743 = a1743 ^ b_inv1743 ^ c1743;
  assign and1743 = a1743 & b1743;
  assign or1743  = a1743 | b1743;
  assign c1744 = (a1743 & b1743) | (a1743 & c1743) | (b1743 & c1743);
  wire c_sub1744;
  assign c_sub1744 = (a1743 & b_inv1743) | (a1743 & c1743) | (b_inv1743 & c1743);
  wire s1744, sub1744, and1744, or1744;
  wire b_inv1744;
  assign b_inv1744 = ~b1744;
  assign s1744  = a1744 ^ b1744 ^ c1744;
  assign sub1744 = a1744 ^ b_inv1744 ^ c1744;
  assign and1744 = a1744 & b1744;
  assign or1744  = a1744 | b1744;
  assign c1745 = (a1744 & b1744) | (a1744 & c1744) | (b1744 & c1744);
  wire c_sub1745;
  assign c_sub1745 = (a1744 & b_inv1744) | (a1744 & c1744) | (b_inv1744 & c1744);
  wire s1745, sub1745, and1745, or1745;
  wire b_inv1745;
  assign b_inv1745 = ~b1745;
  assign s1745  = a1745 ^ b1745 ^ c1745;
  assign sub1745 = a1745 ^ b_inv1745 ^ c1745;
  assign and1745 = a1745 & b1745;
  assign or1745  = a1745 | b1745;
  assign c1746 = (a1745 & b1745) | (a1745 & c1745) | (b1745 & c1745);
  wire c_sub1746;
  assign c_sub1746 = (a1745 & b_inv1745) | (a1745 & c1745) | (b_inv1745 & c1745);
  wire s1746, sub1746, and1746, or1746;
  wire b_inv1746;
  assign b_inv1746 = ~b1746;
  assign s1746  = a1746 ^ b1746 ^ c1746;
  assign sub1746 = a1746 ^ b_inv1746 ^ c1746;
  assign and1746 = a1746 & b1746;
  assign or1746  = a1746 | b1746;
  assign c1747 = (a1746 & b1746) | (a1746 & c1746) | (b1746 & c1746);
  wire c_sub1747;
  assign c_sub1747 = (a1746 & b_inv1746) | (a1746 & c1746) | (b_inv1746 & c1746);
  wire s1747, sub1747, and1747, or1747;
  wire b_inv1747;
  assign b_inv1747 = ~b1747;
  assign s1747  = a1747 ^ b1747 ^ c1747;
  assign sub1747 = a1747 ^ b_inv1747 ^ c1747;
  assign and1747 = a1747 & b1747;
  assign or1747  = a1747 | b1747;
  assign c1748 = (a1747 & b1747) | (a1747 & c1747) | (b1747 & c1747);
  wire c_sub1748;
  assign c_sub1748 = (a1747 & b_inv1747) | (a1747 & c1747) | (b_inv1747 & c1747);
  wire s1748, sub1748, and1748, or1748;
  wire b_inv1748;
  assign b_inv1748 = ~b1748;
  assign s1748  = a1748 ^ b1748 ^ c1748;
  assign sub1748 = a1748 ^ b_inv1748 ^ c1748;
  assign and1748 = a1748 & b1748;
  assign or1748  = a1748 | b1748;
  assign c1749 = (a1748 & b1748) | (a1748 & c1748) | (b1748 & c1748);
  wire c_sub1749;
  assign c_sub1749 = (a1748 & b_inv1748) | (a1748 & c1748) | (b_inv1748 & c1748);
  wire s1749, sub1749, and1749, or1749;
  wire b_inv1749;
  assign b_inv1749 = ~b1749;
  assign s1749  = a1749 ^ b1749 ^ c1749;
  assign sub1749 = a1749 ^ b_inv1749 ^ c1749;
  assign and1749 = a1749 & b1749;
  assign or1749  = a1749 | b1749;
  assign c1750 = (a1749 & b1749) | (a1749 & c1749) | (b1749 & c1749);
  wire c_sub1750;
  assign c_sub1750 = (a1749 & b_inv1749) | (a1749 & c1749) | (b_inv1749 & c1749);
  wire s1750, sub1750, and1750, or1750;
  wire b_inv1750;
  assign b_inv1750 = ~b1750;
  assign s1750  = a1750 ^ b1750 ^ c1750;
  assign sub1750 = a1750 ^ b_inv1750 ^ c1750;
  assign and1750 = a1750 & b1750;
  assign or1750  = a1750 | b1750;
  assign c1751 = (a1750 & b1750) | (a1750 & c1750) | (b1750 & c1750);
  wire c_sub1751;
  assign c_sub1751 = (a1750 & b_inv1750) | (a1750 & c1750) | (b_inv1750 & c1750);
  wire s1751, sub1751, and1751, or1751;
  wire b_inv1751;
  assign b_inv1751 = ~b1751;
  assign s1751  = a1751 ^ b1751 ^ c1751;
  assign sub1751 = a1751 ^ b_inv1751 ^ c1751;
  assign and1751 = a1751 & b1751;
  assign or1751  = a1751 | b1751;
  assign c1752 = (a1751 & b1751) | (a1751 & c1751) | (b1751 & c1751);
  wire c_sub1752;
  assign c_sub1752 = (a1751 & b_inv1751) | (a1751 & c1751) | (b_inv1751 & c1751);
  wire s1752, sub1752, and1752, or1752;
  wire b_inv1752;
  assign b_inv1752 = ~b1752;
  assign s1752  = a1752 ^ b1752 ^ c1752;
  assign sub1752 = a1752 ^ b_inv1752 ^ c1752;
  assign and1752 = a1752 & b1752;
  assign or1752  = a1752 | b1752;
  assign c1753 = (a1752 & b1752) | (a1752 & c1752) | (b1752 & c1752);
  wire c_sub1753;
  assign c_sub1753 = (a1752 & b_inv1752) | (a1752 & c1752) | (b_inv1752 & c1752);
  wire s1753, sub1753, and1753, or1753;
  wire b_inv1753;
  assign b_inv1753 = ~b1753;
  assign s1753  = a1753 ^ b1753 ^ c1753;
  assign sub1753 = a1753 ^ b_inv1753 ^ c1753;
  assign and1753 = a1753 & b1753;
  assign or1753  = a1753 | b1753;
  assign c1754 = (a1753 & b1753) | (a1753 & c1753) | (b1753 & c1753);
  wire c_sub1754;
  assign c_sub1754 = (a1753 & b_inv1753) | (a1753 & c1753) | (b_inv1753 & c1753);
  wire s1754, sub1754, and1754, or1754;
  wire b_inv1754;
  assign b_inv1754 = ~b1754;
  assign s1754  = a1754 ^ b1754 ^ c1754;
  assign sub1754 = a1754 ^ b_inv1754 ^ c1754;
  assign and1754 = a1754 & b1754;
  assign or1754  = a1754 | b1754;
  assign c1755 = (a1754 & b1754) | (a1754 & c1754) | (b1754 & c1754);
  wire c_sub1755;
  assign c_sub1755 = (a1754 & b_inv1754) | (a1754 & c1754) | (b_inv1754 & c1754);
  wire s1755, sub1755, and1755, or1755;
  wire b_inv1755;
  assign b_inv1755 = ~b1755;
  assign s1755  = a1755 ^ b1755 ^ c1755;
  assign sub1755 = a1755 ^ b_inv1755 ^ c1755;
  assign and1755 = a1755 & b1755;
  assign or1755  = a1755 | b1755;
  assign c1756 = (a1755 & b1755) | (a1755 & c1755) | (b1755 & c1755);
  wire c_sub1756;
  assign c_sub1756 = (a1755 & b_inv1755) | (a1755 & c1755) | (b_inv1755 & c1755);
  wire s1756, sub1756, and1756, or1756;
  wire b_inv1756;
  assign b_inv1756 = ~b1756;
  assign s1756  = a1756 ^ b1756 ^ c1756;
  assign sub1756 = a1756 ^ b_inv1756 ^ c1756;
  assign and1756 = a1756 & b1756;
  assign or1756  = a1756 | b1756;
  assign c1757 = (a1756 & b1756) | (a1756 & c1756) | (b1756 & c1756);
  wire c_sub1757;
  assign c_sub1757 = (a1756 & b_inv1756) | (a1756 & c1756) | (b_inv1756 & c1756);
  wire s1757, sub1757, and1757, or1757;
  wire b_inv1757;
  assign b_inv1757 = ~b1757;
  assign s1757  = a1757 ^ b1757 ^ c1757;
  assign sub1757 = a1757 ^ b_inv1757 ^ c1757;
  assign and1757 = a1757 & b1757;
  assign or1757  = a1757 | b1757;
  assign c1758 = (a1757 & b1757) | (a1757 & c1757) | (b1757 & c1757);
  wire c_sub1758;
  assign c_sub1758 = (a1757 & b_inv1757) | (a1757 & c1757) | (b_inv1757 & c1757);
  wire s1758, sub1758, and1758, or1758;
  wire b_inv1758;
  assign b_inv1758 = ~b1758;
  assign s1758  = a1758 ^ b1758 ^ c1758;
  assign sub1758 = a1758 ^ b_inv1758 ^ c1758;
  assign and1758 = a1758 & b1758;
  assign or1758  = a1758 | b1758;
  assign c1759 = (a1758 & b1758) | (a1758 & c1758) | (b1758 & c1758);
  wire c_sub1759;
  assign c_sub1759 = (a1758 & b_inv1758) | (a1758 & c1758) | (b_inv1758 & c1758);
  wire s1759, sub1759, and1759, or1759;
  wire b_inv1759;
  assign b_inv1759 = ~b1759;
  assign s1759  = a1759 ^ b1759 ^ c1759;
  assign sub1759 = a1759 ^ b_inv1759 ^ c1759;
  assign and1759 = a1759 & b1759;
  assign or1759  = a1759 | b1759;
  assign c1760 = (a1759 & b1759) | (a1759 & c1759) | (b1759 & c1759);
  wire c_sub1760;
  assign c_sub1760 = (a1759 & b_inv1759) | (a1759 & c1759) | (b_inv1759 & c1759);
  wire s1760, sub1760, and1760, or1760;
  wire b_inv1760;
  assign b_inv1760 = ~b1760;
  assign s1760  = a1760 ^ b1760 ^ c1760;
  assign sub1760 = a1760 ^ b_inv1760 ^ c1760;
  assign and1760 = a1760 & b1760;
  assign or1760  = a1760 | b1760;
  assign c1761 = (a1760 & b1760) | (a1760 & c1760) | (b1760 & c1760);
  wire c_sub1761;
  assign c_sub1761 = (a1760 & b_inv1760) | (a1760 & c1760) | (b_inv1760 & c1760);
  wire s1761, sub1761, and1761, or1761;
  wire b_inv1761;
  assign b_inv1761 = ~b1761;
  assign s1761  = a1761 ^ b1761 ^ c1761;
  assign sub1761 = a1761 ^ b_inv1761 ^ c1761;
  assign and1761 = a1761 & b1761;
  assign or1761  = a1761 | b1761;
  assign c1762 = (a1761 & b1761) | (a1761 & c1761) | (b1761 & c1761);
  wire c_sub1762;
  assign c_sub1762 = (a1761 & b_inv1761) | (a1761 & c1761) | (b_inv1761 & c1761);
  wire s1762, sub1762, and1762, or1762;
  wire b_inv1762;
  assign b_inv1762 = ~b1762;
  assign s1762  = a1762 ^ b1762 ^ c1762;
  assign sub1762 = a1762 ^ b_inv1762 ^ c1762;
  assign and1762 = a1762 & b1762;
  assign or1762  = a1762 | b1762;
  assign c1763 = (a1762 & b1762) | (a1762 & c1762) | (b1762 & c1762);
  wire c_sub1763;
  assign c_sub1763 = (a1762 & b_inv1762) | (a1762 & c1762) | (b_inv1762 & c1762);
  wire s1763, sub1763, and1763, or1763;
  wire b_inv1763;
  assign b_inv1763 = ~b1763;
  assign s1763  = a1763 ^ b1763 ^ c1763;
  assign sub1763 = a1763 ^ b_inv1763 ^ c1763;
  assign and1763 = a1763 & b1763;
  assign or1763  = a1763 | b1763;
  assign c1764 = (a1763 & b1763) | (a1763 & c1763) | (b1763 & c1763);
  wire c_sub1764;
  assign c_sub1764 = (a1763 & b_inv1763) | (a1763 & c1763) | (b_inv1763 & c1763);
  wire s1764, sub1764, and1764, or1764;
  wire b_inv1764;
  assign b_inv1764 = ~b1764;
  assign s1764  = a1764 ^ b1764 ^ c1764;
  assign sub1764 = a1764 ^ b_inv1764 ^ c1764;
  assign and1764 = a1764 & b1764;
  assign or1764  = a1764 | b1764;
  assign c1765 = (a1764 & b1764) | (a1764 & c1764) | (b1764 & c1764);
  wire c_sub1765;
  assign c_sub1765 = (a1764 & b_inv1764) | (a1764 & c1764) | (b_inv1764 & c1764);
  wire s1765, sub1765, and1765, or1765;
  wire b_inv1765;
  assign b_inv1765 = ~b1765;
  assign s1765  = a1765 ^ b1765 ^ c1765;
  assign sub1765 = a1765 ^ b_inv1765 ^ c1765;
  assign and1765 = a1765 & b1765;
  assign or1765  = a1765 | b1765;
  assign c1766 = (a1765 & b1765) | (a1765 & c1765) | (b1765 & c1765);
  wire c_sub1766;
  assign c_sub1766 = (a1765 & b_inv1765) | (a1765 & c1765) | (b_inv1765 & c1765);
  wire s1766, sub1766, and1766, or1766;
  wire b_inv1766;
  assign b_inv1766 = ~b1766;
  assign s1766  = a1766 ^ b1766 ^ c1766;
  assign sub1766 = a1766 ^ b_inv1766 ^ c1766;
  assign and1766 = a1766 & b1766;
  assign or1766  = a1766 | b1766;
  assign c1767 = (a1766 & b1766) | (a1766 & c1766) | (b1766 & c1766);
  wire c_sub1767;
  assign c_sub1767 = (a1766 & b_inv1766) | (a1766 & c1766) | (b_inv1766 & c1766);
  wire s1767, sub1767, and1767, or1767;
  wire b_inv1767;
  assign b_inv1767 = ~b1767;
  assign s1767  = a1767 ^ b1767 ^ c1767;
  assign sub1767 = a1767 ^ b_inv1767 ^ c1767;
  assign and1767 = a1767 & b1767;
  assign or1767  = a1767 | b1767;
  assign c1768 = (a1767 & b1767) | (a1767 & c1767) | (b1767 & c1767);
  wire c_sub1768;
  assign c_sub1768 = (a1767 & b_inv1767) | (a1767 & c1767) | (b_inv1767 & c1767);
  wire s1768, sub1768, and1768, or1768;
  wire b_inv1768;
  assign b_inv1768 = ~b1768;
  assign s1768  = a1768 ^ b1768 ^ c1768;
  assign sub1768 = a1768 ^ b_inv1768 ^ c1768;
  assign and1768 = a1768 & b1768;
  assign or1768  = a1768 | b1768;
  assign c1769 = (a1768 & b1768) | (a1768 & c1768) | (b1768 & c1768);
  wire c_sub1769;
  assign c_sub1769 = (a1768 & b_inv1768) | (a1768 & c1768) | (b_inv1768 & c1768);
  wire s1769, sub1769, and1769, or1769;
  wire b_inv1769;
  assign b_inv1769 = ~b1769;
  assign s1769  = a1769 ^ b1769 ^ c1769;
  assign sub1769 = a1769 ^ b_inv1769 ^ c1769;
  assign and1769 = a1769 & b1769;
  assign or1769  = a1769 | b1769;
  assign c1770 = (a1769 & b1769) | (a1769 & c1769) | (b1769 & c1769);
  wire c_sub1770;
  assign c_sub1770 = (a1769 & b_inv1769) | (a1769 & c1769) | (b_inv1769 & c1769);
  wire s1770, sub1770, and1770, or1770;
  wire b_inv1770;
  assign b_inv1770 = ~b1770;
  assign s1770  = a1770 ^ b1770 ^ c1770;
  assign sub1770 = a1770 ^ b_inv1770 ^ c1770;
  assign and1770 = a1770 & b1770;
  assign or1770  = a1770 | b1770;
  assign c1771 = (a1770 & b1770) | (a1770 & c1770) | (b1770 & c1770);
  wire c_sub1771;
  assign c_sub1771 = (a1770 & b_inv1770) | (a1770 & c1770) | (b_inv1770 & c1770);
  wire s1771, sub1771, and1771, or1771;
  wire b_inv1771;
  assign b_inv1771 = ~b1771;
  assign s1771  = a1771 ^ b1771 ^ c1771;
  assign sub1771 = a1771 ^ b_inv1771 ^ c1771;
  assign and1771 = a1771 & b1771;
  assign or1771  = a1771 | b1771;
  assign c1772 = (a1771 & b1771) | (a1771 & c1771) | (b1771 & c1771);
  wire c_sub1772;
  assign c_sub1772 = (a1771 & b_inv1771) | (a1771 & c1771) | (b_inv1771 & c1771);
  wire s1772, sub1772, and1772, or1772;
  wire b_inv1772;
  assign b_inv1772 = ~b1772;
  assign s1772  = a1772 ^ b1772 ^ c1772;
  assign sub1772 = a1772 ^ b_inv1772 ^ c1772;
  assign and1772 = a1772 & b1772;
  assign or1772  = a1772 | b1772;
  assign c1773 = (a1772 & b1772) | (a1772 & c1772) | (b1772 & c1772);
  wire c_sub1773;
  assign c_sub1773 = (a1772 & b_inv1772) | (a1772 & c1772) | (b_inv1772 & c1772);
  wire s1773, sub1773, and1773, or1773;
  wire b_inv1773;
  assign b_inv1773 = ~b1773;
  assign s1773  = a1773 ^ b1773 ^ c1773;
  assign sub1773 = a1773 ^ b_inv1773 ^ c1773;
  assign and1773 = a1773 & b1773;
  assign or1773  = a1773 | b1773;
  assign c1774 = (a1773 & b1773) | (a1773 & c1773) | (b1773 & c1773);
  wire c_sub1774;
  assign c_sub1774 = (a1773 & b_inv1773) | (a1773 & c1773) | (b_inv1773 & c1773);
  wire s1774, sub1774, and1774, or1774;
  wire b_inv1774;
  assign b_inv1774 = ~b1774;
  assign s1774  = a1774 ^ b1774 ^ c1774;
  assign sub1774 = a1774 ^ b_inv1774 ^ c1774;
  assign and1774 = a1774 & b1774;
  assign or1774  = a1774 | b1774;
  assign c1775 = (a1774 & b1774) | (a1774 & c1774) | (b1774 & c1774);
  wire c_sub1775;
  assign c_sub1775 = (a1774 & b_inv1774) | (a1774 & c1774) | (b_inv1774 & c1774);
  wire s1775, sub1775, and1775, or1775;
  wire b_inv1775;
  assign b_inv1775 = ~b1775;
  assign s1775  = a1775 ^ b1775 ^ c1775;
  assign sub1775 = a1775 ^ b_inv1775 ^ c1775;
  assign and1775 = a1775 & b1775;
  assign or1775  = a1775 | b1775;
  assign c1776 = (a1775 & b1775) | (a1775 & c1775) | (b1775 & c1775);
  wire c_sub1776;
  assign c_sub1776 = (a1775 & b_inv1775) | (a1775 & c1775) | (b_inv1775 & c1775);
  wire s1776, sub1776, and1776, or1776;
  wire b_inv1776;
  assign b_inv1776 = ~b1776;
  assign s1776  = a1776 ^ b1776 ^ c1776;
  assign sub1776 = a1776 ^ b_inv1776 ^ c1776;
  assign and1776 = a1776 & b1776;
  assign or1776  = a1776 | b1776;
  assign c1777 = (a1776 & b1776) | (a1776 & c1776) | (b1776 & c1776);
  wire c_sub1777;
  assign c_sub1777 = (a1776 & b_inv1776) | (a1776 & c1776) | (b_inv1776 & c1776);
  wire s1777, sub1777, and1777, or1777;
  wire b_inv1777;
  assign b_inv1777 = ~b1777;
  assign s1777  = a1777 ^ b1777 ^ c1777;
  assign sub1777 = a1777 ^ b_inv1777 ^ c1777;
  assign and1777 = a1777 & b1777;
  assign or1777  = a1777 | b1777;
  assign c1778 = (a1777 & b1777) | (a1777 & c1777) | (b1777 & c1777);
  wire c_sub1778;
  assign c_sub1778 = (a1777 & b_inv1777) | (a1777 & c1777) | (b_inv1777 & c1777);
  wire s1778, sub1778, and1778, or1778;
  wire b_inv1778;
  assign b_inv1778 = ~b1778;
  assign s1778  = a1778 ^ b1778 ^ c1778;
  assign sub1778 = a1778 ^ b_inv1778 ^ c1778;
  assign and1778 = a1778 & b1778;
  assign or1778  = a1778 | b1778;
  assign c1779 = (a1778 & b1778) | (a1778 & c1778) | (b1778 & c1778);
  wire c_sub1779;
  assign c_sub1779 = (a1778 & b_inv1778) | (a1778 & c1778) | (b_inv1778 & c1778);
  wire s1779, sub1779, and1779, or1779;
  wire b_inv1779;
  assign b_inv1779 = ~b1779;
  assign s1779  = a1779 ^ b1779 ^ c1779;
  assign sub1779 = a1779 ^ b_inv1779 ^ c1779;
  assign and1779 = a1779 & b1779;
  assign or1779  = a1779 | b1779;
  assign c1780 = (a1779 & b1779) | (a1779 & c1779) | (b1779 & c1779);
  wire c_sub1780;
  assign c_sub1780 = (a1779 & b_inv1779) | (a1779 & c1779) | (b_inv1779 & c1779);
  wire s1780, sub1780, and1780, or1780;
  wire b_inv1780;
  assign b_inv1780 = ~b1780;
  assign s1780  = a1780 ^ b1780 ^ c1780;
  assign sub1780 = a1780 ^ b_inv1780 ^ c1780;
  assign and1780 = a1780 & b1780;
  assign or1780  = a1780 | b1780;
  assign c1781 = (a1780 & b1780) | (a1780 & c1780) | (b1780 & c1780);
  wire c_sub1781;
  assign c_sub1781 = (a1780 & b_inv1780) | (a1780 & c1780) | (b_inv1780 & c1780);
  wire s1781, sub1781, and1781, or1781;
  wire b_inv1781;
  assign b_inv1781 = ~b1781;
  assign s1781  = a1781 ^ b1781 ^ c1781;
  assign sub1781 = a1781 ^ b_inv1781 ^ c1781;
  assign and1781 = a1781 & b1781;
  assign or1781  = a1781 | b1781;
  assign c1782 = (a1781 & b1781) | (a1781 & c1781) | (b1781 & c1781);
  wire c_sub1782;
  assign c_sub1782 = (a1781 & b_inv1781) | (a1781 & c1781) | (b_inv1781 & c1781);
  wire s1782, sub1782, and1782, or1782;
  wire b_inv1782;
  assign b_inv1782 = ~b1782;
  assign s1782  = a1782 ^ b1782 ^ c1782;
  assign sub1782 = a1782 ^ b_inv1782 ^ c1782;
  assign and1782 = a1782 & b1782;
  assign or1782  = a1782 | b1782;
  assign c1783 = (a1782 & b1782) | (a1782 & c1782) | (b1782 & c1782);
  wire c_sub1783;
  assign c_sub1783 = (a1782 & b_inv1782) | (a1782 & c1782) | (b_inv1782 & c1782);
  wire s1783, sub1783, and1783, or1783;
  wire b_inv1783;
  assign b_inv1783 = ~b1783;
  assign s1783  = a1783 ^ b1783 ^ c1783;
  assign sub1783 = a1783 ^ b_inv1783 ^ c1783;
  assign and1783 = a1783 & b1783;
  assign or1783  = a1783 | b1783;
  assign c1784 = (a1783 & b1783) | (a1783 & c1783) | (b1783 & c1783);
  wire c_sub1784;
  assign c_sub1784 = (a1783 & b_inv1783) | (a1783 & c1783) | (b_inv1783 & c1783);
  wire s1784, sub1784, and1784, or1784;
  wire b_inv1784;
  assign b_inv1784 = ~b1784;
  assign s1784  = a1784 ^ b1784 ^ c1784;
  assign sub1784 = a1784 ^ b_inv1784 ^ c1784;
  assign and1784 = a1784 & b1784;
  assign or1784  = a1784 | b1784;
  assign c1785 = (a1784 & b1784) | (a1784 & c1784) | (b1784 & c1784);
  wire c_sub1785;
  assign c_sub1785 = (a1784 & b_inv1784) | (a1784 & c1784) | (b_inv1784 & c1784);
  wire s1785, sub1785, and1785, or1785;
  wire b_inv1785;
  assign b_inv1785 = ~b1785;
  assign s1785  = a1785 ^ b1785 ^ c1785;
  assign sub1785 = a1785 ^ b_inv1785 ^ c1785;
  assign and1785 = a1785 & b1785;
  assign or1785  = a1785 | b1785;
  assign c1786 = (a1785 & b1785) | (a1785 & c1785) | (b1785 & c1785);
  wire c_sub1786;
  assign c_sub1786 = (a1785 & b_inv1785) | (a1785 & c1785) | (b_inv1785 & c1785);
  wire s1786, sub1786, and1786, or1786;
  wire b_inv1786;
  assign b_inv1786 = ~b1786;
  assign s1786  = a1786 ^ b1786 ^ c1786;
  assign sub1786 = a1786 ^ b_inv1786 ^ c1786;
  assign and1786 = a1786 & b1786;
  assign or1786  = a1786 | b1786;
  assign c1787 = (a1786 & b1786) | (a1786 & c1786) | (b1786 & c1786);
  wire c_sub1787;
  assign c_sub1787 = (a1786 & b_inv1786) | (a1786 & c1786) | (b_inv1786 & c1786);
  wire s1787, sub1787, and1787, or1787;
  wire b_inv1787;
  assign b_inv1787 = ~b1787;
  assign s1787  = a1787 ^ b1787 ^ c1787;
  assign sub1787 = a1787 ^ b_inv1787 ^ c1787;
  assign and1787 = a1787 & b1787;
  assign or1787  = a1787 | b1787;
  assign c1788 = (a1787 & b1787) | (a1787 & c1787) | (b1787 & c1787);
  wire c_sub1788;
  assign c_sub1788 = (a1787 & b_inv1787) | (a1787 & c1787) | (b_inv1787 & c1787);
  wire s1788, sub1788, and1788, or1788;
  wire b_inv1788;
  assign b_inv1788 = ~b1788;
  assign s1788  = a1788 ^ b1788 ^ c1788;
  assign sub1788 = a1788 ^ b_inv1788 ^ c1788;
  assign and1788 = a1788 & b1788;
  assign or1788  = a1788 | b1788;
  assign c1789 = (a1788 & b1788) | (a1788 & c1788) | (b1788 & c1788);
  wire c_sub1789;
  assign c_sub1789 = (a1788 & b_inv1788) | (a1788 & c1788) | (b_inv1788 & c1788);
  wire s1789, sub1789, and1789, or1789;
  wire b_inv1789;
  assign b_inv1789 = ~b1789;
  assign s1789  = a1789 ^ b1789 ^ c1789;
  assign sub1789 = a1789 ^ b_inv1789 ^ c1789;
  assign and1789 = a1789 & b1789;
  assign or1789  = a1789 | b1789;
  assign c1790 = (a1789 & b1789) | (a1789 & c1789) | (b1789 & c1789);
  wire c_sub1790;
  assign c_sub1790 = (a1789 & b_inv1789) | (a1789 & c1789) | (b_inv1789 & c1789);
  wire s1790, sub1790, and1790, or1790;
  wire b_inv1790;
  assign b_inv1790 = ~b1790;
  assign s1790  = a1790 ^ b1790 ^ c1790;
  assign sub1790 = a1790 ^ b_inv1790 ^ c1790;
  assign and1790 = a1790 & b1790;
  assign or1790  = a1790 | b1790;
  assign c1791 = (a1790 & b1790) | (a1790 & c1790) | (b1790 & c1790);
  wire c_sub1791;
  assign c_sub1791 = (a1790 & b_inv1790) | (a1790 & c1790) | (b_inv1790 & c1790);
  wire s1791, sub1791, and1791, or1791;
  wire b_inv1791;
  assign b_inv1791 = ~b1791;
  assign s1791  = a1791 ^ b1791 ^ c1791;
  assign sub1791 = a1791 ^ b_inv1791 ^ c1791;
  assign and1791 = a1791 & b1791;
  assign or1791  = a1791 | b1791;
  assign c1792 = (a1791 & b1791) | (a1791 & c1791) | (b1791 & c1791);
  wire c_sub1792;
  assign c_sub1792 = (a1791 & b_inv1791) | (a1791 & c1791) | (b_inv1791 & c1791);
  wire s1792, sub1792, and1792, or1792;
  wire b_inv1792;
  assign b_inv1792 = ~b1792;
  assign s1792  = a1792 ^ b1792 ^ c1792;
  assign sub1792 = a1792 ^ b_inv1792 ^ c1792;
  assign and1792 = a1792 & b1792;
  assign or1792  = a1792 | b1792;
  assign c1793 = (a1792 & b1792) | (a1792 & c1792) | (b1792 & c1792);
  wire c_sub1793;
  assign c_sub1793 = (a1792 & b_inv1792) | (a1792 & c1792) | (b_inv1792 & c1792);
  wire s1793, sub1793, and1793, or1793;
  wire b_inv1793;
  assign b_inv1793 = ~b1793;
  assign s1793  = a1793 ^ b1793 ^ c1793;
  assign sub1793 = a1793 ^ b_inv1793 ^ c1793;
  assign and1793 = a1793 & b1793;
  assign or1793  = a1793 | b1793;
  assign c1794 = (a1793 & b1793) | (a1793 & c1793) | (b1793 & c1793);
  wire c_sub1794;
  assign c_sub1794 = (a1793 & b_inv1793) | (a1793 & c1793) | (b_inv1793 & c1793);
  wire s1794, sub1794, and1794, or1794;
  wire b_inv1794;
  assign b_inv1794 = ~b1794;
  assign s1794  = a1794 ^ b1794 ^ c1794;
  assign sub1794 = a1794 ^ b_inv1794 ^ c1794;
  assign and1794 = a1794 & b1794;
  assign or1794  = a1794 | b1794;
  assign c1795 = (a1794 & b1794) | (a1794 & c1794) | (b1794 & c1794);
  wire c_sub1795;
  assign c_sub1795 = (a1794 & b_inv1794) | (a1794 & c1794) | (b_inv1794 & c1794);
  wire s1795, sub1795, and1795, or1795;
  wire b_inv1795;
  assign b_inv1795 = ~b1795;
  assign s1795  = a1795 ^ b1795 ^ c1795;
  assign sub1795 = a1795 ^ b_inv1795 ^ c1795;
  assign and1795 = a1795 & b1795;
  assign or1795  = a1795 | b1795;
  assign c1796 = (a1795 & b1795) | (a1795 & c1795) | (b1795 & c1795);
  wire c_sub1796;
  assign c_sub1796 = (a1795 & b_inv1795) | (a1795 & c1795) | (b_inv1795 & c1795);
  wire s1796, sub1796, and1796, or1796;
  wire b_inv1796;
  assign b_inv1796 = ~b1796;
  assign s1796  = a1796 ^ b1796 ^ c1796;
  assign sub1796 = a1796 ^ b_inv1796 ^ c1796;
  assign and1796 = a1796 & b1796;
  assign or1796  = a1796 | b1796;
  assign c1797 = (a1796 & b1796) | (a1796 & c1796) | (b1796 & c1796);
  wire c_sub1797;
  assign c_sub1797 = (a1796 & b_inv1796) | (a1796 & c1796) | (b_inv1796 & c1796);
  wire s1797, sub1797, and1797, or1797;
  wire b_inv1797;
  assign b_inv1797 = ~b1797;
  assign s1797  = a1797 ^ b1797 ^ c1797;
  assign sub1797 = a1797 ^ b_inv1797 ^ c1797;
  assign and1797 = a1797 & b1797;
  assign or1797  = a1797 | b1797;
  assign c1798 = (a1797 & b1797) | (a1797 & c1797) | (b1797 & c1797);
  wire c_sub1798;
  assign c_sub1798 = (a1797 & b_inv1797) | (a1797 & c1797) | (b_inv1797 & c1797);
  wire s1798, sub1798, and1798, or1798;
  wire b_inv1798;
  assign b_inv1798 = ~b1798;
  assign s1798  = a1798 ^ b1798 ^ c1798;
  assign sub1798 = a1798 ^ b_inv1798 ^ c1798;
  assign and1798 = a1798 & b1798;
  assign or1798  = a1798 | b1798;
  assign c1799 = (a1798 & b1798) | (a1798 & c1798) | (b1798 & c1798);
  wire c_sub1799;
  assign c_sub1799 = (a1798 & b_inv1798) | (a1798 & c1798) | (b_inv1798 & c1798);
  wire s1799, sub1799, and1799, or1799;
  wire b_inv1799;
  assign b_inv1799 = ~b1799;
  assign s1799  = a1799 ^ b1799 ^ c1799;
  assign sub1799 = a1799 ^ b_inv1799 ^ c1799;
  assign and1799 = a1799 & b1799;
  assign or1799  = a1799 | b1799;
  assign c1800 = (a1799 & b1799) | (a1799 & c1799) | (b1799 & c1799);
  wire c_sub1800;
  assign c_sub1800 = (a1799 & b_inv1799) | (a1799 & c1799) | (b_inv1799 & c1799);
  wire s1800, sub1800, and1800, or1800;
  wire b_inv1800;
  assign b_inv1800 = ~b1800;
  assign s1800  = a1800 ^ b1800 ^ c1800;
  assign sub1800 = a1800 ^ b_inv1800 ^ c1800;
  assign and1800 = a1800 & b1800;
  assign or1800  = a1800 | b1800;
  assign c1801 = (a1800 & b1800) | (a1800 & c1800) | (b1800 & c1800);
  wire c_sub1801;
  assign c_sub1801 = (a1800 & b_inv1800) | (a1800 & c1800) | (b_inv1800 & c1800);
  wire s1801, sub1801, and1801, or1801;
  wire b_inv1801;
  assign b_inv1801 = ~b1801;
  assign s1801  = a1801 ^ b1801 ^ c1801;
  assign sub1801 = a1801 ^ b_inv1801 ^ c1801;
  assign and1801 = a1801 & b1801;
  assign or1801  = a1801 | b1801;
  assign c1802 = (a1801 & b1801) | (a1801 & c1801) | (b1801 & c1801);
  wire c_sub1802;
  assign c_sub1802 = (a1801 & b_inv1801) | (a1801 & c1801) | (b_inv1801 & c1801);
  wire s1802, sub1802, and1802, or1802;
  wire b_inv1802;
  assign b_inv1802 = ~b1802;
  assign s1802  = a1802 ^ b1802 ^ c1802;
  assign sub1802 = a1802 ^ b_inv1802 ^ c1802;
  assign and1802 = a1802 & b1802;
  assign or1802  = a1802 | b1802;
  assign c1803 = (a1802 & b1802) | (a1802 & c1802) | (b1802 & c1802);
  wire c_sub1803;
  assign c_sub1803 = (a1802 & b_inv1802) | (a1802 & c1802) | (b_inv1802 & c1802);
  wire s1803, sub1803, and1803, or1803;
  wire b_inv1803;
  assign b_inv1803 = ~b1803;
  assign s1803  = a1803 ^ b1803 ^ c1803;
  assign sub1803 = a1803 ^ b_inv1803 ^ c1803;
  assign and1803 = a1803 & b1803;
  assign or1803  = a1803 | b1803;
  assign c1804 = (a1803 & b1803) | (a1803 & c1803) | (b1803 & c1803);
  wire c_sub1804;
  assign c_sub1804 = (a1803 & b_inv1803) | (a1803 & c1803) | (b_inv1803 & c1803);
  wire s1804, sub1804, and1804, or1804;
  wire b_inv1804;
  assign b_inv1804 = ~b1804;
  assign s1804  = a1804 ^ b1804 ^ c1804;
  assign sub1804 = a1804 ^ b_inv1804 ^ c1804;
  assign and1804 = a1804 & b1804;
  assign or1804  = a1804 | b1804;
  assign c1805 = (a1804 & b1804) | (a1804 & c1804) | (b1804 & c1804);
  wire c_sub1805;
  assign c_sub1805 = (a1804 & b_inv1804) | (a1804 & c1804) | (b_inv1804 & c1804);
  wire s1805, sub1805, and1805, or1805;
  wire b_inv1805;
  assign b_inv1805 = ~b1805;
  assign s1805  = a1805 ^ b1805 ^ c1805;
  assign sub1805 = a1805 ^ b_inv1805 ^ c1805;
  assign and1805 = a1805 & b1805;
  assign or1805  = a1805 | b1805;
  assign c1806 = (a1805 & b1805) | (a1805 & c1805) | (b1805 & c1805);
  wire c_sub1806;
  assign c_sub1806 = (a1805 & b_inv1805) | (a1805 & c1805) | (b_inv1805 & c1805);
  wire s1806, sub1806, and1806, or1806;
  wire b_inv1806;
  assign b_inv1806 = ~b1806;
  assign s1806  = a1806 ^ b1806 ^ c1806;
  assign sub1806 = a1806 ^ b_inv1806 ^ c1806;
  assign and1806 = a1806 & b1806;
  assign or1806  = a1806 | b1806;
  assign c1807 = (a1806 & b1806) | (a1806 & c1806) | (b1806 & c1806);
  wire c_sub1807;
  assign c_sub1807 = (a1806 & b_inv1806) | (a1806 & c1806) | (b_inv1806 & c1806);
  wire s1807, sub1807, and1807, or1807;
  wire b_inv1807;
  assign b_inv1807 = ~b1807;
  assign s1807  = a1807 ^ b1807 ^ c1807;
  assign sub1807 = a1807 ^ b_inv1807 ^ c1807;
  assign and1807 = a1807 & b1807;
  assign or1807  = a1807 | b1807;
  assign c1808 = (a1807 & b1807) | (a1807 & c1807) | (b1807 & c1807);
  wire c_sub1808;
  assign c_sub1808 = (a1807 & b_inv1807) | (a1807 & c1807) | (b_inv1807 & c1807);
  wire s1808, sub1808, and1808, or1808;
  wire b_inv1808;
  assign b_inv1808 = ~b1808;
  assign s1808  = a1808 ^ b1808 ^ c1808;
  assign sub1808 = a1808 ^ b_inv1808 ^ c1808;
  assign and1808 = a1808 & b1808;
  assign or1808  = a1808 | b1808;
  assign c1809 = (a1808 & b1808) | (a1808 & c1808) | (b1808 & c1808);
  wire c_sub1809;
  assign c_sub1809 = (a1808 & b_inv1808) | (a1808 & c1808) | (b_inv1808 & c1808);
  wire s1809, sub1809, and1809, or1809;
  wire b_inv1809;
  assign b_inv1809 = ~b1809;
  assign s1809  = a1809 ^ b1809 ^ c1809;
  assign sub1809 = a1809 ^ b_inv1809 ^ c1809;
  assign and1809 = a1809 & b1809;
  assign or1809  = a1809 | b1809;
  assign c1810 = (a1809 & b1809) | (a1809 & c1809) | (b1809 & c1809);
  wire c_sub1810;
  assign c_sub1810 = (a1809 & b_inv1809) | (a1809 & c1809) | (b_inv1809 & c1809);
  wire s1810, sub1810, and1810, or1810;
  wire b_inv1810;
  assign b_inv1810 = ~b1810;
  assign s1810  = a1810 ^ b1810 ^ c1810;
  assign sub1810 = a1810 ^ b_inv1810 ^ c1810;
  assign and1810 = a1810 & b1810;
  assign or1810  = a1810 | b1810;
  assign c1811 = (a1810 & b1810) | (a1810 & c1810) | (b1810 & c1810);
  wire c_sub1811;
  assign c_sub1811 = (a1810 & b_inv1810) | (a1810 & c1810) | (b_inv1810 & c1810);
  wire s1811, sub1811, and1811, or1811;
  wire b_inv1811;
  assign b_inv1811 = ~b1811;
  assign s1811  = a1811 ^ b1811 ^ c1811;
  assign sub1811 = a1811 ^ b_inv1811 ^ c1811;
  assign and1811 = a1811 & b1811;
  assign or1811  = a1811 | b1811;
  assign c1812 = (a1811 & b1811) | (a1811 & c1811) | (b1811 & c1811);
  wire c_sub1812;
  assign c_sub1812 = (a1811 & b_inv1811) | (a1811 & c1811) | (b_inv1811 & c1811);
  wire s1812, sub1812, and1812, or1812;
  wire b_inv1812;
  assign b_inv1812 = ~b1812;
  assign s1812  = a1812 ^ b1812 ^ c1812;
  assign sub1812 = a1812 ^ b_inv1812 ^ c1812;
  assign and1812 = a1812 & b1812;
  assign or1812  = a1812 | b1812;
  assign c1813 = (a1812 & b1812) | (a1812 & c1812) | (b1812 & c1812);
  wire c_sub1813;
  assign c_sub1813 = (a1812 & b_inv1812) | (a1812 & c1812) | (b_inv1812 & c1812);
  wire s1813, sub1813, and1813, or1813;
  wire b_inv1813;
  assign b_inv1813 = ~b1813;
  assign s1813  = a1813 ^ b1813 ^ c1813;
  assign sub1813 = a1813 ^ b_inv1813 ^ c1813;
  assign and1813 = a1813 & b1813;
  assign or1813  = a1813 | b1813;
  assign c1814 = (a1813 & b1813) | (a1813 & c1813) | (b1813 & c1813);
  wire c_sub1814;
  assign c_sub1814 = (a1813 & b_inv1813) | (a1813 & c1813) | (b_inv1813 & c1813);
  wire s1814, sub1814, and1814, or1814;
  wire b_inv1814;
  assign b_inv1814 = ~b1814;
  assign s1814  = a1814 ^ b1814 ^ c1814;
  assign sub1814 = a1814 ^ b_inv1814 ^ c1814;
  assign and1814 = a1814 & b1814;
  assign or1814  = a1814 | b1814;
  assign c1815 = (a1814 & b1814) | (a1814 & c1814) | (b1814 & c1814);
  wire c_sub1815;
  assign c_sub1815 = (a1814 & b_inv1814) | (a1814 & c1814) | (b_inv1814 & c1814);
  wire s1815, sub1815, and1815, or1815;
  wire b_inv1815;
  assign b_inv1815 = ~b1815;
  assign s1815  = a1815 ^ b1815 ^ c1815;
  assign sub1815 = a1815 ^ b_inv1815 ^ c1815;
  assign and1815 = a1815 & b1815;
  assign or1815  = a1815 | b1815;
  assign c1816 = (a1815 & b1815) | (a1815 & c1815) | (b1815 & c1815);
  wire c_sub1816;
  assign c_sub1816 = (a1815 & b_inv1815) | (a1815 & c1815) | (b_inv1815 & c1815);
  wire s1816, sub1816, and1816, or1816;
  wire b_inv1816;
  assign b_inv1816 = ~b1816;
  assign s1816  = a1816 ^ b1816 ^ c1816;
  assign sub1816 = a1816 ^ b_inv1816 ^ c1816;
  assign and1816 = a1816 & b1816;
  assign or1816  = a1816 | b1816;
  assign c1817 = (a1816 & b1816) | (a1816 & c1816) | (b1816 & c1816);
  wire c_sub1817;
  assign c_sub1817 = (a1816 & b_inv1816) | (a1816 & c1816) | (b_inv1816 & c1816);
  wire s1817, sub1817, and1817, or1817;
  wire b_inv1817;
  assign b_inv1817 = ~b1817;
  assign s1817  = a1817 ^ b1817 ^ c1817;
  assign sub1817 = a1817 ^ b_inv1817 ^ c1817;
  assign and1817 = a1817 & b1817;
  assign or1817  = a1817 | b1817;
  assign c1818 = (a1817 & b1817) | (a1817 & c1817) | (b1817 & c1817);
  wire c_sub1818;
  assign c_sub1818 = (a1817 & b_inv1817) | (a1817 & c1817) | (b_inv1817 & c1817);
  wire s1818, sub1818, and1818, or1818;
  wire b_inv1818;
  assign b_inv1818 = ~b1818;
  assign s1818  = a1818 ^ b1818 ^ c1818;
  assign sub1818 = a1818 ^ b_inv1818 ^ c1818;
  assign and1818 = a1818 & b1818;
  assign or1818  = a1818 | b1818;
  assign c1819 = (a1818 & b1818) | (a1818 & c1818) | (b1818 & c1818);
  wire c_sub1819;
  assign c_sub1819 = (a1818 & b_inv1818) | (a1818 & c1818) | (b_inv1818 & c1818);
  wire s1819, sub1819, and1819, or1819;
  wire b_inv1819;
  assign b_inv1819 = ~b1819;
  assign s1819  = a1819 ^ b1819 ^ c1819;
  assign sub1819 = a1819 ^ b_inv1819 ^ c1819;
  assign and1819 = a1819 & b1819;
  assign or1819  = a1819 | b1819;
  assign c1820 = (a1819 & b1819) | (a1819 & c1819) | (b1819 & c1819);
  wire c_sub1820;
  assign c_sub1820 = (a1819 & b_inv1819) | (a1819 & c1819) | (b_inv1819 & c1819);
  wire s1820, sub1820, and1820, or1820;
  wire b_inv1820;
  assign b_inv1820 = ~b1820;
  assign s1820  = a1820 ^ b1820 ^ c1820;
  assign sub1820 = a1820 ^ b_inv1820 ^ c1820;
  assign and1820 = a1820 & b1820;
  assign or1820  = a1820 | b1820;
  assign c1821 = (a1820 & b1820) | (a1820 & c1820) | (b1820 & c1820);
  wire c_sub1821;
  assign c_sub1821 = (a1820 & b_inv1820) | (a1820 & c1820) | (b_inv1820 & c1820);
  wire s1821, sub1821, and1821, or1821;
  wire b_inv1821;
  assign b_inv1821 = ~b1821;
  assign s1821  = a1821 ^ b1821 ^ c1821;
  assign sub1821 = a1821 ^ b_inv1821 ^ c1821;
  assign and1821 = a1821 & b1821;
  assign or1821  = a1821 | b1821;
  assign c1822 = (a1821 & b1821) | (a1821 & c1821) | (b1821 & c1821);
  wire c_sub1822;
  assign c_sub1822 = (a1821 & b_inv1821) | (a1821 & c1821) | (b_inv1821 & c1821);
  wire s1822, sub1822, and1822, or1822;
  wire b_inv1822;
  assign b_inv1822 = ~b1822;
  assign s1822  = a1822 ^ b1822 ^ c1822;
  assign sub1822 = a1822 ^ b_inv1822 ^ c1822;
  assign and1822 = a1822 & b1822;
  assign or1822  = a1822 | b1822;
  assign c1823 = (a1822 & b1822) | (a1822 & c1822) | (b1822 & c1822);
  wire c_sub1823;
  assign c_sub1823 = (a1822 & b_inv1822) | (a1822 & c1822) | (b_inv1822 & c1822);
  wire s1823, sub1823, and1823, or1823;
  wire b_inv1823;
  assign b_inv1823 = ~b1823;
  assign s1823  = a1823 ^ b1823 ^ c1823;
  assign sub1823 = a1823 ^ b_inv1823 ^ c1823;
  assign and1823 = a1823 & b1823;
  assign or1823  = a1823 | b1823;
  assign c1824 = (a1823 & b1823) | (a1823 & c1823) | (b1823 & c1823);
  wire c_sub1824;
  assign c_sub1824 = (a1823 & b_inv1823) | (a1823 & c1823) | (b_inv1823 & c1823);
  wire s1824, sub1824, and1824, or1824;
  wire b_inv1824;
  assign b_inv1824 = ~b1824;
  assign s1824  = a1824 ^ b1824 ^ c1824;
  assign sub1824 = a1824 ^ b_inv1824 ^ c1824;
  assign and1824 = a1824 & b1824;
  assign or1824  = a1824 | b1824;
  assign c1825 = (a1824 & b1824) | (a1824 & c1824) | (b1824 & c1824);
  wire c_sub1825;
  assign c_sub1825 = (a1824 & b_inv1824) | (a1824 & c1824) | (b_inv1824 & c1824);
  wire s1825, sub1825, and1825, or1825;
  wire b_inv1825;
  assign b_inv1825 = ~b1825;
  assign s1825  = a1825 ^ b1825 ^ c1825;
  assign sub1825 = a1825 ^ b_inv1825 ^ c1825;
  assign and1825 = a1825 & b1825;
  assign or1825  = a1825 | b1825;
  assign c1826 = (a1825 & b1825) | (a1825 & c1825) | (b1825 & c1825);
  wire c_sub1826;
  assign c_sub1826 = (a1825 & b_inv1825) | (a1825 & c1825) | (b_inv1825 & c1825);
  wire s1826, sub1826, and1826, or1826;
  wire b_inv1826;
  assign b_inv1826 = ~b1826;
  assign s1826  = a1826 ^ b1826 ^ c1826;
  assign sub1826 = a1826 ^ b_inv1826 ^ c1826;
  assign and1826 = a1826 & b1826;
  assign or1826  = a1826 | b1826;
  assign c1827 = (a1826 & b1826) | (a1826 & c1826) | (b1826 & c1826);
  wire c_sub1827;
  assign c_sub1827 = (a1826 & b_inv1826) | (a1826 & c1826) | (b_inv1826 & c1826);
  wire s1827, sub1827, and1827, or1827;
  wire b_inv1827;
  assign b_inv1827 = ~b1827;
  assign s1827  = a1827 ^ b1827 ^ c1827;
  assign sub1827 = a1827 ^ b_inv1827 ^ c1827;
  assign and1827 = a1827 & b1827;
  assign or1827  = a1827 | b1827;
  assign c1828 = (a1827 & b1827) | (a1827 & c1827) | (b1827 & c1827);
  wire c_sub1828;
  assign c_sub1828 = (a1827 & b_inv1827) | (a1827 & c1827) | (b_inv1827 & c1827);
  wire s1828, sub1828, and1828, or1828;
  wire b_inv1828;
  assign b_inv1828 = ~b1828;
  assign s1828  = a1828 ^ b1828 ^ c1828;
  assign sub1828 = a1828 ^ b_inv1828 ^ c1828;
  assign and1828 = a1828 & b1828;
  assign or1828  = a1828 | b1828;
  assign c1829 = (a1828 & b1828) | (a1828 & c1828) | (b1828 & c1828);
  wire c_sub1829;
  assign c_sub1829 = (a1828 & b_inv1828) | (a1828 & c1828) | (b_inv1828 & c1828);
  wire s1829, sub1829, and1829, or1829;
  wire b_inv1829;
  assign b_inv1829 = ~b1829;
  assign s1829  = a1829 ^ b1829 ^ c1829;
  assign sub1829 = a1829 ^ b_inv1829 ^ c1829;
  assign and1829 = a1829 & b1829;
  assign or1829  = a1829 | b1829;
  assign c1830 = (a1829 & b1829) | (a1829 & c1829) | (b1829 & c1829);
  wire c_sub1830;
  assign c_sub1830 = (a1829 & b_inv1829) | (a1829 & c1829) | (b_inv1829 & c1829);
  wire s1830, sub1830, and1830, or1830;
  wire b_inv1830;
  assign b_inv1830 = ~b1830;
  assign s1830  = a1830 ^ b1830 ^ c1830;
  assign sub1830 = a1830 ^ b_inv1830 ^ c1830;
  assign and1830 = a1830 & b1830;
  assign or1830  = a1830 | b1830;
  assign c1831 = (a1830 & b1830) | (a1830 & c1830) | (b1830 & c1830);
  wire c_sub1831;
  assign c_sub1831 = (a1830 & b_inv1830) | (a1830 & c1830) | (b_inv1830 & c1830);
  wire s1831, sub1831, and1831, or1831;
  wire b_inv1831;
  assign b_inv1831 = ~b1831;
  assign s1831  = a1831 ^ b1831 ^ c1831;
  assign sub1831 = a1831 ^ b_inv1831 ^ c1831;
  assign and1831 = a1831 & b1831;
  assign or1831  = a1831 | b1831;
  assign c1832 = (a1831 & b1831) | (a1831 & c1831) | (b1831 & c1831);
  wire c_sub1832;
  assign c_sub1832 = (a1831 & b_inv1831) | (a1831 & c1831) | (b_inv1831 & c1831);
  wire s1832, sub1832, and1832, or1832;
  wire b_inv1832;
  assign b_inv1832 = ~b1832;
  assign s1832  = a1832 ^ b1832 ^ c1832;
  assign sub1832 = a1832 ^ b_inv1832 ^ c1832;
  assign and1832 = a1832 & b1832;
  assign or1832  = a1832 | b1832;
  assign c1833 = (a1832 & b1832) | (a1832 & c1832) | (b1832 & c1832);
  wire c_sub1833;
  assign c_sub1833 = (a1832 & b_inv1832) | (a1832 & c1832) | (b_inv1832 & c1832);
  wire s1833, sub1833, and1833, or1833;
  wire b_inv1833;
  assign b_inv1833 = ~b1833;
  assign s1833  = a1833 ^ b1833 ^ c1833;
  assign sub1833 = a1833 ^ b_inv1833 ^ c1833;
  assign and1833 = a1833 & b1833;
  assign or1833  = a1833 | b1833;
  assign c1834 = (a1833 & b1833) | (a1833 & c1833) | (b1833 & c1833);
  wire c_sub1834;
  assign c_sub1834 = (a1833 & b_inv1833) | (a1833 & c1833) | (b_inv1833 & c1833);
  wire s1834, sub1834, and1834, or1834;
  wire b_inv1834;
  assign b_inv1834 = ~b1834;
  assign s1834  = a1834 ^ b1834 ^ c1834;
  assign sub1834 = a1834 ^ b_inv1834 ^ c1834;
  assign and1834 = a1834 & b1834;
  assign or1834  = a1834 | b1834;
  assign c1835 = (a1834 & b1834) | (a1834 & c1834) | (b1834 & c1834);
  wire c_sub1835;
  assign c_sub1835 = (a1834 & b_inv1834) | (a1834 & c1834) | (b_inv1834 & c1834);
  wire s1835, sub1835, and1835, or1835;
  wire b_inv1835;
  assign b_inv1835 = ~b1835;
  assign s1835  = a1835 ^ b1835 ^ c1835;
  assign sub1835 = a1835 ^ b_inv1835 ^ c1835;
  assign and1835 = a1835 & b1835;
  assign or1835  = a1835 | b1835;
  assign c1836 = (a1835 & b1835) | (a1835 & c1835) | (b1835 & c1835);
  wire c_sub1836;
  assign c_sub1836 = (a1835 & b_inv1835) | (a1835 & c1835) | (b_inv1835 & c1835);
  wire s1836, sub1836, and1836, or1836;
  wire b_inv1836;
  assign b_inv1836 = ~b1836;
  assign s1836  = a1836 ^ b1836 ^ c1836;
  assign sub1836 = a1836 ^ b_inv1836 ^ c1836;
  assign and1836 = a1836 & b1836;
  assign or1836  = a1836 | b1836;
  assign c1837 = (a1836 & b1836) | (a1836 & c1836) | (b1836 & c1836);
  wire c_sub1837;
  assign c_sub1837 = (a1836 & b_inv1836) | (a1836 & c1836) | (b_inv1836 & c1836);
  wire s1837, sub1837, and1837, or1837;
  wire b_inv1837;
  assign b_inv1837 = ~b1837;
  assign s1837  = a1837 ^ b1837 ^ c1837;
  assign sub1837 = a1837 ^ b_inv1837 ^ c1837;
  assign and1837 = a1837 & b1837;
  assign or1837  = a1837 | b1837;
  assign c1838 = (a1837 & b1837) | (a1837 & c1837) | (b1837 & c1837);
  wire c_sub1838;
  assign c_sub1838 = (a1837 & b_inv1837) | (a1837 & c1837) | (b_inv1837 & c1837);
  wire s1838, sub1838, and1838, or1838;
  wire b_inv1838;
  assign b_inv1838 = ~b1838;
  assign s1838  = a1838 ^ b1838 ^ c1838;
  assign sub1838 = a1838 ^ b_inv1838 ^ c1838;
  assign and1838 = a1838 & b1838;
  assign or1838  = a1838 | b1838;
  assign c1839 = (a1838 & b1838) | (a1838 & c1838) | (b1838 & c1838);
  wire c_sub1839;
  assign c_sub1839 = (a1838 & b_inv1838) | (a1838 & c1838) | (b_inv1838 & c1838);
  wire s1839, sub1839, and1839, or1839;
  wire b_inv1839;
  assign b_inv1839 = ~b1839;
  assign s1839  = a1839 ^ b1839 ^ c1839;
  assign sub1839 = a1839 ^ b_inv1839 ^ c1839;
  assign and1839 = a1839 & b1839;
  assign or1839  = a1839 | b1839;
  assign c1840 = (a1839 & b1839) | (a1839 & c1839) | (b1839 & c1839);
  wire c_sub1840;
  assign c_sub1840 = (a1839 & b_inv1839) | (a1839 & c1839) | (b_inv1839 & c1839);
  wire s1840, sub1840, and1840, or1840;
  wire b_inv1840;
  assign b_inv1840 = ~b1840;
  assign s1840  = a1840 ^ b1840 ^ c1840;
  assign sub1840 = a1840 ^ b_inv1840 ^ c1840;
  assign and1840 = a1840 & b1840;
  assign or1840  = a1840 | b1840;
  assign c1841 = (a1840 & b1840) | (a1840 & c1840) | (b1840 & c1840);
  wire c_sub1841;
  assign c_sub1841 = (a1840 & b_inv1840) | (a1840 & c1840) | (b_inv1840 & c1840);
  wire s1841, sub1841, and1841, or1841;
  wire b_inv1841;
  assign b_inv1841 = ~b1841;
  assign s1841  = a1841 ^ b1841 ^ c1841;
  assign sub1841 = a1841 ^ b_inv1841 ^ c1841;
  assign and1841 = a1841 & b1841;
  assign or1841  = a1841 | b1841;
  assign c1842 = (a1841 & b1841) | (a1841 & c1841) | (b1841 & c1841);
  wire c_sub1842;
  assign c_sub1842 = (a1841 & b_inv1841) | (a1841 & c1841) | (b_inv1841 & c1841);
  wire s1842, sub1842, and1842, or1842;
  wire b_inv1842;
  assign b_inv1842 = ~b1842;
  assign s1842  = a1842 ^ b1842 ^ c1842;
  assign sub1842 = a1842 ^ b_inv1842 ^ c1842;
  assign and1842 = a1842 & b1842;
  assign or1842  = a1842 | b1842;
  assign c1843 = (a1842 & b1842) | (a1842 & c1842) | (b1842 & c1842);
  wire c_sub1843;
  assign c_sub1843 = (a1842 & b_inv1842) | (a1842 & c1842) | (b_inv1842 & c1842);
  wire s1843, sub1843, and1843, or1843;
  wire b_inv1843;
  assign b_inv1843 = ~b1843;
  assign s1843  = a1843 ^ b1843 ^ c1843;
  assign sub1843 = a1843 ^ b_inv1843 ^ c1843;
  assign and1843 = a1843 & b1843;
  assign or1843  = a1843 | b1843;
  assign c1844 = (a1843 & b1843) | (a1843 & c1843) | (b1843 & c1843);
  wire c_sub1844;
  assign c_sub1844 = (a1843 & b_inv1843) | (a1843 & c1843) | (b_inv1843 & c1843);
  wire s1844, sub1844, and1844, or1844;
  wire b_inv1844;
  assign b_inv1844 = ~b1844;
  assign s1844  = a1844 ^ b1844 ^ c1844;
  assign sub1844 = a1844 ^ b_inv1844 ^ c1844;
  assign and1844 = a1844 & b1844;
  assign or1844  = a1844 | b1844;
  assign c1845 = (a1844 & b1844) | (a1844 & c1844) | (b1844 & c1844);
  wire c_sub1845;
  assign c_sub1845 = (a1844 & b_inv1844) | (a1844 & c1844) | (b_inv1844 & c1844);
  wire s1845, sub1845, and1845, or1845;
  wire b_inv1845;
  assign b_inv1845 = ~b1845;
  assign s1845  = a1845 ^ b1845 ^ c1845;
  assign sub1845 = a1845 ^ b_inv1845 ^ c1845;
  assign and1845 = a1845 & b1845;
  assign or1845  = a1845 | b1845;
  assign c1846 = (a1845 & b1845) | (a1845 & c1845) | (b1845 & c1845);
  wire c_sub1846;
  assign c_sub1846 = (a1845 & b_inv1845) | (a1845 & c1845) | (b_inv1845 & c1845);
  wire s1846, sub1846, and1846, or1846;
  wire b_inv1846;
  assign b_inv1846 = ~b1846;
  assign s1846  = a1846 ^ b1846 ^ c1846;
  assign sub1846 = a1846 ^ b_inv1846 ^ c1846;
  assign and1846 = a1846 & b1846;
  assign or1846  = a1846 | b1846;
  assign c1847 = (a1846 & b1846) | (a1846 & c1846) | (b1846 & c1846);
  wire c_sub1847;
  assign c_sub1847 = (a1846 & b_inv1846) | (a1846 & c1846) | (b_inv1846 & c1846);
  wire s1847, sub1847, and1847, or1847;
  wire b_inv1847;
  assign b_inv1847 = ~b1847;
  assign s1847  = a1847 ^ b1847 ^ c1847;
  assign sub1847 = a1847 ^ b_inv1847 ^ c1847;
  assign and1847 = a1847 & b1847;
  assign or1847  = a1847 | b1847;
  assign c1848 = (a1847 & b1847) | (a1847 & c1847) | (b1847 & c1847);
  wire c_sub1848;
  assign c_sub1848 = (a1847 & b_inv1847) | (a1847 & c1847) | (b_inv1847 & c1847);
  wire s1848, sub1848, and1848, or1848;
  wire b_inv1848;
  assign b_inv1848 = ~b1848;
  assign s1848  = a1848 ^ b1848 ^ c1848;
  assign sub1848 = a1848 ^ b_inv1848 ^ c1848;
  assign and1848 = a1848 & b1848;
  assign or1848  = a1848 | b1848;
  assign c1849 = (a1848 & b1848) | (a1848 & c1848) | (b1848 & c1848);
  wire c_sub1849;
  assign c_sub1849 = (a1848 & b_inv1848) | (a1848 & c1848) | (b_inv1848 & c1848);
  wire s1849, sub1849, and1849, or1849;
  wire b_inv1849;
  assign b_inv1849 = ~b1849;
  assign s1849  = a1849 ^ b1849 ^ c1849;
  assign sub1849 = a1849 ^ b_inv1849 ^ c1849;
  assign and1849 = a1849 & b1849;
  assign or1849  = a1849 | b1849;
  assign c1850 = (a1849 & b1849) | (a1849 & c1849) | (b1849 & c1849);
  wire c_sub1850;
  assign c_sub1850 = (a1849 & b_inv1849) | (a1849 & c1849) | (b_inv1849 & c1849);
  wire s1850, sub1850, and1850, or1850;
  wire b_inv1850;
  assign b_inv1850 = ~b1850;
  assign s1850  = a1850 ^ b1850 ^ c1850;
  assign sub1850 = a1850 ^ b_inv1850 ^ c1850;
  assign and1850 = a1850 & b1850;
  assign or1850  = a1850 | b1850;
  assign c1851 = (a1850 & b1850) | (a1850 & c1850) | (b1850 & c1850);
  wire c_sub1851;
  assign c_sub1851 = (a1850 & b_inv1850) | (a1850 & c1850) | (b_inv1850 & c1850);
  wire s1851, sub1851, and1851, or1851;
  wire b_inv1851;
  assign b_inv1851 = ~b1851;
  assign s1851  = a1851 ^ b1851 ^ c1851;
  assign sub1851 = a1851 ^ b_inv1851 ^ c1851;
  assign and1851 = a1851 & b1851;
  assign or1851  = a1851 | b1851;
  assign c1852 = (a1851 & b1851) | (a1851 & c1851) | (b1851 & c1851);
  wire c_sub1852;
  assign c_sub1852 = (a1851 & b_inv1851) | (a1851 & c1851) | (b_inv1851 & c1851);
  wire s1852, sub1852, and1852, or1852;
  wire b_inv1852;
  assign b_inv1852 = ~b1852;
  assign s1852  = a1852 ^ b1852 ^ c1852;
  assign sub1852 = a1852 ^ b_inv1852 ^ c1852;
  assign and1852 = a1852 & b1852;
  assign or1852  = a1852 | b1852;
  assign c1853 = (a1852 & b1852) | (a1852 & c1852) | (b1852 & c1852);
  wire c_sub1853;
  assign c_sub1853 = (a1852 & b_inv1852) | (a1852 & c1852) | (b_inv1852 & c1852);
  wire s1853, sub1853, and1853, or1853;
  wire b_inv1853;
  assign b_inv1853 = ~b1853;
  assign s1853  = a1853 ^ b1853 ^ c1853;
  assign sub1853 = a1853 ^ b_inv1853 ^ c1853;
  assign and1853 = a1853 & b1853;
  assign or1853  = a1853 | b1853;
  assign c1854 = (a1853 & b1853) | (a1853 & c1853) | (b1853 & c1853);
  wire c_sub1854;
  assign c_sub1854 = (a1853 & b_inv1853) | (a1853 & c1853) | (b_inv1853 & c1853);
  wire s1854, sub1854, and1854, or1854;
  wire b_inv1854;
  assign b_inv1854 = ~b1854;
  assign s1854  = a1854 ^ b1854 ^ c1854;
  assign sub1854 = a1854 ^ b_inv1854 ^ c1854;
  assign and1854 = a1854 & b1854;
  assign or1854  = a1854 | b1854;
  assign c1855 = (a1854 & b1854) | (a1854 & c1854) | (b1854 & c1854);
  wire c_sub1855;
  assign c_sub1855 = (a1854 & b_inv1854) | (a1854 & c1854) | (b_inv1854 & c1854);
  wire s1855, sub1855, and1855, or1855;
  wire b_inv1855;
  assign b_inv1855 = ~b1855;
  assign s1855  = a1855 ^ b1855 ^ c1855;
  assign sub1855 = a1855 ^ b_inv1855 ^ c1855;
  assign and1855 = a1855 & b1855;
  assign or1855  = a1855 | b1855;
  assign c1856 = (a1855 & b1855) | (a1855 & c1855) | (b1855 & c1855);
  wire c_sub1856;
  assign c_sub1856 = (a1855 & b_inv1855) | (a1855 & c1855) | (b_inv1855 & c1855);
  wire s1856, sub1856, and1856, or1856;
  wire b_inv1856;
  assign b_inv1856 = ~b1856;
  assign s1856  = a1856 ^ b1856 ^ c1856;
  assign sub1856 = a1856 ^ b_inv1856 ^ c1856;
  assign and1856 = a1856 & b1856;
  assign or1856  = a1856 | b1856;
  assign c1857 = (a1856 & b1856) | (a1856 & c1856) | (b1856 & c1856);
  wire c_sub1857;
  assign c_sub1857 = (a1856 & b_inv1856) | (a1856 & c1856) | (b_inv1856 & c1856);
  wire s1857, sub1857, and1857, or1857;
  wire b_inv1857;
  assign b_inv1857 = ~b1857;
  assign s1857  = a1857 ^ b1857 ^ c1857;
  assign sub1857 = a1857 ^ b_inv1857 ^ c1857;
  assign and1857 = a1857 & b1857;
  assign or1857  = a1857 | b1857;
  assign c1858 = (a1857 & b1857) | (a1857 & c1857) | (b1857 & c1857);
  wire c_sub1858;
  assign c_sub1858 = (a1857 & b_inv1857) | (a1857 & c1857) | (b_inv1857 & c1857);
  wire s1858, sub1858, and1858, or1858;
  wire b_inv1858;
  assign b_inv1858 = ~b1858;
  assign s1858  = a1858 ^ b1858 ^ c1858;
  assign sub1858 = a1858 ^ b_inv1858 ^ c1858;
  assign and1858 = a1858 & b1858;
  assign or1858  = a1858 | b1858;
  assign c1859 = (a1858 & b1858) | (a1858 & c1858) | (b1858 & c1858);
  wire c_sub1859;
  assign c_sub1859 = (a1858 & b_inv1858) | (a1858 & c1858) | (b_inv1858 & c1858);
  wire s1859, sub1859, and1859, or1859;
  wire b_inv1859;
  assign b_inv1859 = ~b1859;
  assign s1859  = a1859 ^ b1859 ^ c1859;
  assign sub1859 = a1859 ^ b_inv1859 ^ c1859;
  assign and1859 = a1859 & b1859;
  assign or1859  = a1859 | b1859;
  assign c1860 = (a1859 & b1859) | (a1859 & c1859) | (b1859 & c1859);
  wire c_sub1860;
  assign c_sub1860 = (a1859 & b_inv1859) | (a1859 & c1859) | (b_inv1859 & c1859);
  wire s1860, sub1860, and1860, or1860;
  wire b_inv1860;
  assign b_inv1860 = ~b1860;
  assign s1860  = a1860 ^ b1860 ^ c1860;
  assign sub1860 = a1860 ^ b_inv1860 ^ c1860;
  assign and1860 = a1860 & b1860;
  assign or1860  = a1860 | b1860;
  assign c1861 = (a1860 & b1860) | (a1860 & c1860) | (b1860 & c1860);
  wire c_sub1861;
  assign c_sub1861 = (a1860 & b_inv1860) | (a1860 & c1860) | (b_inv1860 & c1860);
  wire s1861, sub1861, and1861, or1861;
  wire b_inv1861;
  assign b_inv1861 = ~b1861;
  assign s1861  = a1861 ^ b1861 ^ c1861;
  assign sub1861 = a1861 ^ b_inv1861 ^ c1861;
  assign and1861 = a1861 & b1861;
  assign or1861  = a1861 | b1861;
  assign c1862 = (a1861 & b1861) | (a1861 & c1861) | (b1861 & c1861);
  wire c_sub1862;
  assign c_sub1862 = (a1861 & b_inv1861) | (a1861 & c1861) | (b_inv1861 & c1861);
  wire s1862, sub1862, and1862, or1862;
  wire b_inv1862;
  assign b_inv1862 = ~b1862;
  assign s1862  = a1862 ^ b1862 ^ c1862;
  assign sub1862 = a1862 ^ b_inv1862 ^ c1862;
  assign and1862 = a1862 & b1862;
  assign or1862  = a1862 | b1862;
  assign c1863 = (a1862 & b1862) | (a1862 & c1862) | (b1862 & c1862);
  wire c_sub1863;
  assign c_sub1863 = (a1862 & b_inv1862) | (a1862 & c1862) | (b_inv1862 & c1862);
  wire s1863, sub1863, and1863, or1863;
  wire b_inv1863;
  assign b_inv1863 = ~b1863;
  assign s1863  = a1863 ^ b1863 ^ c1863;
  assign sub1863 = a1863 ^ b_inv1863 ^ c1863;
  assign and1863 = a1863 & b1863;
  assign or1863  = a1863 | b1863;
  assign c1864 = (a1863 & b1863) | (a1863 & c1863) | (b1863 & c1863);
  wire c_sub1864;
  assign c_sub1864 = (a1863 & b_inv1863) | (a1863 & c1863) | (b_inv1863 & c1863);
  wire s1864, sub1864, and1864, or1864;
  wire b_inv1864;
  assign b_inv1864 = ~b1864;
  assign s1864  = a1864 ^ b1864 ^ c1864;
  assign sub1864 = a1864 ^ b_inv1864 ^ c1864;
  assign and1864 = a1864 & b1864;
  assign or1864  = a1864 | b1864;
  assign c1865 = (a1864 & b1864) | (a1864 & c1864) | (b1864 & c1864);
  wire c_sub1865;
  assign c_sub1865 = (a1864 & b_inv1864) | (a1864 & c1864) | (b_inv1864 & c1864);
  wire s1865, sub1865, and1865, or1865;
  wire b_inv1865;
  assign b_inv1865 = ~b1865;
  assign s1865  = a1865 ^ b1865 ^ c1865;
  assign sub1865 = a1865 ^ b_inv1865 ^ c1865;
  assign and1865 = a1865 & b1865;
  assign or1865  = a1865 | b1865;
  assign c1866 = (a1865 & b1865) | (a1865 & c1865) | (b1865 & c1865);
  wire c_sub1866;
  assign c_sub1866 = (a1865 & b_inv1865) | (a1865 & c1865) | (b_inv1865 & c1865);
  wire s1866, sub1866, and1866, or1866;
  wire b_inv1866;
  assign b_inv1866 = ~b1866;
  assign s1866  = a1866 ^ b1866 ^ c1866;
  assign sub1866 = a1866 ^ b_inv1866 ^ c1866;
  assign and1866 = a1866 & b1866;
  assign or1866  = a1866 | b1866;
  assign c1867 = (a1866 & b1866) | (a1866 & c1866) | (b1866 & c1866);
  wire c_sub1867;
  assign c_sub1867 = (a1866 & b_inv1866) | (a1866 & c1866) | (b_inv1866 & c1866);
  wire s1867, sub1867, and1867, or1867;
  wire b_inv1867;
  assign b_inv1867 = ~b1867;
  assign s1867  = a1867 ^ b1867 ^ c1867;
  assign sub1867 = a1867 ^ b_inv1867 ^ c1867;
  assign and1867 = a1867 & b1867;
  assign or1867  = a1867 | b1867;
  assign c1868 = (a1867 & b1867) | (a1867 & c1867) | (b1867 & c1867);
  wire c_sub1868;
  assign c_sub1868 = (a1867 & b_inv1867) | (a1867 & c1867) | (b_inv1867 & c1867);
  wire s1868, sub1868, and1868, or1868;
  wire b_inv1868;
  assign b_inv1868 = ~b1868;
  assign s1868  = a1868 ^ b1868 ^ c1868;
  assign sub1868 = a1868 ^ b_inv1868 ^ c1868;
  assign and1868 = a1868 & b1868;
  assign or1868  = a1868 | b1868;
  assign c1869 = (a1868 & b1868) | (a1868 & c1868) | (b1868 & c1868);
  wire c_sub1869;
  assign c_sub1869 = (a1868 & b_inv1868) | (a1868 & c1868) | (b_inv1868 & c1868);
  wire s1869, sub1869, and1869, or1869;
  wire b_inv1869;
  assign b_inv1869 = ~b1869;
  assign s1869  = a1869 ^ b1869 ^ c1869;
  assign sub1869 = a1869 ^ b_inv1869 ^ c1869;
  assign and1869 = a1869 & b1869;
  assign or1869  = a1869 | b1869;
  assign c1870 = (a1869 & b1869) | (a1869 & c1869) | (b1869 & c1869);
  wire c_sub1870;
  assign c_sub1870 = (a1869 & b_inv1869) | (a1869 & c1869) | (b_inv1869 & c1869);
  wire s1870, sub1870, and1870, or1870;
  wire b_inv1870;
  assign b_inv1870 = ~b1870;
  assign s1870  = a1870 ^ b1870 ^ c1870;
  assign sub1870 = a1870 ^ b_inv1870 ^ c1870;
  assign and1870 = a1870 & b1870;
  assign or1870  = a1870 | b1870;
  assign c1871 = (a1870 & b1870) | (a1870 & c1870) | (b1870 & c1870);
  wire c_sub1871;
  assign c_sub1871 = (a1870 & b_inv1870) | (a1870 & c1870) | (b_inv1870 & c1870);
  wire s1871, sub1871, and1871, or1871;
  wire b_inv1871;
  assign b_inv1871 = ~b1871;
  assign s1871  = a1871 ^ b1871 ^ c1871;
  assign sub1871 = a1871 ^ b_inv1871 ^ c1871;
  assign and1871 = a1871 & b1871;
  assign or1871  = a1871 | b1871;
  assign c1872 = (a1871 & b1871) | (a1871 & c1871) | (b1871 & c1871);
  wire c_sub1872;
  assign c_sub1872 = (a1871 & b_inv1871) | (a1871 & c1871) | (b_inv1871 & c1871);
  wire s1872, sub1872, and1872, or1872;
  wire b_inv1872;
  assign b_inv1872 = ~b1872;
  assign s1872  = a1872 ^ b1872 ^ c1872;
  assign sub1872 = a1872 ^ b_inv1872 ^ c1872;
  assign and1872 = a1872 & b1872;
  assign or1872  = a1872 | b1872;
  assign c1873 = (a1872 & b1872) | (a1872 & c1872) | (b1872 & c1872);
  wire c_sub1873;
  assign c_sub1873 = (a1872 & b_inv1872) | (a1872 & c1872) | (b_inv1872 & c1872);
  wire s1873, sub1873, and1873, or1873;
  wire b_inv1873;
  assign b_inv1873 = ~b1873;
  assign s1873  = a1873 ^ b1873 ^ c1873;
  assign sub1873 = a1873 ^ b_inv1873 ^ c1873;
  assign and1873 = a1873 & b1873;
  assign or1873  = a1873 | b1873;
  assign c1874 = (a1873 & b1873) | (a1873 & c1873) | (b1873 & c1873);
  wire c_sub1874;
  assign c_sub1874 = (a1873 & b_inv1873) | (a1873 & c1873) | (b_inv1873 & c1873);
  wire s1874, sub1874, and1874, or1874;
  wire b_inv1874;
  assign b_inv1874 = ~b1874;
  assign s1874  = a1874 ^ b1874 ^ c1874;
  assign sub1874 = a1874 ^ b_inv1874 ^ c1874;
  assign and1874 = a1874 & b1874;
  assign or1874  = a1874 | b1874;
  assign c1875 = (a1874 & b1874) | (a1874 & c1874) | (b1874 & c1874);
  wire c_sub1875;
  assign c_sub1875 = (a1874 & b_inv1874) | (a1874 & c1874) | (b_inv1874 & c1874);
  wire s1875, sub1875, and1875, or1875;
  wire b_inv1875;
  assign b_inv1875 = ~b1875;
  assign s1875  = a1875 ^ b1875 ^ c1875;
  assign sub1875 = a1875 ^ b_inv1875 ^ c1875;
  assign and1875 = a1875 & b1875;
  assign or1875  = a1875 | b1875;
  assign c1876 = (a1875 & b1875) | (a1875 & c1875) | (b1875 & c1875);
  wire c_sub1876;
  assign c_sub1876 = (a1875 & b_inv1875) | (a1875 & c1875) | (b_inv1875 & c1875);
  wire s1876, sub1876, and1876, or1876;
  wire b_inv1876;
  assign b_inv1876 = ~b1876;
  assign s1876  = a1876 ^ b1876 ^ c1876;
  assign sub1876 = a1876 ^ b_inv1876 ^ c1876;
  assign and1876 = a1876 & b1876;
  assign or1876  = a1876 | b1876;
  assign c1877 = (a1876 & b1876) | (a1876 & c1876) | (b1876 & c1876);
  wire c_sub1877;
  assign c_sub1877 = (a1876 & b_inv1876) | (a1876 & c1876) | (b_inv1876 & c1876);
  wire s1877, sub1877, and1877, or1877;
  wire b_inv1877;
  assign b_inv1877 = ~b1877;
  assign s1877  = a1877 ^ b1877 ^ c1877;
  assign sub1877 = a1877 ^ b_inv1877 ^ c1877;
  assign and1877 = a1877 & b1877;
  assign or1877  = a1877 | b1877;
  assign c1878 = (a1877 & b1877) | (a1877 & c1877) | (b1877 & c1877);
  wire c_sub1878;
  assign c_sub1878 = (a1877 & b_inv1877) | (a1877 & c1877) | (b_inv1877 & c1877);
  wire s1878, sub1878, and1878, or1878;
  wire b_inv1878;
  assign b_inv1878 = ~b1878;
  assign s1878  = a1878 ^ b1878 ^ c1878;
  assign sub1878 = a1878 ^ b_inv1878 ^ c1878;
  assign and1878 = a1878 & b1878;
  assign or1878  = a1878 | b1878;
  assign c1879 = (a1878 & b1878) | (a1878 & c1878) | (b1878 & c1878);
  wire c_sub1879;
  assign c_sub1879 = (a1878 & b_inv1878) | (a1878 & c1878) | (b_inv1878 & c1878);
  wire s1879, sub1879, and1879, or1879;
  wire b_inv1879;
  assign b_inv1879 = ~b1879;
  assign s1879  = a1879 ^ b1879 ^ c1879;
  assign sub1879 = a1879 ^ b_inv1879 ^ c1879;
  assign and1879 = a1879 & b1879;
  assign or1879  = a1879 | b1879;
  assign c1880 = (a1879 & b1879) | (a1879 & c1879) | (b1879 & c1879);
  wire c_sub1880;
  assign c_sub1880 = (a1879 & b_inv1879) | (a1879 & c1879) | (b_inv1879 & c1879);
  wire s1880, sub1880, and1880, or1880;
  wire b_inv1880;
  assign b_inv1880 = ~b1880;
  assign s1880  = a1880 ^ b1880 ^ c1880;
  assign sub1880 = a1880 ^ b_inv1880 ^ c1880;
  assign and1880 = a1880 & b1880;
  assign or1880  = a1880 | b1880;
  assign c1881 = (a1880 & b1880) | (a1880 & c1880) | (b1880 & c1880);
  wire c_sub1881;
  assign c_sub1881 = (a1880 & b_inv1880) | (a1880 & c1880) | (b_inv1880 & c1880);
  wire s1881, sub1881, and1881, or1881;
  wire b_inv1881;
  assign b_inv1881 = ~b1881;
  assign s1881  = a1881 ^ b1881 ^ c1881;
  assign sub1881 = a1881 ^ b_inv1881 ^ c1881;
  assign and1881 = a1881 & b1881;
  assign or1881  = a1881 | b1881;
  assign c1882 = (a1881 & b1881) | (a1881 & c1881) | (b1881 & c1881);
  wire c_sub1882;
  assign c_sub1882 = (a1881 & b_inv1881) | (a1881 & c1881) | (b_inv1881 & c1881);
  wire s1882, sub1882, and1882, or1882;
  wire b_inv1882;
  assign b_inv1882 = ~b1882;
  assign s1882  = a1882 ^ b1882 ^ c1882;
  assign sub1882 = a1882 ^ b_inv1882 ^ c1882;
  assign and1882 = a1882 & b1882;
  assign or1882  = a1882 | b1882;
  assign c1883 = (a1882 & b1882) | (a1882 & c1882) | (b1882 & c1882);
  wire c_sub1883;
  assign c_sub1883 = (a1882 & b_inv1882) | (a1882 & c1882) | (b_inv1882 & c1882);
  wire s1883, sub1883, and1883, or1883;
  wire b_inv1883;
  assign b_inv1883 = ~b1883;
  assign s1883  = a1883 ^ b1883 ^ c1883;
  assign sub1883 = a1883 ^ b_inv1883 ^ c1883;
  assign and1883 = a1883 & b1883;
  assign or1883  = a1883 | b1883;
  assign c1884 = (a1883 & b1883) | (a1883 & c1883) | (b1883 & c1883);
  wire c_sub1884;
  assign c_sub1884 = (a1883 & b_inv1883) | (a1883 & c1883) | (b_inv1883 & c1883);
  wire s1884, sub1884, and1884, or1884;
  wire b_inv1884;
  assign b_inv1884 = ~b1884;
  assign s1884  = a1884 ^ b1884 ^ c1884;
  assign sub1884 = a1884 ^ b_inv1884 ^ c1884;
  assign and1884 = a1884 & b1884;
  assign or1884  = a1884 | b1884;
  assign c1885 = (a1884 & b1884) | (a1884 & c1884) | (b1884 & c1884);
  wire c_sub1885;
  assign c_sub1885 = (a1884 & b_inv1884) | (a1884 & c1884) | (b_inv1884 & c1884);
  wire s1885, sub1885, and1885, or1885;
  wire b_inv1885;
  assign b_inv1885 = ~b1885;
  assign s1885  = a1885 ^ b1885 ^ c1885;
  assign sub1885 = a1885 ^ b_inv1885 ^ c1885;
  assign and1885 = a1885 & b1885;
  assign or1885  = a1885 | b1885;
  assign c1886 = (a1885 & b1885) | (a1885 & c1885) | (b1885 & c1885);
  wire c_sub1886;
  assign c_sub1886 = (a1885 & b_inv1885) | (a1885 & c1885) | (b_inv1885 & c1885);
  wire s1886, sub1886, and1886, or1886;
  wire b_inv1886;
  assign b_inv1886 = ~b1886;
  assign s1886  = a1886 ^ b1886 ^ c1886;
  assign sub1886 = a1886 ^ b_inv1886 ^ c1886;
  assign and1886 = a1886 & b1886;
  assign or1886  = a1886 | b1886;
  assign c1887 = (a1886 & b1886) | (a1886 & c1886) | (b1886 & c1886);
  wire c_sub1887;
  assign c_sub1887 = (a1886 & b_inv1886) | (a1886 & c1886) | (b_inv1886 & c1886);
  wire s1887, sub1887, and1887, or1887;
  wire b_inv1887;
  assign b_inv1887 = ~b1887;
  assign s1887  = a1887 ^ b1887 ^ c1887;
  assign sub1887 = a1887 ^ b_inv1887 ^ c1887;
  assign and1887 = a1887 & b1887;
  assign or1887  = a1887 | b1887;
  assign c1888 = (a1887 & b1887) | (a1887 & c1887) | (b1887 & c1887);
  wire c_sub1888;
  assign c_sub1888 = (a1887 & b_inv1887) | (a1887 & c1887) | (b_inv1887 & c1887);
  wire s1888, sub1888, and1888, or1888;
  wire b_inv1888;
  assign b_inv1888 = ~b1888;
  assign s1888  = a1888 ^ b1888 ^ c1888;
  assign sub1888 = a1888 ^ b_inv1888 ^ c1888;
  assign and1888 = a1888 & b1888;
  assign or1888  = a1888 | b1888;
  assign c1889 = (a1888 & b1888) | (a1888 & c1888) | (b1888 & c1888);
  wire c_sub1889;
  assign c_sub1889 = (a1888 & b_inv1888) | (a1888 & c1888) | (b_inv1888 & c1888);
  wire s1889, sub1889, and1889, or1889;
  wire b_inv1889;
  assign b_inv1889 = ~b1889;
  assign s1889  = a1889 ^ b1889 ^ c1889;
  assign sub1889 = a1889 ^ b_inv1889 ^ c1889;
  assign and1889 = a1889 & b1889;
  assign or1889  = a1889 | b1889;
  assign c1890 = (a1889 & b1889) | (a1889 & c1889) | (b1889 & c1889);
  wire c_sub1890;
  assign c_sub1890 = (a1889 & b_inv1889) | (a1889 & c1889) | (b_inv1889 & c1889);
  wire s1890, sub1890, and1890, or1890;
  wire b_inv1890;
  assign b_inv1890 = ~b1890;
  assign s1890  = a1890 ^ b1890 ^ c1890;
  assign sub1890 = a1890 ^ b_inv1890 ^ c1890;
  assign and1890 = a1890 & b1890;
  assign or1890  = a1890 | b1890;
  assign c1891 = (a1890 & b1890) | (a1890 & c1890) | (b1890 & c1890);
  wire c_sub1891;
  assign c_sub1891 = (a1890 & b_inv1890) | (a1890 & c1890) | (b_inv1890 & c1890);
  wire s1891, sub1891, and1891, or1891;
  wire b_inv1891;
  assign b_inv1891 = ~b1891;
  assign s1891  = a1891 ^ b1891 ^ c1891;
  assign sub1891 = a1891 ^ b_inv1891 ^ c1891;
  assign and1891 = a1891 & b1891;
  assign or1891  = a1891 | b1891;
  assign c1892 = (a1891 & b1891) | (a1891 & c1891) | (b1891 & c1891);
  wire c_sub1892;
  assign c_sub1892 = (a1891 & b_inv1891) | (a1891 & c1891) | (b_inv1891 & c1891);
  wire s1892, sub1892, and1892, or1892;
  wire b_inv1892;
  assign b_inv1892 = ~b1892;
  assign s1892  = a1892 ^ b1892 ^ c1892;
  assign sub1892 = a1892 ^ b_inv1892 ^ c1892;
  assign and1892 = a1892 & b1892;
  assign or1892  = a1892 | b1892;
  assign c1893 = (a1892 & b1892) | (a1892 & c1892) | (b1892 & c1892);
  wire c_sub1893;
  assign c_sub1893 = (a1892 & b_inv1892) | (a1892 & c1892) | (b_inv1892 & c1892);
  wire s1893, sub1893, and1893, or1893;
  wire b_inv1893;
  assign b_inv1893 = ~b1893;
  assign s1893  = a1893 ^ b1893 ^ c1893;
  assign sub1893 = a1893 ^ b_inv1893 ^ c1893;
  assign and1893 = a1893 & b1893;
  assign or1893  = a1893 | b1893;
  assign c1894 = (a1893 & b1893) | (a1893 & c1893) | (b1893 & c1893);
  wire c_sub1894;
  assign c_sub1894 = (a1893 & b_inv1893) | (a1893 & c1893) | (b_inv1893 & c1893);
  wire s1894, sub1894, and1894, or1894;
  wire b_inv1894;
  assign b_inv1894 = ~b1894;
  assign s1894  = a1894 ^ b1894 ^ c1894;
  assign sub1894 = a1894 ^ b_inv1894 ^ c1894;
  assign and1894 = a1894 & b1894;
  assign or1894  = a1894 | b1894;
  assign c1895 = (a1894 & b1894) | (a1894 & c1894) | (b1894 & c1894);
  wire c_sub1895;
  assign c_sub1895 = (a1894 & b_inv1894) | (a1894 & c1894) | (b_inv1894 & c1894);
  wire s1895, sub1895, and1895, or1895;
  wire b_inv1895;
  assign b_inv1895 = ~b1895;
  assign s1895  = a1895 ^ b1895 ^ c1895;
  assign sub1895 = a1895 ^ b_inv1895 ^ c1895;
  assign and1895 = a1895 & b1895;
  assign or1895  = a1895 | b1895;
  assign c1896 = (a1895 & b1895) | (a1895 & c1895) | (b1895 & c1895);
  wire c_sub1896;
  assign c_sub1896 = (a1895 & b_inv1895) | (a1895 & c1895) | (b_inv1895 & c1895);
  wire s1896, sub1896, and1896, or1896;
  wire b_inv1896;
  assign b_inv1896 = ~b1896;
  assign s1896  = a1896 ^ b1896 ^ c1896;
  assign sub1896 = a1896 ^ b_inv1896 ^ c1896;
  assign and1896 = a1896 & b1896;
  assign or1896  = a1896 | b1896;
  assign c1897 = (a1896 & b1896) | (a1896 & c1896) | (b1896 & c1896);
  wire c_sub1897;
  assign c_sub1897 = (a1896 & b_inv1896) | (a1896 & c1896) | (b_inv1896 & c1896);
  wire s1897, sub1897, and1897, or1897;
  wire b_inv1897;
  assign b_inv1897 = ~b1897;
  assign s1897  = a1897 ^ b1897 ^ c1897;
  assign sub1897 = a1897 ^ b_inv1897 ^ c1897;
  assign and1897 = a1897 & b1897;
  assign or1897  = a1897 | b1897;
  assign c1898 = (a1897 & b1897) | (a1897 & c1897) | (b1897 & c1897);
  wire c_sub1898;
  assign c_sub1898 = (a1897 & b_inv1897) | (a1897 & c1897) | (b_inv1897 & c1897);
  wire s1898, sub1898, and1898, or1898;
  wire b_inv1898;
  assign b_inv1898 = ~b1898;
  assign s1898  = a1898 ^ b1898 ^ c1898;
  assign sub1898 = a1898 ^ b_inv1898 ^ c1898;
  assign and1898 = a1898 & b1898;
  assign or1898  = a1898 | b1898;
  assign c1899 = (a1898 & b1898) | (a1898 & c1898) | (b1898 & c1898);
  wire c_sub1899;
  assign c_sub1899 = (a1898 & b_inv1898) | (a1898 & c1898) | (b_inv1898 & c1898);
  wire s1899, sub1899, and1899, or1899;
  wire b_inv1899;
  assign b_inv1899 = ~b1899;
  assign s1899  = a1899 ^ b1899 ^ c1899;
  assign sub1899 = a1899 ^ b_inv1899 ^ c1899;
  assign and1899 = a1899 & b1899;
  assign or1899  = a1899 | b1899;
  assign c1900 = (a1899 & b1899) | (a1899 & c1899) | (b1899 & c1899);
  wire c_sub1900;
  assign c_sub1900 = (a1899 & b_inv1899) | (a1899 & c1899) | (b_inv1899 & c1899);
  wire s1900, sub1900, and1900, or1900;
  wire b_inv1900;
  assign b_inv1900 = ~b1900;
  assign s1900  = a1900 ^ b1900 ^ c1900;
  assign sub1900 = a1900 ^ b_inv1900 ^ c1900;
  assign and1900 = a1900 & b1900;
  assign or1900  = a1900 | b1900;
  assign c1901 = (a1900 & b1900) | (a1900 & c1900) | (b1900 & c1900);
  wire c_sub1901;
  assign c_sub1901 = (a1900 & b_inv1900) | (a1900 & c1900) | (b_inv1900 & c1900);
  wire s1901, sub1901, and1901, or1901;
  wire b_inv1901;
  assign b_inv1901 = ~b1901;
  assign s1901  = a1901 ^ b1901 ^ c1901;
  assign sub1901 = a1901 ^ b_inv1901 ^ c1901;
  assign and1901 = a1901 & b1901;
  assign or1901  = a1901 | b1901;
  assign c1902 = (a1901 & b1901) | (a1901 & c1901) | (b1901 & c1901);
  wire c_sub1902;
  assign c_sub1902 = (a1901 & b_inv1901) | (a1901 & c1901) | (b_inv1901 & c1901);
  wire s1902, sub1902, and1902, or1902;
  wire b_inv1902;
  assign b_inv1902 = ~b1902;
  assign s1902  = a1902 ^ b1902 ^ c1902;
  assign sub1902 = a1902 ^ b_inv1902 ^ c1902;
  assign and1902 = a1902 & b1902;
  assign or1902  = a1902 | b1902;
  assign c1903 = (a1902 & b1902) | (a1902 & c1902) | (b1902 & c1902);
  wire c_sub1903;
  assign c_sub1903 = (a1902 & b_inv1902) | (a1902 & c1902) | (b_inv1902 & c1902);
  wire s1903, sub1903, and1903, or1903;
  wire b_inv1903;
  assign b_inv1903 = ~b1903;
  assign s1903  = a1903 ^ b1903 ^ c1903;
  assign sub1903 = a1903 ^ b_inv1903 ^ c1903;
  assign and1903 = a1903 & b1903;
  assign or1903  = a1903 | b1903;
  assign c1904 = (a1903 & b1903) | (a1903 & c1903) | (b1903 & c1903);
  wire c_sub1904;
  assign c_sub1904 = (a1903 & b_inv1903) | (a1903 & c1903) | (b_inv1903 & c1903);
  wire s1904, sub1904, and1904, or1904;
  wire b_inv1904;
  assign b_inv1904 = ~b1904;
  assign s1904  = a1904 ^ b1904 ^ c1904;
  assign sub1904 = a1904 ^ b_inv1904 ^ c1904;
  assign and1904 = a1904 & b1904;
  assign or1904  = a1904 | b1904;
  assign c1905 = (a1904 & b1904) | (a1904 & c1904) | (b1904 & c1904);
  wire c_sub1905;
  assign c_sub1905 = (a1904 & b_inv1904) | (a1904 & c1904) | (b_inv1904 & c1904);
  wire s1905, sub1905, and1905, or1905;
  wire b_inv1905;
  assign b_inv1905 = ~b1905;
  assign s1905  = a1905 ^ b1905 ^ c1905;
  assign sub1905 = a1905 ^ b_inv1905 ^ c1905;
  assign and1905 = a1905 & b1905;
  assign or1905  = a1905 | b1905;
  assign c1906 = (a1905 & b1905) | (a1905 & c1905) | (b1905 & c1905);
  wire c_sub1906;
  assign c_sub1906 = (a1905 & b_inv1905) | (a1905 & c1905) | (b_inv1905 & c1905);
  wire s1906, sub1906, and1906, or1906;
  wire b_inv1906;
  assign b_inv1906 = ~b1906;
  assign s1906  = a1906 ^ b1906 ^ c1906;
  assign sub1906 = a1906 ^ b_inv1906 ^ c1906;
  assign and1906 = a1906 & b1906;
  assign or1906  = a1906 | b1906;
  assign c1907 = (a1906 & b1906) | (a1906 & c1906) | (b1906 & c1906);
  wire c_sub1907;
  assign c_sub1907 = (a1906 & b_inv1906) | (a1906 & c1906) | (b_inv1906 & c1906);
  wire s1907, sub1907, and1907, or1907;
  wire b_inv1907;
  assign b_inv1907 = ~b1907;
  assign s1907  = a1907 ^ b1907 ^ c1907;
  assign sub1907 = a1907 ^ b_inv1907 ^ c1907;
  assign and1907 = a1907 & b1907;
  assign or1907  = a1907 | b1907;
  assign c1908 = (a1907 & b1907) | (a1907 & c1907) | (b1907 & c1907);
  wire c_sub1908;
  assign c_sub1908 = (a1907 & b_inv1907) | (a1907 & c1907) | (b_inv1907 & c1907);
  wire s1908, sub1908, and1908, or1908;
  wire b_inv1908;
  assign b_inv1908 = ~b1908;
  assign s1908  = a1908 ^ b1908 ^ c1908;
  assign sub1908 = a1908 ^ b_inv1908 ^ c1908;
  assign and1908 = a1908 & b1908;
  assign or1908  = a1908 | b1908;
  assign c1909 = (a1908 & b1908) | (a1908 & c1908) | (b1908 & c1908);
  wire c_sub1909;
  assign c_sub1909 = (a1908 & b_inv1908) | (a1908 & c1908) | (b_inv1908 & c1908);
  wire s1909, sub1909, and1909, or1909;
  wire b_inv1909;
  assign b_inv1909 = ~b1909;
  assign s1909  = a1909 ^ b1909 ^ c1909;
  assign sub1909 = a1909 ^ b_inv1909 ^ c1909;
  assign and1909 = a1909 & b1909;
  assign or1909  = a1909 | b1909;
  assign c1910 = (a1909 & b1909) | (a1909 & c1909) | (b1909 & c1909);
  wire c_sub1910;
  assign c_sub1910 = (a1909 & b_inv1909) | (a1909 & c1909) | (b_inv1909 & c1909);
  wire s1910, sub1910, and1910, or1910;
  wire b_inv1910;
  assign b_inv1910 = ~b1910;
  assign s1910  = a1910 ^ b1910 ^ c1910;
  assign sub1910 = a1910 ^ b_inv1910 ^ c1910;
  assign and1910 = a1910 & b1910;
  assign or1910  = a1910 | b1910;
  assign c1911 = (a1910 & b1910) | (a1910 & c1910) | (b1910 & c1910);
  wire c_sub1911;
  assign c_sub1911 = (a1910 & b_inv1910) | (a1910 & c1910) | (b_inv1910 & c1910);
  wire s1911, sub1911, and1911, or1911;
  wire b_inv1911;
  assign b_inv1911 = ~b1911;
  assign s1911  = a1911 ^ b1911 ^ c1911;
  assign sub1911 = a1911 ^ b_inv1911 ^ c1911;
  assign and1911 = a1911 & b1911;
  assign or1911  = a1911 | b1911;
  assign c1912 = (a1911 & b1911) | (a1911 & c1911) | (b1911 & c1911);
  wire c_sub1912;
  assign c_sub1912 = (a1911 & b_inv1911) | (a1911 & c1911) | (b_inv1911 & c1911);
  wire s1912, sub1912, and1912, or1912;
  wire b_inv1912;
  assign b_inv1912 = ~b1912;
  assign s1912  = a1912 ^ b1912 ^ c1912;
  assign sub1912 = a1912 ^ b_inv1912 ^ c1912;
  assign and1912 = a1912 & b1912;
  assign or1912  = a1912 | b1912;
  assign c1913 = (a1912 & b1912) | (a1912 & c1912) | (b1912 & c1912);
  wire c_sub1913;
  assign c_sub1913 = (a1912 & b_inv1912) | (a1912 & c1912) | (b_inv1912 & c1912);
  wire s1913, sub1913, and1913, or1913;
  wire b_inv1913;
  assign b_inv1913 = ~b1913;
  assign s1913  = a1913 ^ b1913 ^ c1913;
  assign sub1913 = a1913 ^ b_inv1913 ^ c1913;
  assign and1913 = a1913 & b1913;
  assign or1913  = a1913 | b1913;
  assign c1914 = (a1913 & b1913) | (a1913 & c1913) | (b1913 & c1913);
  wire c_sub1914;
  assign c_sub1914 = (a1913 & b_inv1913) | (a1913 & c1913) | (b_inv1913 & c1913);
  wire s1914, sub1914, and1914, or1914;
  wire b_inv1914;
  assign b_inv1914 = ~b1914;
  assign s1914  = a1914 ^ b1914 ^ c1914;
  assign sub1914 = a1914 ^ b_inv1914 ^ c1914;
  assign and1914 = a1914 & b1914;
  assign or1914  = a1914 | b1914;
  assign c1915 = (a1914 & b1914) | (a1914 & c1914) | (b1914 & c1914);
  wire c_sub1915;
  assign c_sub1915 = (a1914 & b_inv1914) | (a1914 & c1914) | (b_inv1914 & c1914);
  wire s1915, sub1915, and1915, or1915;
  wire b_inv1915;
  assign b_inv1915 = ~b1915;
  assign s1915  = a1915 ^ b1915 ^ c1915;
  assign sub1915 = a1915 ^ b_inv1915 ^ c1915;
  assign and1915 = a1915 & b1915;
  assign or1915  = a1915 | b1915;
  assign c1916 = (a1915 & b1915) | (a1915 & c1915) | (b1915 & c1915);
  wire c_sub1916;
  assign c_sub1916 = (a1915 & b_inv1915) | (a1915 & c1915) | (b_inv1915 & c1915);
  wire s1916, sub1916, and1916, or1916;
  wire b_inv1916;
  assign b_inv1916 = ~b1916;
  assign s1916  = a1916 ^ b1916 ^ c1916;
  assign sub1916 = a1916 ^ b_inv1916 ^ c1916;
  assign and1916 = a1916 & b1916;
  assign or1916  = a1916 | b1916;
  assign c1917 = (a1916 & b1916) | (a1916 & c1916) | (b1916 & c1916);
  wire c_sub1917;
  assign c_sub1917 = (a1916 & b_inv1916) | (a1916 & c1916) | (b_inv1916 & c1916);
  wire s1917, sub1917, and1917, or1917;
  wire b_inv1917;
  assign b_inv1917 = ~b1917;
  assign s1917  = a1917 ^ b1917 ^ c1917;
  assign sub1917 = a1917 ^ b_inv1917 ^ c1917;
  assign and1917 = a1917 & b1917;
  assign or1917  = a1917 | b1917;
  assign c1918 = (a1917 & b1917) | (a1917 & c1917) | (b1917 & c1917);
  wire c_sub1918;
  assign c_sub1918 = (a1917 & b_inv1917) | (a1917 & c1917) | (b_inv1917 & c1917);
  wire s1918, sub1918, and1918, or1918;
  wire b_inv1918;
  assign b_inv1918 = ~b1918;
  assign s1918  = a1918 ^ b1918 ^ c1918;
  assign sub1918 = a1918 ^ b_inv1918 ^ c1918;
  assign and1918 = a1918 & b1918;
  assign or1918  = a1918 | b1918;
  assign c1919 = (a1918 & b1918) | (a1918 & c1918) | (b1918 & c1918);
  wire c_sub1919;
  assign c_sub1919 = (a1918 & b_inv1918) | (a1918 & c1918) | (b_inv1918 & c1918);
  wire s1919, sub1919, and1919, or1919;
  wire b_inv1919;
  assign b_inv1919 = ~b1919;
  assign s1919  = a1919 ^ b1919 ^ c1919;
  assign sub1919 = a1919 ^ b_inv1919 ^ c1919;
  assign and1919 = a1919 & b1919;
  assign or1919  = a1919 | b1919;
  assign c1920 = (a1919 & b1919) | (a1919 & c1919) | (b1919 & c1919);
  wire c_sub1920;
  assign c_sub1920 = (a1919 & b_inv1919) | (a1919 & c1919) | (b_inv1919 & c1919);
  wire s1920, sub1920, and1920, or1920;
  wire b_inv1920;
  assign b_inv1920 = ~b1920;
  assign s1920  = a1920 ^ b1920 ^ c1920;
  assign sub1920 = a1920 ^ b_inv1920 ^ c1920;
  assign and1920 = a1920 & b1920;
  assign or1920  = a1920 | b1920;
  assign c1921 = (a1920 & b1920) | (a1920 & c1920) | (b1920 & c1920);
  wire c_sub1921;
  assign c_sub1921 = (a1920 & b_inv1920) | (a1920 & c1920) | (b_inv1920 & c1920);
  wire s1921, sub1921, and1921, or1921;
  wire b_inv1921;
  assign b_inv1921 = ~b1921;
  assign s1921  = a1921 ^ b1921 ^ c1921;
  assign sub1921 = a1921 ^ b_inv1921 ^ c1921;
  assign and1921 = a1921 & b1921;
  assign or1921  = a1921 | b1921;
  assign c1922 = (a1921 & b1921) | (a1921 & c1921) | (b1921 & c1921);
  wire c_sub1922;
  assign c_sub1922 = (a1921 & b_inv1921) | (a1921 & c1921) | (b_inv1921 & c1921);
  wire s1922, sub1922, and1922, or1922;
  wire b_inv1922;
  assign b_inv1922 = ~b1922;
  assign s1922  = a1922 ^ b1922 ^ c1922;
  assign sub1922 = a1922 ^ b_inv1922 ^ c1922;
  assign and1922 = a1922 & b1922;
  assign or1922  = a1922 | b1922;
  assign c1923 = (a1922 & b1922) | (a1922 & c1922) | (b1922 & c1922);
  wire c_sub1923;
  assign c_sub1923 = (a1922 & b_inv1922) | (a1922 & c1922) | (b_inv1922 & c1922);
  wire s1923, sub1923, and1923, or1923;
  wire b_inv1923;
  assign b_inv1923 = ~b1923;
  assign s1923  = a1923 ^ b1923 ^ c1923;
  assign sub1923 = a1923 ^ b_inv1923 ^ c1923;
  assign and1923 = a1923 & b1923;
  assign or1923  = a1923 | b1923;
  assign c1924 = (a1923 & b1923) | (a1923 & c1923) | (b1923 & c1923);
  wire c_sub1924;
  assign c_sub1924 = (a1923 & b_inv1923) | (a1923 & c1923) | (b_inv1923 & c1923);
  wire s1924, sub1924, and1924, or1924;
  wire b_inv1924;
  assign b_inv1924 = ~b1924;
  assign s1924  = a1924 ^ b1924 ^ c1924;
  assign sub1924 = a1924 ^ b_inv1924 ^ c1924;
  assign and1924 = a1924 & b1924;
  assign or1924  = a1924 | b1924;
  assign c1925 = (a1924 & b1924) | (a1924 & c1924) | (b1924 & c1924);
  wire c_sub1925;
  assign c_sub1925 = (a1924 & b_inv1924) | (a1924 & c1924) | (b_inv1924 & c1924);
  wire s1925, sub1925, and1925, or1925;
  wire b_inv1925;
  assign b_inv1925 = ~b1925;
  assign s1925  = a1925 ^ b1925 ^ c1925;
  assign sub1925 = a1925 ^ b_inv1925 ^ c1925;
  assign and1925 = a1925 & b1925;
  assign or1925  = a1925 | b1925;
  assign c1926 = (a1925 & b1925) | (a1925 & c1925) | (b1925 & c1925);
  wire c_sub1926;
  assign c_sub1926 = (a1925 & b_inv1925) | (a1925 & c1925) | (b_inv1925 & c1925);
  wire s1926, sub1926, and1926, or1926;
  wire b_inv1926;
  assign b_inv1926 = ~b1926;
  assign s1926  = a1926 ^ b1926 ^ c1926;
  assign sub1926 = a1926 ^ b_inv1926 ^ c1926;
  assign and1926 = a1926 & b1926;
  assign or1926  = a1926 | b1926;
  assign c1927 = (a1926 & b1926) | (a1926 & c1926) | (b1926 & c1926);
  wire c_sub1927;
  assign c_sub1927 = (a1926 & b_inv1926) | (a1926 & c1926) | (b_inv1926 & c1926);
  wire s1927, sub1927, and1927, or1927;
  wire b_inv1927;
  assign b_inv1927 = ~b1927;
  assign s1927  = a1927 ^ b1927 ^ c1927;
  assign sub1927 = a1927 ^ b_inv1927 ^ c1927;
  assign and1927 = a1927 & b1927;
  assign or1927  = a1927 | b1927;
  assign c1928 = (a1927 & b1927) | (a1927 & c1927) | (b1927 & c1927);
  wire c_sub1928;
  assign c_sub1928 = (a1927 & b_inv1927) | (a1927 & c1927) | (b_inv1927 & c1927);
  wire s1928, sub1928, and1928, or1928;
  wire b_inv1928;
  assign b_inv1928 = ~b1928;
  assign s1928  = a1928 ^ b1928 ^ c1928;
  assign sub1928 = a1928 ^ b_inv1928 ^ c1928;
  assign and1928 = a1928 & b1928;
  assign or1928  = a1928 | b1928;
  assign c1929 = (a1928 & b1928) | (a1928 & c1928) | (b1928 & c1928);
  wire c_sub1929;
  assign c_sub1929 = (a1928 & b_inv1928) | (a1928 & c1928) | (b_inv1928 & c1928);
  wire s1929, sub1929, and1929, or1929;
  wire b_inv1929;
  assign b_inv1929 = ~b1929;
  assign s1929  = a1929 ^ b1929 ^ c1929;
  assign sub1929 = a1929 ^ b_inv1929 ^ c1929;
  assign and1929 = a1929 & b1929;
  assign or1929  = a1929 | b1929;
  assign c1930 = (a1929 & b1929) | (a1929 & c1929) | (b1929 & c1929);
  wire c_sub1930;
  assign c_sub1930 = (a1929 & b_inv1929) | (a1929 & c1929) | (b_inv1929 & c1929);
  wire s1930, sub1930, and1930, or1930;
  wire b_inv1930;
  assign b_inv1930 = ~b1930;
  assign s1930  = a1930 ^ b1930 ^ c1930;
  assign sub1930 = a1930 ^ b_inv1930 ^ c1930;
  assign and1930 = a1930 & b1930;
  assign or1930  = a1930 | b1930;
  assign c1931 = (a1930 & b1930) | (a1930 & c1930) | (b1930 & c1930);
  wire c_sub1931;
  assign c_sub1931 = (a1930 & b_inv1930) | (a1930 & c1930) | (b_inv1930 & c1930);
  wire s1931, sub1931, and1931, or1931;
  wire b_inv1931;
  assign b_inv1931 = ~b1931;
  assign s1931  = a1931 ^ b1931 ^ c1931;
  assign sub1931 = a1931 ^ b_inv1931 ^ c1931;
  assign and1931 = a1931 & b1931;
  assign or1931  = a1931 | b1931;
  assign c1932 = (a1931 & b1931) | (a1931 & c1931) | (b1931 & c1931);
  wire c_sub1932;
  assign c_sub1932 = (a1931 & b_inv1931) | (a1931 & c1931) | (b_inv1931 & c1931);
  wire s1932, sub1932, and1932, or1932;
  wire b_inv1932;
  assign b_inv1932 = ~b1932;
  assign s1932  = a1932 ^ b1932 ^ c1932;
  assign sub1932 = a1932 ^ b_inv1932 ^ c1932;
  assign and1932 = a1932 & b1932;
  assign or1932  = a1932 | b1932;
  assign c1933 = (a1932 & b1932) | (a1932 & c1932) | (b1932 & c1932);
  wire c_sub1933;
  assign c_sub1933 = (a1932 & b_inv1932) | (a1932 & c1932) | (b_inv1932 & c1932);
  wire s1933, sub1933, and1933, or1933;
  wire b_inv1933;
  assign b_inv1933 = ~b1933;
  assign s1933  = a1933 ^ b1933 ^ c1933;
  assign sub1933 = a1933 ^ b_inv1933 ^ c1933;
  assign and1933 = a1933 & b1933;
  assign or1933  = a1933 | b1933;
  assign c1934 = (a1933 & b1933) | (a1933 & c1933) | (b1933 & c1933);
  wire c_sub1934;
  assign c_sub1934 = (a1933 & b_inv1933) | (a1933 & c1933) | (b_inv1933 & c1933);
  wire s1934, sub1934, and1934, or1934;
  wire b_inv1934;
  assign b_inv1934 = ~b1934;
  assign s1934  = a1934 ^ b1934 ^ c1934;
  assign sub1934 = a1934 ^ b_inv1934 ^ c1934;
  assign and1934 = a1934 & b1934;
  assign or1934  = a1934 | b1934;
  assign c1935 = (a1934 & b1934) | (a1934 & c1934) | (b1934 & c1934);
  wire c_sub1935;
  assign c_sub1935 = (a1934 & b_inv1934) | (a1934 & c1934) | (b_inv1934 & c1934);
  wire s1935, sub1935, and1935, or1935;
  wire b_inv1935;
  assign b_inv1935 = ~b1935;
  assign s1935  = a1935 ^ b1935 ^ c1935;
  assign sub1935 = a1935 ^ b_inv1935 ^ c1935;
  assign and1935 = a1935 & b1935;
  assign or1935  = a1935 | b1935;
  assign c1936 = (a1935 & b1935) | (a1935 & c1935) | (b1935 & c1935);
  wire c_sub1936;
  assign c_sub1936 = (a1935 & b_inv1935) | (a1935 & c1935) | (b_inv1935 & c1935);
  wire s1936, sub1936, and1936, or1936;
  wire b_inv1936;
  assign b_inv1936 = ~b1936;
  assign s1936  = a1936 ^ b1936 ^ c1936;
  assign sub1936 = a1936 ^ b_inv1936 ^ c1936;
  assign and1936 = a1936 & b1936;
  assign or1936  = a1936 | b1936;
  assign c1937 = (a1936 & b1936) | (a1936 & c1936) | (b1936 & c1936);
  wire c_sub1937;
  assign c_sub1937 = (a1936 & b_inv1936) | (a1936 & c1936) | (b_inv1936 & c1936);
  wire s1937, sub1937, and1937, or1937;
  wire b_inv1937;
  assign b_inv1937 = ~b1937;
  assign s1937  = a1937 ^ b1937 ^ c1937;
  assign sub1937 = a1937 ^ b_inv1937 ^ c1937;
  assign and1937 = a1937 & b1937;
  assign or1937  = a1937 | b1937;
  assign c1938 = (a1937 & b1937) | (a1937 & c1937) | (b1937 & c1937);
  wire c_sub1938;
  assign c_sub1938 = (a1937 & b_inv1937) | (a1937 & c1937) | (b_inv1937 & c1937);
  wire s1938, sub1938, and1938, or1938;
  wire b_inv1938;
  assign b_inv1938 = ~b1938;
  assign s1938  = a1938 ^ b1938 ^ c1938;
  assign sub1938 = a1938 ^ b_inv1938 ^ c1938;
  assign and1938 = a1938 & b1938;
  assign or1938  = a1938 | b1938;
  assign c1939 = (a1938 & b1938) | (a1938 & c1938) | (b1938 & c1938);
  wire c_sub1939;
  assign c_sub1939 = (a1938 & b_inv1938) | (a1938 & c1938) | (b_inv1938 & c1938);
  wire s1939, sub1939, and1939, or1939;
  wire b_inv1939;
  assign b_inv1939 = ~b1939;
  assign s1939  = a1939 ^ b1939 ^ c1939;
  assign sub1939 = a1939 ^ b_inv1939 ^ c1939;
  assign and1939 = a1939 & b1939;
  assign or1939  = a1939 | b1939;
  assign c1940 = (a1939 & b1939) | (a1939 & c1939) | (b1939 & c1939);
  wire c_sub1940;
  assign c_sub1940 = (a1939 & b_inv1939) | (a1939 & c1939) | (b_inv1939 & c1939);
  wire s1940, sub1940, and1940, or1940;
  wire b_inv1940;
  assign b_inv1940 = ~b1940;
  assign s1940  = a1940 ^ b1940 ^ c1940;
  assign sub1940 = a1940 ^ b_inv1940 ^ c1940;
  assign and1940 = a1940 & b1940;
  assign or1940  = a1940 | b1940;
  assign c1941 = (a1940 & b1940) | (a1940 & c1940) | (b1940 & c1940);
  wire c_sub1941;
  assign c_sub1941 = (a1940 & b_inv1940) | (a1940 & c1940) | (b_inv1940 & c1940);
  wire s1941, sub1941, and1941, or1941;
  wire b_inv1941;
  assign b_inv1941 = ~b1941;
  assign s1941  = a1941 ^ b1941 ^ c1941;
  assign sub1941 = a1941 ^ b_inv1941 ^ c1941;
  assign and1941 = a1941 & b1941;
  assign or1941  = a1941 | b1941;
  assign c1942 = (a1941 & b1941) | (a1941 & c1941) | (b1941 & c1941);
  wire c_sub1942;
  assign c_sub1942 = (a1941 & b_inv1941) | (a1941 & c1941) | (b_inv1941 & c1941);
  wire s1942, sub1942, and1942, or1942;
  wire b_inv1942;
  assign b_inv1942 = ~b1942;
  assign s1942  = a1942 ^ b1942 ^ c1942;
  assign sub1942 = a1942 ^ b_inv1942 ^ c1942;
  assign and1942 = a1942 & b1942;
  assign or1942  = a1942 | b1942;
  assign c1943 = (a1942 & b1942) | (a1942 & c1942) | (b1942 & c1942);
  wire c_sub1943;
  assign c_sub1943 = (a1942 & b_inv1942) | (a1942 & c1942) | (b_inv1942 & c1942);
  wire s1943, sub1943, and1943, or1943;
  wire b_inv1943;
  assign b_inv1943 = ~b1943;
  assign s1943  = a1943 ^ b1943 ^ c1943;
  assign sub1943 = a1943 ^ b_inv1943 ^ c1943;
  assign and1943 = a1943 & b1943;
  assign or1943  = a1943 | b1943;
  assign c1944 = (a1943 & b1943) | (a1943 & c1943) | (b1943 & c1943);
  wire c_sub1944;
  assign c_sub1944 = (a1943 & b_inv1943) | (a1943 & c1943) | (b_inv1943 & c1943);
  wire s1944, sub1944, and1944, or1944;
  wire b_inv1944;
  assign b_inv1944 = ~b1944;
  assign s1944  = a1944 ^ b1944 ^ c1944;
  assign sub1944 = a1944 ^ b_inv1944 ^ c1944;
  assign and1944 = a1944 & b1944;
  assign or1944  = a1944 | b1944;
  assign c1945 = (a1944 & b1944) | (a1944 & c1944) | (b1944 & c1944);
  wire c_sub1945;
  assign c_sub1945 = (a1944 & b_inv1944) | (a1944 & c1944) | (b_inv1944 & c1944);
  wire s1945, sub1945, and1945, or1945;
  wire b_inv1945;
  assign b_inv1945 = ~b1945;
  assign s1945  = a1945 ^ b1945 ^ c1945;
  assign sub1945 = a1945 ^ b_inv1945 ^ c1945;
  assign and1945 = a1945 & b1945;
  assign or1945  = a1945 | b1945;
  assign c1946 = (a1945 & b1945) | (a1945 & c1945) | (b1945 & c1945);
  wire c_sub1946;
  assign c_sub1946 = (a1945 & b_inv1945) | (a1945 & c1945) | (b_inv1945 & c1945);
  wire s1946, sub1946, and1946, or1946;
  wire b_inv1946;
  assign b_inv1946 = ~b1946;
  assign s1946  = a1946 ^ b1946 ^ c1946;
  assign sub1946 = a1946 ^ b_inv1946 ^ c1946;
  assign and1946 = a1946 & b1946;
  assign or1946  = a1946 | b1946;
  assign c1947 = (a1946 & b1946) | (a1946 & c1946) | (b1946 & c1946);
  wire c_sub1947;
  assign c_sub1947 = (a1946 & b_inv1946) | (a1946 & c1946) | (b_inv1946 & c1946);
  wire s1947, sub1947, and1947, or1947;
  wire b_inv1947;
  assign b_inv1947 = ~b1947;
  assign s1947  = a1947 ^ b1947 ^ c1947;
  assign sub1947 = a1947 ^ b_inv1947 ^ c1947;
  assign and1947 = a1947 & b1947;
  assign or1947  = a1947 | b1947;
  assign c1948 = (a1947 & b1947) | (a1947 & c1947) | (b1947 & c1947);
  wire c_sub1948;
  assign c_sub1948 = (a1947 & b_inv1947) | (a1947 & c1947) | (b_inv1947 & c1947);
  wire s1948, sub1948, and1948, or1948;
  wire b_inv1948;
  assign b_inv1948 = ~b1948;
  assign s1948  = a1948 ^ b1948 ^ c1948;
  assign sub1948 = a1948 ^ b_inv1948 ^ c1948;
  assign and1948 = a1948 & b1948;
  assign or1948  = a1948 | b1948;
  assign c1949 = (a1948 & b1948) | (a1948 & c1948) | (b1948 & c1948);
  wire c_sub1949;
  assign c_sub1949 = (a1948 & b_inv1948) | (a1948 & c1948) | (b_inv1948 & c1948);
  wire s1949, sub1949, and1949, or1949;
  wire b_inv1949;
  assign b_inv1949 = ~b1949;
  assign s1949  = a1949 ^ b1949 ^ c1949;
  assign sub1949 = a1949 ^ b_inv1949 ^ c1949;
  assign and1949 = a1949 & b1949;
  assign or1949  = a1949 | b1949;
  assign c1950 = (a1949 & b1949) | (a1949 & c1949) | (b1949 & c1949);
  wire c_sub1950;
  assign c_sub1950 = (a1949 & b_inv1949) | (a1949 & c1949) | (b_inv1949 & c1949);
  wire s1950, sub1950, and1950, or1950;
  wire b_inv1950;
  assign b_inv1950 = ~b1950;
  assign s1950  = a1950 ^ b1950 ^ c1950;
  assign sub1950 = a1950 ^ b_inv1950 ^ c1950;
  assign and1950 = a1950 & b1950;
  assign or1950  = a1950 | b1950;
  assign c1951 = (a1950 & b1950) | (a1950 & c1950) | (b1950 & c1950);
  wire c_sub1951;
  assign c_sub1951 = (a1950 & b_inv1950) | (a1950 & c1950) | (b_inv1950 & c1950);
  wire s1951, sub1951, and1951, or1951;
  wire b_inv1951;
  assign b_inv1951 = ~b1951;
  assign s1951  = a1951 ^ b1951 ^ c1951;
  assign sub1951 = a1951 ^ b_inv1951 ^ c1951;
  assign and1951 = a1951 & b1951;
  assign or1951  = a1951 | b1951;
  assign c1952 = (a1951 & b1951) | (a1951 & c1951) | (b1951 & c1951);
  wire c_sub1952;
  assign c_sub1952 = (a1951 & b_inv1951) | (a1951 & c1951) | (b_inv1951 & c1951);
  wire s1952, sub1952, and1952, or1952;
  wire b_inv1952;
  assign b_inv1952 = ~b1952;
  assign s1952  = a1952 ^ b1952 ^ c1952;
  assign sub1952 = a1952 ^ b_inv1952 ^ c1952;
  assign and1952 = a1952 & b1952;
  assign or1952  = a1952 | b1952;
  assign c1953 = (a1952 & b1952) | (a1952 & c1952) | (b1952 & c1952);
  wire c_sub1953;
  assign c_sub1953 = (a1952 & b_inv1952) | (a1952 & c1952) | (b_inv1952 & c1952);
  wire s1953, sub1953, and1953, or1953;
  wire b_inv1953;
  assign b_inv1953 = ~b1953;
  assign s1953  = a1953 ^ b1953 ^ c1953;
  assign sub1953 = a1953 ^ b_inv1953 ^ c1953;
  assign and1953 = a1953 & b1953;
  assign or1953  = a1953 | b1953;
  assign c1954 = (a1953 & b1953) | (a1953 & c1953) | (b1953 & c1953);
  wire c_sub1954;
  assign c_sub1954 = (a1953 & b_inv1953) | (a1953 & c1953) | (b_inv1953 & c1953);
  wire s1954, sub1954, and1954, or1954;
  wire b_inv1954;
  assign b_inv1954 = ~b1954;
  assign s1954  = a1954 ^ b1954 ^ c1954;
  assign sub1954 = a1954 ^ b_inv1954 ^ c1954;
  assign and1954 = a1954 & b1954;
  assign or1954  = a1954 | b1954;
  assign c1955 = (a1954 & b1954) | (a1954 & c1954) | (b1954 & c1954);
  wire c_sub1955;
  assign c_sub1955 = (a1954 & b_inv1954) | (a1954 & c1954) | (b_inv1954 & c1954);
  wire s1955, sub1955, and1955, or1955;
  wire b_inv1955;
  assign b_inv1955 = ~b1955;
  assign s1955  = a1955 ^ b1955 ^ c1955;
  assign sub1955 = a1955 ^ b_inv1955 ^ c1955;
  assign and1955 = a1955 & b1955;
  assign or1955  = a1955 | b1955;
  assign c1956 = (a1955 & b1955) | (a1955 & c1955) | (b1955 & c1955);
  wire c_sub1956;
  assign c_sub1956 = (a1955 & b_inv1955) | (a1955 & c1955) | (b_inv1955 & c1955);
  wire s1956, sub1956, and1956, or1956;
  wire b_inv1956;
  assign b_inv1956 = ~b1956;
  assign s1956  = a1956 ^ b1956 ^ c1956;
  assign sub1956 = a1956 ^ b_inv1956 ^ c1956;
  assign and1956 = a1956 & b1956;
  assign or1956  = a1956 | b1956;
  assign c1957 = (a1956 & b1956) | (a1956 & c1956) | (b1956 & c1956);
  wire c_sub1957;
  assign c_sub1957 = (a1956 & b_inv1956) | (a1956 & c1956) | (b_inv1956 & c1956);
  wire s1957, sub1957, and1957, or1957;
  wire b_inv1957;
  assign b_inv1957 = ~b1957;
  assign s1957  = a1957 ^ b1957 ^ c1957;
  assign sub1957 = a1957 ^ b_inv1957 ^ c1957;
  assign and1957 = a1957 & b1957;
  assign or1957  = a1957 | b1957;
  assign c1958 = (a1957 & b1957) | (a1957 & c1957) | (b1957 & c1957);
  wire c_sub1958;
  assign c_sub1958 = (a1957 & b_inv1957) | (a1957 & c1957) | (b_inv1957 & c1957);
  wire s1958, sub1958, and1958, or1958;
  wire b_inv1958;
  assign b_inv1958 = ~b1958;
  assign s1958  = a1958 ^ b1958 ^ c1958;
  assign sub1958 = a1958 ^ b_inv1958 ^ c1958;
  assign and1958 = a1958 & b1958;
  assign or1958  = a1958 | b1958;
  assign c1959 = (a1958 & b1958) | (a1958 & c1958) | (b1958 & c1958);
  wire c_sub1959;
  assign c_sub1959 = (a1958 & b_inv1958) | (a1958 & c1958) | (b_inv1958 & c1958);
  wire s1959, sub1959, and1959, or1959;
  wire b_inv1959;
  assign b_inv1959 = ~b1959;
  assign s1959  = a1959 ^ b1959 ^ c1959;
  assign sub1959 = a1959 ^ b_inv1959 ^ c1959;
  assign and1959 = a1959 & b1959;
  assign or1959  = a1959 | b1959;
  assign c1960 = (a1959 & b1959) | (a1959 & c1959) | (b1959 & c1959);
  wire c_sub1960;
  assign c_sub1960 = (a1959 & b_inv1959) | (a1959 & c1959) | (b_inv1959 & c1959);
  wire s1960, sub1960, and1960, or1960;
  wire b_inv1960;
  assign b_inv1960 = ~b1960;
  assign s1960  = a1960 ^ b1960 ^ c1960;
  assign sub1960 = a1960 ^ b_inv1960 ^ c1960;
  assign and1960 = a1960 & b1960;
  assign or1960  = a1960 | b1960;
  assign c1961 = (a1960 & b1960) | (a1960 & c1960) | (b1960 & c1960);
  wire c_sub1961;
  assign c_sub1961 = (a1960 & b_inv1960) | (a1960 & c1960) | (b_inv1960 & c1960);
  wire s1961, sub1961, and1961, or1961;
  wire b_inv1961;
  assign b_inv1961 = ~b1961;
  assign s1961  = a1961 ^ b1961 ^ c1961;
  assign sub1961 = a1961 ^ b_inv1961 ^ c1961;
  assign and1961 = a1961 & b1961;
  assign or1961  = a1961 | b1961;
  assign c1962 = (a1961 & b1961) | (a1961 & c1961) | (b1961 & c1961);
  wire c_sub1962;
  assign c_sub1962 = (a1961 & b_inv1961) | (a1961 & c1961) | (b_inv1961 & c1961);
  wire s1962, sub1962, and1962, or1962;
  wire b_inv1962;
  assign b_inv1962 = ~b1962;
  assign s1962  = a1962 ^ b1962 ^ c1962;
  assign sub1962 = a1962 ^ b_inv1962 ^ c1962;
  assign and1962 = a1962 & b1962;
  assign or1962  = a1962 | b1962;
  assign c1963 = (a1962 & b1962) | (a1962 & c1962) | (b1962 & c1962);
  wire c_sub1963;
  assign c_sub1963 = (a1962 & b_inv1962) | (a1962 & c1962) | (b_inv1962 & c1962);
  wire s1963, sub1963, and1963, or1963;
  wire b_inv1963;
  assign b_inv1963 = ~b1963;
  assign s1963  = a1963 ^ b1963 ^ c1963;
  assign sub1963 = a1963 ^ b_inv1963 ^ c1963;
  assign and1963 = a1963 & b1963;
  assign or1963  = a1963 | b1963;
  assign c1964 = (a1963 & b1963) | (a1963 & c1963) | (b1963 & c1963);
  wire c_sub1964;
  assign c_sub1964 = (a1963 & b_inv1963) | (a1963 & c1963) | (b_inv1963 & c1963);
  wire s1964, sub1964, and1964, or1964;
  wire b_inv1964;
  assign b_inv1964 = ~b1964;
  assign s1964  = a1964 ^ b1964 ^ c1964;
  assign sub1964 = a1964 ^ b_inv1964 ^ c1964;
  assign and1964 = a1964 & b1964;
  assign or1964  = a1964 | b1964;
  assign c1965 = (a1964 & b1964) | (a1964 & c1964) | (b1964 & c1964);
  wire c_sub1965;
  assign c_sub1965 = (a1964 & b_inv1964) | (a1964 & c1964) | (b_inv1964 & c1964);
  wire s1965, sub1965, and1965, or1965;
  wire b_inv1965;
  assign b_inv1965 = ~b1965;
  assign s1965  = a1965 ^ b1965 ^ c1965;
  assign sub1965 = a1965 ^ b_inv1965 ^ c1965;
  assign and1965 = a1965 & b1965;
  assign or1965  = a1965 | b1965;
  assign c1966 = (a1965 & b1965) | (a1965 & c1965) | (b1965 & c1965);
  wire c_sub1966;
  assign c_sub1966 = (a1965 & b_inv1965) | (a1965 & c1965) | (b_inv1965 & c1965);
  wire s1966, sub1966, and1966, or1966;
  wire b_inv1966;
  assign b_inv1966 = ~b1966;
  assign s1966  = a1966 ^ b1966 ^ c1966;
  assign sub1966 = a1966 ^ b_inv1966 ^ c1966;
  assign and1966 = a1966 & b1966;
  assign or1966  = a1966 | b1966;
  assign c1967 = (a1966 & b1966) | (a1966 & c1966) | (b1966 & c1966);
  wire c_sub1967;
  assign c_sub1967 = (a1966 & b_inv1966) | (a1966 & c1966) | (b_inv1966 & c1966);
  wire s1967, sub1967, and1967, or1967;
  wire b_inv1967;
  assign b_inv1967 = ~b1967;
  assign s1967  = a1967 ^ b1967 ^ c1967;
  assign sub1967 = a1967 ^ b_inv1967 ^ c1967;
  assign and1967 = a1967 & b1967;
  assign or1967  = a1967 | b1967;
  assign c1968 = (a1967 & b1967) | (a1967 & c1967) | (b1967 & c1967);
  wire c_sub1968;
  assign c_sub1968 = (a1967 & b_inv1967) | (a1967 & c1967) | (b_inv1967 & c1967);
  wire s1968, sub1968, and1968, or1968;
  wire b_inv1968;
  assign b_inv1968 = ~b1968;
  assign s1968  = a1968 ^ b1968 ^ c1968;
  assign sub1968 = a1968 ^ b_inv1968 ^ c1968;
  assign and1968 = a1968 & b1968;
  assign or1968  = a1968 | b1968;
  assign c1969 = (a1968 & b1968) | (a1968 & c1968) | (b1968 & c1968);
  wire c_sub1969;
  assign c_sub1969 = (a1968 & b_inv1968) | (a1968 & c1968) | (b_inv1968 & c1968);
  wire s1969, sub1969, and1969, or1969;
  wire b_inv1969;
  assign b_inv1969 = ~b1969;
  assign s1969  = a1969 ^ b1969 ^ c1969;
  assign sub1969 = a1969 ^ b_inv1969 ^ c1969;
  assign and1969 = a1969 & b1969;
  assign or1969  = a1969 | b1969;
  assign c1970 = (a1969 & b1969) | (a1969 & c1969) | (b1969 & c1969);
  wire c_sub1970;
  assign c_sub1970 = (a1969 & b_inv1969) | (a1969 & c1969) | (b_inv1969 & c1969);
  wire s1970, sub1970, and1970, or1970;
  wire b_inv1970;
  assign b_inv1970 = ~b1970;
  assign s1970  = a1970 ^ b1970 ^ c1970;
  assign sub1970 = a1970 ^ b_inv1970 ^ c1970;
  assign and1970 = a1970 & b1970;
  assign or1970  = a1970 | b1970;
  assign c1971 = (a1970 & b1970) | (a1970 & c1970) | (b1970 & c1970);
  wire c_sub1971;
  assign c_sub1971 = (a1970 & b_inv1970) | (a1970 & c1970) | (b_inv1970 & c1970);
  wire s1971, sub1971, and1971, or1971;
  wire b_inv1971;
  assign b_inv1971 = ~b1971;
  assign s1971  = a1971 ^ b1971 ^ c1971;
  assign sub1971 = a1971 ^ b_inv1971 ^ c1971;
  assign and1971 = a1971 & b1971;
  assign or1971  = a1971 | b1971;
  assign c1972 = (a1971 & b1971) | (a1971 & c1971) | (b1971 & c1971);
  wire c_sub1972;
  assign c_sub1972 = (a1971 & b_inv1971) | (a1971 & c1971) | (b_inv1971 & c1971);
  wire s1972, sub1972, and1972, or1972;
  wire b_inv1972;
  assign b_inv1972 = ~b1972;
  assign s1972  = a1972 ^ b1972 ^ c1972;
  assign sub1972 = a1972 ^ b_inv1972 ^ c1972;
  assign and1972 = a1972 & b1972;
  assign or1972  = a1972 | b1972;
  assign c1973 = (a1972 & b1972) | (a1972 & c1972) | (b1972 & c1972);
  wire c_sub1973;
  assign c_sub1973 = (a1972 & b_inv1972) | (a1972 & c1972) | (b_inv1972 & c1972);
  wire s1973, sub1973, and1973, or1973;
  wire b_inv1973;
  assign b_inv1973 = ~b1973;
  assign s1973  = a1973 ^ b1973 ^ c1973;
  assign sub1973 = a1973 ^ b_inv1973 ^ c1973;
  assign and1973 = a1973 & b1973;
  assign or1973  = a1973 | b1973;
  assign c1974 = (a1973 & b1973) | (a1973 & c1973) | (b1973 & c1973);
  wire c_sub1974;
  assign c_sub1974 = (a1973 & b_inv1973) | (a1973 & c1973) | (b_inv1973 & c1973);
  wire s1974, sub1974, and1974, or1974;
  wire b_inv1974;
  assign b_inv1974 = ~b1974;
  assign s1974  = a1974 ^ b1974 ^ c1974;
  assign sub1974 = a1974 ^ b_inv1974 ^ c1974;
  assign and1974 = a1974 & b1974;
  assign or1974  = a1974 | b1974;
  assign c1975 = (a1974 & b1974) | (a1974 & c1974) | (b1974 & c1974);
  wire c_sub1975;
  assign c_sub1975 = (a1974 & b_inv1974) | (a1974 & c1974) | (b_inv1974 & c1974);
  wire s1975, sub1975, and1975, or1975;
  wire b_inv1975;
  assign b_inv1975 = ~b1975;
  assign s1975  = a1975 ^ b1975 ^ c1975;
  assign sub1975 = a1975 ^ b_inv1975 ^ c1975;
  assign and1975 = a1975 & b1975;
  assign or1975  = a1975 | b1975;
  assign c1976 = (a1975 & b1975) | (a1975 & c1975) | (b1975 & c1975);
  wire c_sub1976;
  assign c_sub1976 = (a1975 & b_inv1975) | (a1975 & c1975) | (b_inv1975 & c1975);
  wire s1976, sub1976, and1976, or1976;
  wire b_inv1976;
  assign b_inv1976 = ~b1976;
  assign s1976  = a1976 ^ b1976 ^ c1976;
  assign sub1976 = a1976 ^ b_inv1976 ^ c1976;
  assign and1976 = a1976 & b1976;
  assign or1976  = a1976 | b1976;
  assign c1977 = (a1976 & b1976) | (a1976 & c1976) | (b1976 & c1976);
  wire c_sub1977;
  assign c_sub1977 = (a1976 & b_inv1976) | (a1976 & c1976) | (b_inv1976 & c1976);
  wire s1977, sub1977, and1977, or1977;
  wire b_inv1977;
  assign b_inv1977 = ~b1977;
  assign s1977  = a1977 ^ b1977 ^ c1977;
  assign sub1977 = a1977 ^ b_inv1977 ^ c1977;
  assign and1977 = a1977 & b1977;
  assign or1977  = a1977 | b1977;
  assign c1978 = (a1977 & b1977) | (a1977 & c1977) | (b1977 & c1977);
  wire c_sub1978;
  assign c_sub1978 = (a1977 & b_inv1977) | (a1977 & c1977) | (b_inv1977 & c1977);
  wire s1978, sub1978, and1978, or1978;
  wire b_inv1978;
  assign b_inv1978 = ~b1978;
  assign s1978  = a1978 ^ b1978 ^ c1978;
  assign sub1978 = a1978 ^ b_inv1978 ^ c1978;
  assign and1978 = a1978 & b1978;
  assign or1978  = a1978 | b1978;
  assign c1979 = (a1978 & b1978) | (a1978 & c1978) | (b1978 & c1978);
  wire c_sub1979;
  assign c_sub1979 = (a1978 & b_inv1978) | (a1978 & c1978) | (b_inv1978 & c1978);
  wire s1979, sub1979, and1979, or1979;
  wire b_inv1979;
  assign b_inv1979 = ~b1979;
  assign s1979  = a1979 ^ b1979 ^ c1979;
  assign sub1979 = a1979 ^ b_inv1979 ^ c1979;
  assign and1979 = a1979 & b1979;
  assign or1979  = a1979 | b1979;
  assign c1980 = (a1979 & b1979) | (a1979 & c1979) | (b1979 & c1979);
  wire c_sub1980;
  assign c_sub1980 = (a1979 & b_inv1979) | (a1979 & c1979) | (b_inv1979 & c1979);
  wire s1980, sub1980, and1980, or1980;
  wire b_inv1980;
  assign b_inv1980 = ~b1980;
  assign s1980  = a1980 ^ b1980 ^ c1980;
  assign sub1980 = a1980 ^ b_inv1980 ^ c1980;
  assign and1980 = a1980 & b1980;
  assign or1980  = a1980 | b1980;
  assign c1981 = (a1980 & b1980) | (a1980 & c1980) | (b1980 & c1980);
  wire c_sub1981;
  assign c_sub1981 = (a1980 & b_inv1980) | (a1980 & c1980) | (b_inv1980 & c1980);
  wire s1981, sub1981, and1981, or1981;
  wire b_inv1981;
  assign b_inv1981 = ~b1981;
  assign s1981  = a1981 ^ b1981 ^ c1981;
  assign sub1981 = a1981 ^ b_inv1981 ^ c1981;
  assign and1981 = a1981 & b1981;
  assign or1981  = a1981 | b1981;
  assign c1982 = (a1981 & b1981) | (a1981 & c1981) | (b1981 & c1981);
  wire c_sub1982;
  assign c_sub1982 = (a1981 & b_inv1981) | (a1981 & c1981) | (b_inv1981 & c1981);
  wire s1982, sub1982, and1982, or1982;
  wire b_inv1982;
  assign b_inv1982 = ~b1982;
  assign s1982  = a1982 ^ b1982 ^ c1982;
  assign sub1982 = a1982 ^ b_inv1982 ^ c1982;
  assign and1982 = a1982 & b1982;
  assign or1982  = a1982 | b1982;
  assign c1983 = (a1982 & b1982) | (a1982 & c1982) | (b1982 & c1982);
  wire c_sub1983;
  assign c_sub1983 = (a1982 & b_inv1982) | (a1982 & c1982) | (b_inv1982 & c1982);
  wire s1983, sub1983, and1983, or1983;
  wire b_inv1983;
  assign b_inv1983 = ~b1983;
  assign s1983  = a1983 ^ b1983 ^ c1983;
  assign sub1983 = a1983 ^ b_inv1983 ^ c1983;
  assign and1983 = a1983 & b1983;
  assign or1983  = a1983 | b1983;
  assign c1984 = (a1983 & b1983) | (a1983 & c1983) | (b1983 & c1983);
  wire c_sub1984;
  assign c_sub1984 = (a1983 & b_inv1983) | (a1983 & c1983) | (b_inv1983 & c1983);
  wire s1984, sub1984, and1984, or1984;
  wire b_inv1984;
  assign b_inv1984 = ~b1984;
  assign s1984  = a1984 ^ b1984 ^ c1984;
  assign sub1984 = a1984 ^ b_inv1984 ^ c1984;
  assign and1984 = a1984 & b1984;
  assign or1984  = a1984 | b1984;
  assign c1985 = (a1984 & b1984) | (a1984 & c1984) | (b1984 & c1984);
  wire c_sub1985;
  assign c_sub1985 = (a1984 & b_inv1984) | (a1984 & c1984) | (b_inv1984 & c1984);
  wire s1985, sub1985, and1985, or1985;
  wire b_inv1985;
  assign b_inv1985 = ~b1985;
  assign s1985  = a1985 ^ b1985 ^ c1985;
  assign sub1985 = a1985 ^ b_inv1985 ^ c1985;
  assign and1985 = a1985 & b1985;
  assign or1985  = a1985 | b1985;
  assign c1986 = (a1985 & b1985) | (a1985 & c1985) | (b1985 & c1985);
  wire c_sub1986;
  assign c_sub1986 = (a1985 & b_inv1985) | (a1985 & c1985) | (b_inv1985 & c1985);
  wire s1986, sub1986, and1986, or1986;
  wire b_inv1986;
  assign b_inv1986 = ~b1986;
  assign s1986  = a1986 ^ b1986 ^ c1986;
  assign sub1986 = a1986 ^ b_inv1986 ^ c1986;
  assign and1986 = a1986 & b1986;
  assign or1986  = a1986 | b1986;
  assign c1987 = (a1986 & b1986) | (a1986 & c1986) | (b1986 & c1986);
  wire c_sub1987;
  assign c_sub1987 = (a1986 & b_inv1986) | (a1986 & c1986) | (b_inv1986 & c1986);
  wire s1987, sub1987, and1987, or1987;
  wire b_inv1987;
  assign b_inv1987 = ~b1987;
  assign s1987  = a1987 ^ b1987 ^ c1987;
  assign sub1987 = a1987 ^ b_inv1987 ^ c1987;
  assign and1987 = a1987 & b1987;
  assign or1987  = a1987 | b1987;
  assign c1988 = (a1987 & b1987) | (a1987 & c1987) | (b1987 & c1987);
  wire c_sub1988;
  assign c_sub1988 = (a1987 & b_inv1987) | (a1987 & c1987) | (b_inv1987 & c1987);
  wire s1988, sub1988, and1988, or1988;
  wire b_inv1988;
  assign b_inv1988 = ~b1988;
  assign s1988  = a1988 ^ b1988 ^ c1988;
  assign sub1988 = a1988 ^ b_inv1988 ^ c1988;
  assign and1988 = a1988 & b1988;
  assign or1988  = a1988 | b1988;
  assign c1989 = (a1988 & b1988) | (a1988 & c1988) | (b1988 & c1988);
  wire c_sub1989;
  assign c_sub1989 = (a1988 & b_inv1988) | (a1988 & c1988) | (b_inv1988 & c1988);
  wire s1989, sub1989, and1989, or1989;
  wire b_inv1989;
  assign b_inv1989 = ~b1989;
  assign s1989  = a1989 ^ b1989 ^ c1989;
  assign sub1989 = a1989 ^ b_inv1989 ^ c1989;
  assign and1989 = a1989 & b1989;
  assign or1989  = a1989 | b1989;
  assign c1990 = (a1989 & b1989) | (a1989 & c1989) | (b1989 & c1989);
  wire c_sub1990;
  assign c_sub1990 = (a1989 & b_inv1989) | (a1989 & c1989) | (b_inv1989 & c1989);
  wire s1990, sub1990, and1990, or1990;
  wire b_inv1990;
  assign b_inv1990 = ~b1990;
  assign s1990  = a1990 ^ b1990 ^ c1990;
  assign sub1990 = a1990 ^ b_inv1990 ^ c1990;
  assign and1990 = a1990 & b1990;
  assign or1990  = a1990 | b1990;
  assign c1991 = (a1990 & b1990) | (a1990 & c1990) | (b1990 & c1990);
  wire c_sub1991;
  assign c_sub1991 = (a1990 & b_inv1990) | (a1990 & c1990) | (b_inv1990 & c1990);
  wire s1991, sub1991, and1991, or1991;
  wire b_inv1991;
  assign b_inv1991 = ~b1991;
  assign s1991  = a1991 ^ b1991 ^ c1991;
  assign sub1991 = a1991 ^ b_inv1991 ^ c1991;
  assign and1991 = a1991 & b1991;
  assign or1991  = a1991 | b1991;
  assign c1992 = (a1991 & b1991) | (a1991 & c1991) | (b1991 & c1991);
  wire c_sub1992;
  assign c_sub1992 = (a1991 & b_inv1991) | (a1991 & c1991) | (b_inv1991 & c1991);
  wire s1992, sub1992, and1992, or1992;
  wire b_inv1992;
  assign b_inv1992 = ~b1992;
  assign s1992  = a1992 ^ b1992 ^ c1992;
  assign sub1992 = a1992 ^ b_inv1992 ^ c1992;
  assign and1992 = a1992 & b1992;
  assign or1992  = a1992 | b1992;
  assign c1993 = (a1992 & b1992) | (a1992 & c1992) | (b1992 & c1992);
  wire c_sub1993;
  assign c_sub1993 = (a1992 & b_inv1992) | (a1992 & c1992) | (b_inv1992 & c1992);
  wire s1993, sub1993, and1993, or1993;
  wire b_inv1993;
  assign b_inv1993 = ~b1993;
  assign s1993  = a1993 ^ b1993 ^ c1993;
  assign sub1993 = a1993 ^ b_inv1993 ^ c1993;
  assign and1993 = a1993 & b1993;
  assign or1993  = a1993 | b1993;
  assign c1994 = (a1993 & b1993) | (a1993 & c1993) | (b1993 & c1993);
  wire c_sub1994;
  assign c_sub1994 = (a1993 & b_inv1993) | (a1993 & c1993) | (b_inv1993 & c1993);
  wire s1994, sub1994, and1994, or1994;
  wire b_inv1994;
  assign b_inv1994 = ~b1994;
  assign s1994  = a1994 ^ b1994 ^ c1994;
  assign sub1994 = a1994 ^ b_inv1994 ^ c1994;
  assign and1994 = a1994 & b1994;
  assign or1994  = a1994 | b1994;
  assign c1995 = (a1994 & b1994) | (a1994 & c1994) | (b1994 & c1994);
  wire c_sub1995;
  assign c_sub1995 = (a1994 & b_inv1994) | (a1994 & c1994) | (b_inv1994 & c1994);
  wire s1995, sub1995, and1995, or1995;
  wire b_inv1995;
  assign b_inv1995 = ~b1995;
  assign s1995  = a1995 ^ b1995 ^ c1995;
  assign sub1995 = a1995 ^ b_inv1995 ^ c1995;
  assign and1995 = a1995 & b1995;
  assign or1995  = a1995 | b1995;
  assign c1996 = (a1995 & b1995) | (a1995 & c1995) | (b1995 & c1995);
  wire c_sub1996;
  assign c_sub1996 = (a1995 & b_inv1995) | (a1995 & c1995) | (b_inv1995 & c1995);
  wire s1996, sub1996, and1996, or1996;
  wire b_inv1996;
  assign b_inv1996 = ~b1996;
  assign s1996  = a1996 ^ b1996 ^ c1996;
  assign sub1996 = a1996 ^ b_inv1996 ^ c1996;
  assign and1996 = a1996 & b1996;
  assign or1996  = a1996 | b1996;
  assign c1997 = (a1996 & b1996) | (a1996 & c1996) | (b1996 & c1996);
  wire c_sub1997;
  assign c_sub1997 = (a1996 & b_inv1996) | (a1996 & c1996) | (b_inv1996 & c1996);
  wire s1997, sub1997, and1997, or1997;
  wire b_inv1997;
  assign b_inv1997 = ~b1997;
  assign s1997  = a1997 ^ b1997 ^ c1997;
  assign sub1997 = a1997 ^ b_inv1997 ^ c1997;
  assign and1997 = a1997 & b1997;
  assign or1997  = a1997 | b1997;
  assign c1998 = (a1997 & b1997) | (a1997 & c1997) | (b1997 & c1997);
  wire c_sub1998;
  assign c_sub1998 = (a1997 & b_inv1997) | (a1997 & c1997) | (b_inv1997 & c1997);
  wire s1998, sub1998, and1998, or1998;
  wire b_inv1998;
  assign b_inv1998 = ~b1998;
  assign s1998  = a1998 ^ b1998 ^ c1998;
  assign sub1998 = a1998 ^ b_inv1998 ^ c1998;
  assign and1998 = a1998 & b1998;
  assign or1998  = a1998 | b1998;
  assign c1999 = (a1998 & b1998) | (a1998 & c1998) | (b1998 & c1998);
  wire c_sub1999;
  assign c_sub1999 = (a1998 & b_inv1998) | (a1998 & c1998) | (b_inv1998 & c1998);
  wire s1999, sub1999, and1999, or1999;
  wire b_inv1999;
  assign b_inv1999 = ~b1999;
  assign s1999  = a1999 ^ b1999 ^ c1999;
  assign sub1999 = a1999 ^ b_inv1999 ^ c1999;
  assign and1999 = a1999 & b1999;
  assign or1999  = a1999 | b1999;
  assign c2000 = (a1999 & b1999) | (a1999 & c1999) | (b1999 & c1999);
  wire c_sub2000;
  assign c_sub2000 = (a1999 & b_inv1999) | (a1999 & c1999) | (b_inv1999 & c1999);
  wire s2000, sub2000, and2000, or2000;
  wire b_inv2000;
  assign b_inv2000 = ~b2000;
  assign s2000  = a2000 ^ b2000 ^ c2000;
  assign sub2000 = a2000 ^ b_inv2000 ^ c2000;
  assign and2000 = a2000 & b2000;
  assign or2000  = a2000 | b2000;
  assign c2001 = (a2000 & b2000) | (a2000 & c2000) | (b2000 & c2000);
  wire c_sub2001;
  assign c_sub2001 = (a2000 & b_inv2000) | (a2000 & c2000) | (b_inv2000 & c2000);
  wire s2001, sub2001, and2001, or2001;
  wire b_inv2001;
  assign b_inv2001 = ~b2001;
  assign s2001  = a2001 ^ b2001 ^ c2001;
  assign sub2001 = a2001 ^ b_inv2001 ^ c2001;
  assign and2001 = a2001 & b2001;
  assign or2001  = a2001 | b2001;
  assign c2002 = (a2001 & b2001) | (a2001 & c2001) | (b2001 & c2001);
  wire c_sub2002;
  assign c_sub2002 = (a2001 & b_inv2001) | (a2001 & c2001) | (b_inv2001 & c2001);
  wire s2002, sub2002, and2002, or2002;
  wire b_inv2002;
  assign b_inv2002 = ~b2002;
  assign s2002  = a2002 ^ b2002 ^ c2002;
  assign sub2002 = a2002 ^ b_inv2002 ^ c2002;
  assign and2002 = a2002 & b2002;
  assign or2002  = a2002 | b2002;
  assign c2003 = (a2002 & b2002) | (a2002 & c2002) | (b2002 & c2002);
  wire c_sub2003;
  assign c_sub2003 = (a2002 & b_inv2002) | (a2002 & c2002) | (b_inv2002 & c2002);
  wire s2003, sub2003, and2003, or2003;
  wire b_inv2003;
  assign b_inv2003 = ~b2003;
  assign s2003  = a2003 ^ b2003 ^ c2003;
  assign sub2003 = a2003 ^ b_inv2003 ^ c2003;
  assign and2003 = a2003 & b2003;
  assign or2003  = a2003 | b2003;
  assign c2004 = (a2003 & b2003) | (a2003 & c2003) | (b2003 & c2003);
  wire c_sub2004;
  assign c_sub2004 = (a2003 & b_inv2003) | (a2003 & c2003) | (b_inv2003 & c2003);
  wire s2004, sub2004, and2004, or2004;
  wire b_inv2004;
  assign b_inv2004 = ~b2004;
  assign s2004  = a2004 ^ b2004 ^ c2004;
  assign sub2004 = a2004 ^ b_inv2004 ^ c2004;
  assign and2004 = a2004 & b2004;
  assign or2004  = a2004 | b2004;
  assign c2005 = (a2004 & b2004) | (a2004 & c2004) | (b2004 & c2004);
  wire c_sub2005;
  assign c_sub2005 = (a2004 & b_inv2004) | (a2004 & c2004) | (b_inv2004 & c2004);
  wire s2005, sub2005, and2005, or2005;
  wire b_inv2005;
  assign b_inv2005 = ~b2005;
  assign s2005  = a2005 ^ b2005 ^ c2005;
  assign sub2005 = a2005 ^ b_inv2005 ^ c2005;
  assign and2005 = a2005 & b2005;
  assign or2005  = a2005 | b2005;
  assign c2006 = (a2005 & b2005) | (a2005 & c2005) | (b2005 & c2005);
  wire c_sub2006;
  assign c_sub2006 = (a2005 & b_inv2005) | (a2005 & c2005) | (b_inv2005 & c2005);
  wire s2006, sub2006, and2006, or2006;
  wire b_inv2006;
  assign b_inv2006 = ~b2006;
  assign s2006  = a2006 ^ b2006 ^ c2006;
  assign sub2006 = a2006 ^ b_inv2006 ^ c2006;
  assign and2006 = a2006 & b2006;
  assign or2006  = a2006 | b2006;
  assign c2007 = (a2006 & b2006) | (a2006 & c2006) | (b2006 & c2006);
  wire c_sub2007;
  assign c_sub2007 = (a2006 & b_inv2006) | (a2006 & c2006) | (b_inv2006 & c2006);
  wire s2007, sub2007, and2007, or2007;
  wire b_inv2007;
  assign b_inv2007 = ~b2007;
  assign s2007  = a2007 ^ b2007 ^ c2007;
  assign sub2007 = a2007 ^ b_inv2007 ^ c2007;
  assign and2007 = a2007 & b2007;
  assign or2007  = a2007 | b2007;
  assign c2008 = (a2007 & b2007) | (a2007 & c2007) | (b2007 & c2007);
  wire c_sub2008;
  assign c_sub2008 = (a2007 & b_inv2007) | (a2007 & c2007) | (b_inv2007 & c2007);
  wire s2008, sub2008, and2008, or2008;
  wire b_inv2008;
  assign b_inv2008 = ~b2008;
  assign s2008  = a2008 ^ b2008 ^ c2008;
  assign sub2008 = a2008 ^ b_inv2008 ^ c2008;
  assign and2008 = a2008 & b2008;
  assign or2008  = a2008 | b2008;
  assign c2009 = (a2008 & b2008) | (a2008 & c2008) | (b2008 & c2008);
  wire c_sub2009;
  assign c_sub2009 = (a2008 & b_inv2008) | (a2008 & c2008) | (b_inv2008 & c2008);
  wire s2009, sub2009, and2009, or2009;
  wire b_inv2009;
  assign b_inv2009 = ~b2009;
  assign s2009  = a2009 ^ b2009 ^ c2009;
  assign sub2009 = a2009 ^ b_inv2009 ^ c2009;
  assign and2009 = a2009 & b2009;
  assign or2009  = a2009 | b2009;
  assign c2010 = (a2009 & b2009) | (a2009 & c2009) | (b2009 & c2009);
  wire c_sub2010;
  assign c_sub2010 = (a2009 & b_inv2009) | (a2009 & c2009) | (b_inv2009 & c2009);
  wire s2010, sub2010, and2010, or2010;
  wire b_inv2010;
  assign b_inv2010 = ~b2010;
  assign s2010  = a2010 ^ b2010 ^ c2010;
  assign sub2010 = a2010 ^ b_inv2010 ^ c2010;
  assign and2010 = a2010 & b2010;
  assign or2010  = a2010 | b2010;
  assign c2011 = (a2010 & b2010) | (a2010 & c2010) | (b2010 & c2010);
  wire c_sub2011;
  assign c_sub2011 = (a2010 & b_inv2010) | (a2010 & c2010) | (b_inv2010 & c2010);
  wire s2011, sub2011, and2011, or2011;
  wire b_inv2011;
  assign b_inv2011 = ~b2011;
  assign s2011  = a2011 ^ b2011 ^ c2011;
  assign sub2011 = a2011 ^ b_inv2011 ^ c2011;
  assign and2011 = a2011 & b2011;
  assign or2011  = a2011 | b2011;
  assign c2012 = (a2011 & b2011) | (a2011 & c2011) | (b2011 & c2011);
  wire c_sub2012;
  assign c_sub2012 = (a2011 & b_inv2011) | (a2011 & c2011) | (b_inv2011 & c2011);
  wire s2012, sub2012, and2012, or2012;
  wire b_inv2012;
  assign b_inv2012 = ~b2012;
  assign s2012  = a2012 ^ b2012 ^ c2012;
  assign sub2012 = a2012 ^ b_inv2012 ^ c2012;
  assign and2012 = a2012 & b2012;
  assign or2012  = a2012 | b2012;
  assign c2013 = (a2012 & b2012) | (a2012 & c2012) | (b2012 & c2012);
  wire c_sub2013;
  assign c_sub2013 = (a2012 & b_inv2012) | (a2012 & c2012) | (b_inv2012 & c2012);
  wire s2013, sub2013, and2013, or2013;
  wire b_inv2013;
  assign b_inv2013 = ~b2013;
  assign s2013  = a2013 ^ b2013 ^ c2013;
  assign sub2013 = a2013 ^ b_inv2013 ^ c2013;
  assign and2013 = a2013 & b2013;
  assign or2013  = a2013 | b2013;
  assign c2014 = (a2013 & b2013) | (a2013 & c2013) | (b2013 & c2013);
  wire c_sub2014;
  assign c_sub2014 = (a2013 & b_inv2013) | (a2013 & c2013) | (b_inv2013 & c2013);
  wire s2014, sub2014, and2014, or2014;
  wire b_inv2014;
  assign b_inv2014 = ~b2014;
  assign s2014  = a2014 ^ b2014 ^ c2014;
  assign sub2014 = a2014 ^ b_inv2014 ^ c2014;
  assign and2014 = a2014 & b2014;
  assign or2014  = a2014 | b2014;
  assign c2015 = (a2014 & b2014) | (a2014 & c2014) | (b2014 & c2014);
  wire c_sub2015;
  assign c_sub2015 = (a2014 & b_inv2014) | (a2014 & c2014) | (b_inv2014 & c2014);
  wire s2015, sub2015, and2015, or2015;
  wire b_inv2015;
  assign b_inv2015 = ~b2015;
  assign s2015  = a2015 ^ b2015 ^ c2015;
  assign sub2015 = a2015 ^ b_inv2015 ^ c2015;
  assign and2015 = a2015 & b2015;
  assign or2015  = a2015 | b2015;
  assign c2016 = (a2015 & b2015) | (a2015 & c2015) | (b2015 & c2015);
  wire c_sub2016;
  assign c_sub2016 = (a2015 & b_inv2015) | (a2015 & c2015) | (b_inv2015 & c2015);
  wire s2016, sub2016, and2016, or2016;
  wire b_inv2016;
  assign b_inv2016 = ~b2016;
  assign s2016  = a2016 ^ b2016 ^ c2016;
  assign sub2016 = a2016 ^ b_inv2016 ^ c2016;
  assign and2016 = a2016 & b2016;
  assign or2016  = a2016 | b2016;
  assign c2017 = (a2016 & b2016) | (a2016 & c2016) | (b2016 & c2016);
  wire c_sub2017;
  assign c_sub2017 = (a2016 & b_inv2016) | (a2016 & c2016) | (b_inv2016 & c2016);
  wire s2017, sub2017, and2017, or2017;
  wire b_inv2017;
  assign b_inv2017 = ~b2017;
  assign s2017  = a2017 ^ b2017 ^ c2017;
  assign sub2017 = a2017 ^ b_inv2017 ^ c2017;
  assign and2017 = a2017 & b2017;
  assign or2017  = a2017 | b2017;
  assign c2018 = (a2017 & b2017) | (a2017 & c2017) | (b2017 & c2017);
  wire c_sub2018;
  assign c_sub2018 = (a2017 & b_inv2017) | (a2017 & c2017) | (b_inv2017 & c2017);
  wire s2018, sub2018, and2018, or2018;
  wire b_inv2018;
  assign b_inv2018 = ~b2018;
  assign s2018  = a2018 ^ b2018 ^ c2018;
  assign sub2018 = a2018 ^ b_inv2018 ^ c2018;
  assign and2018 = a2018 & b2018;
  assign or2018  = a2018 | b2018;
  assign c2019 = (a2018 & b2018) | (a2018 & c2018) | (b2018 & c2018);
  wire c_sub2019;
  assign c_sub2019 = (a2018 & b_inv2018) | (a2018 & c2018) | (b_inv2018 & c2018);
  wire s2019, sub2019, and2019, or2019;
  wire b_inv2019;
  assign b_inv2019 = ~b2019;
  assign s2019  = a2019 ^ b2019 ^ c2019;
  assign sub2019 = a2019 ^ b_inv2019 ^ c2019;
  assign and2019 = a2019 & b2019;
  assign or2019  = a2019 | b2019;
  assign c2020 = (a2019 & b2019) | (a2019 & c2019) | (b2019 & c2019);
  wire c_sub2020;
  assign c_sub2020 = (a2019 & b_inv2019) | (a2019 & c2019) | (b_inv2019 & c2019);
  wire s2020, sub2020, and2020, or2020;
  wire b_inv2020;
  assign b_inv2020 = ~b2020;
  assign s2020  = a2020 ^ b2020 ^ c2020;
  assign sub2020 = a2020 ^ b_inv2020 ^ c2020;
  assign and2020 = a2020 & b2020;
  assign or2020  = a2020 | b2020;
  assign c2021 = (a2020 & b2020) | (a2020 & c2020) | (b2020 & c2020);
  wire c_sub2021;
  assign c_sub2021 = (a2020 & b_inv2020) | (a2020 & c2020) | (b_inv2020 & c2020);
  wire s2021, sub2021, and2021, or2021;
  wire b_inv2021;
  assign b_inv2021 = ~b2021;
  assign s2021  = a2021 ^ b2021 ^ c2021;
  assign sub2021 = a2021 ^ b_inv2021 ^ c2021;
  assign and2021 = a2021 & b2021;
  assign or2021  = a2021 | b2021;
  assign c2022 = (a2021 & b2021) | (a2021 & c2021) | (b2021 & c2021);
  wire c_sub2022;
  assign c_sub2022 = (a2021 & b_inv2021) | (a2021 & c2021) | (b_inv2021 & c2021);
  wire s2022, sub2022, and2022, or2022;
  wire b_inv2022;
  assign b_inv2022 = ~b2022;
  assign s2022  = a2022 ^ b2022 ^ c2022;
  assign sub2022 = a2022 ^ b_inv2022 ^ c2022;
  assign and2022 = a2022 & b2022;
  assign or2022  = a2022 | b2022;
  assign c2023 = (a2022 & b2022) | (a2022 & c2022) | (b2022 & c2022);
  wire c_sub2023;
  assign c_sub2023 = (a2022 & b_inv2022) | (a2022 & c2022) | (b_inv2022 & c2022);
  wire s2023, sub2023, and2023, or2023;
  wire b_inv2023;
  assign b_inv2023 = ~b2023;
  assign s2023  = a2023 ^ b2023 ^ c2023;
  assign sub2023 = a2023 ^ b_inv2023 ^ c2023;
  assign and2023 = a2023 & b2023;
  assign or2023  = a2023 | b2023;
  assign c2024 = (a2023 & b2023) | (a2023 & c2023) | (b2023 & c2023);
  wire c_sub2024;
  assign c_sub2024 = (a2023 & b_inv2023) | (a2023 & c2023) | (b_inv2023 & c2023);
  wire s2024, sub2024, and2024, or2024;
  wire b_inv2024;
  assign b_inv2024 = ~b2024;
  assign s2024  = a2024 ^ b2024 ^ c2024;
  assign sub2024 = a2024 ^ b_inv2024 ^ c2024;
  assign and2024 = a2024 & b2024;
  assign or2024  = a2024 | b2024;
  assign c2025 = (a2024 & b2024) | (a2024 & c2024) | (b2024 & c2024);
  wire c_sub2025;
  assign c_sub2025 = (a2024 & b_inv2024) | (a2024 & c2024) | (b_inv2024 & c2024);
  wire s2025, sub2025, and2025, or2025;
  wire b_inv2025;
  assign b_inv2025 = ~b2025;
  assign s2025  = a2025 ^ b2025 ^ c2025;
  assign sub2025 = a2025 ^ b_inv2025 ^ c2025;
  assign and2025 = a2025 & b2025;
  assign or2025  = a2025 | b2025;
  assign c2026 = (a2025 & b2025) | (a2025 & c2025) | (b2025 & c2025);
  wire c_sub2026;
  assign c_sub2026 = (a2025 & b_inv2025) | (a2025 & c2025) | (b_inv2025 & c2025);
  wire s2026, sub2026, and2026, or2026;
  wire b_inv2026;
  assign b_inv2026 = ~b2026;
  assign s2026  = a2026 ^ b2026 ^ c2026;
  assign sub2026 = a2026 ^ b_inv2026 ^ c2026;
  assign and2026 = a2026 & b2026;
  assign or2026  = a2026 | b2026;
  assign c2027 = (a2026 & b2026) | (a2026 & c2026) | (b2026 & c2026);
  wire c_sub2027;
  assign c_sub2027 = (a2026 & b_inv2026) | (a2026 & c2026) | (b_inv2026 & c2026);
  wire s2027, sub2027, and2027, or2027;
  wire b_inv2027;
  assign b_inv2027 = ~b2027;
  assign s2027  = a2027 ^ b2027 ^ c2027;
  assign sub2027 = a2027 ^ b_inv2027 ^ c2027;
  assign and2027 = a2027 & b2027;
  assign or2027  = a2027 | b2027;
  assign c2028 = (a2027 & b2027) | (a2027 & c2027) | (b2027 & c2027);
  wire c_sub2028;
  assign c_sub2028 = (a2027 & b_inv2027) | (a2027 & c2027) | (b_inv2027 & c2027);
  wire s2028, sub2028, and2028, or2028;
  wire b_inv2028;
  assign b_inv2028 = ~b2028;
  assign s2028  = a2028 ^ b2028 ^ c2028;
  assign sub2028 = a2028 ^ b_inv2028 ^ c2028;
  assign and2028 = a2028 & b2028;
  assign or2028  = a2028 | b2028;
  assign c2029 = (a2028 & b2028) | (a2028 & c2028) | (b2028 & c2028);
  wire c_sub2029;
  assign c_sub2029 = (a2028 & b_inv2028) | (a2028 & c2028) | (b_inv2028 & c2028);
  wire s2029, sub2029, and2029, or2029;
  wire b_inv2029;
  assign b_inv2029 = ~b2029;
  assign s2029  = a2029 ^ b2029 ^ c2029;
  assign sub2029 = a2029 ^ b_inv2029 ^ c2029;
  assign and2029 = a2029 & b2029;
  assign or2029  = a2029 | b2029;
  assign c2030 = (a2029 & b2029) | (a2029 & c2029) | (b2029 & c2029);
  wire c_sub2030;
  assign c_sub2030 = (a2029 & b_inv2029) | (a2029 & c2029) | (b_inv2029 & c2029);
  wire s2030, sub2030, and2030, or2030;
  wire b_inv2030;
  assign b_inv2030 = ~b2030;
  assign s2030  = a2030 ^ b2030 ^ c2030;
  assign sub2030 = a2030 ^ b_inv2030 ^ c2030;
  assign and2030 = a2030 & b2030;
  assign or2030  = a2030 | b2030;
  assign c2031 = (a2030 & b2030) | (a2030 & c2030) | (b2030 & c2030);
  wire c_sub2031;
  assign c_sub2031 = (a2030 & b_inv2030) | (a2030 & c2030) | (b_inv2030 & c2030);
  wire s2031, sub2031, and2031, or2031;
  wire b_inv2031;
  assign b_inv2031 = ~b2031;
  assign s2031  = a2031 ^ b2031 ^ c2031;
  assign sub2031 = a2031 ^ b_inv2031 ^ c2031;
  assign and2031 = a2031 & b2031;
  assign or2031  = a2031 | b2031;
  assign c2032 = (a2031 & b2031) | (a2031 & c2031) | (b2031 & c2031);
  wire c_sub2032;
  assign c_sub2032 = (a2031 & b_inv2031) | (a2031 & c2031) | (b_inv2031 & c2031);
  wire s2032, sub2032, and2032, or2032;
  wire b_inv2032;
  assign b_inv2032 = ~b2032;
  assign s2032  = a2032 ^ b2032 ^ c2032;
  assign sub2032 = a2032 ^ b_inv2032 ^ c2032;
  assign and2032 = a2032 & b2032;
  assign or2032  = a2032 | b2032;
  assign c2033 = (a2032 & b2032) | (a2032 & c2032) | (b2032 & c2032);
  wire c_sub2033;
  assign c_sub2033 = (a2032 & b_inv2032) | (a2032 & c2032) | (b_inv2032 & c2032);
  wire s2033, sub2033, and2033, or2033;
  wire b_inv2033;
  assign b_inv2033 = ~b2033;
  assign s2033  = a2033 ^ b2033 ^ c2033;
  assign sub2033 = a2033 ^ b_inv2033 ^ c2033;
  assign and2033 = a2033 & b2033;
  assign or2033  = a2033 | b2033;
  assign c2034 = (a2033 & b2033) | (a2033 & c2033) | (b2033 & c2033);
  wire c_sub2034;
  assign c_sub2034 = (a2033 & b_inv2033) | (a2033 & c2033) | (b_inv2033 & c2033);
  wire s2034, sub2034, and2034, or2034;
  wire b_inv2034;
  assign b_inv2034 = ~b2034;
  assign s2034  = a2034 ^ b2034 ^ c2034;
  assign sub2034 = a2034 ^ b_inv2034 ^ c2034;
  assign and2034 = a2034 & b2034;
  assign or2034  = a2034 | b2034;
  assign c2035 = (a2034 & b2034) | (a2034 & c2034) | (b2034 & c2034);
  wire c_sub2035;
  assign c_sub2035 = (a2034 & b_inv2034) | (a2034 & c2034) | (b_inv2034 & c2034);
  wire s2035, sub2035, and2035, or2035;
  wire b_inv2035;
  assign b_inv2035 = ~b2035;
  assign s2035  = a2035 ^ b2035 ^ c2035;
  assign sub2035 = a2035 ^ b_inv2035 ^ c2035;
  assign and2035 = a2035 & b2035;
  assign or2035  = a2035 | b2035;
  assign c2036 = (a2035 & b2035) | (a2035 & c2035) | (b2035 & c2035);
  wire c_sub2036;
  assign c_sub2036 = (a2035 & b_inv2035) | (a2035 & c2035) | (b_inv2035 & c2035);
  wire s2036, sub2036, and2036, or2036;
  wire b_inv2036;
  assign b_inv2036 = ~b2036;
  assign s2036  = a2036 ^ b2036 ^ c2036;
  assign sub2036 = a2036 ^ b_inv2036 ^ c2036;
  assign and2036 = a2036 & b2036;
  assign or2036  = a2036 | b2036;
  assign c2037 = (a2036 & b2036) | (a2036 & c2036) | (b2036 & c2036);
  wire c_sub2037;
  assign c_sub2037 = (a2036 & b_inv2036) | (a2036 & c2036) | (b_inv2036 & c2036);
  wire s2037, sub2037, and2037, or2037;
  wire b_inv2037;
  assign b_inv2037 = ~b2037;
  assign s2037  = a2037 ^ b2037 ^ c2037;
  assign sub2037 = a2037 ^ b_inv2037 ^ c2037;
  assign and2037 = a2037 & b2037;
  assign or2037  = a2037 | b2037;
  assign c2038 = (a2037 & b2037) | (a2037 & c2037) | (b2037 & c2037);
  wire c_sub2038;
  assign c_sub2038 = (a2037 & b_inv2037) | (a2037 & c2037) | (b_inv2037 & c2037);
  wire s2038, sub2038, and2038, or2038;
  wire b_inv2038;
  assign b_inv2038 = ~b2038;
  assign s2038  = a2038 ^ b2038 ^ c2038;
  assign sub2038 = a2038 ^ b_inv2038 ^ c2038;
  assign and2038 = a2038 & b2038;
  assign or2038  = a2038 | b2038;
  assign c2039 = (a2038 & b2038) | (a2038 & c2038) | (b2038 & c2038);
  wire c_sub2039;
  assign c_sub2039 = (a2038 & b_inv2038) | (a2038 & c2038) | (b_inv2038 & c2038);
  wire s2039, sub2039, and2039, or2039;
  wire b_inv2039;
  assign b_inv2039 = ~b2039;
  assign s2039  = a2039 ^ b2039 ^ c2039;
  assign sub2039 = a2039 ^ b_inv2039 ^ c2039;
  assign and2039 = a2039 & b2039;
  assign or2039  = a2039 | b2039;
  assign c2040 = (a2039 & b2039) | (a2039 & c2039) | (b2039 & c2039);
  wire c_sub2040;
  assign c_sub2040 = (a2039 & b_inv2039) | (a2039 & c2039) | (b_inv2039 & c2039);
  wire s2040, sub2040, and2040, or2040;
  wire b_inv2040;
  assign b_inv2040 = ~b2040;
  assign s2040  = a2040 ^ b2040 ^ c2040;
  assign sub2040 = a2040 ^ b_inv2040 ^ c2040;
  assign and2040 = a2040 & b2040;
  assign or2040  = a2040 | b2040;
  assign c2041 = (a2040 & b2040) | (a2040 & c2040) | (b2040 & c2040);
  wire c_sub2041;
  assign c_sub2041 = (a2040 & b_inv2040) | (a2040 & c2040) | (b_inv2040 & c2040);
  wire s2041, sub2041, and2041, or2041;
  wire b_inv2041;
  assign b_inv2041 = ~b2041;
  assign s2041  = a2041 ^ b2041 ^ c2041;
  assign sub2041 = a2041 ^ b_inv2041 ^ c2041;
  assign and2041 = a2041 & b2041;
  assign or2041  = a2041 | b2041;
  assign c2042 = (a2041 & b2041) | (a2041 & c2041) | (b2041 & c2041);
  wire c_sub2042;
  assign c_sub2042 = (a2041 & b_inv2041) | (a2041 & c2041) | (b_inv2041 & c2041);
  wire s2042, sub2042, and2042, or2042;
  wire b_inv2042;
  assign b_inv2042 = ~b2042;
  assign s2042  = a2042 ^ b2042 ^ c2042;
  assign sub2042 = a2042 ^ b_inv2042 ^ c2042;
  assign and2042 = a2042 & b2042;
  assign or2042  = a2042 | b2042;
  assign c2043 = (a2042 & b2042) | (a2042 & c2042) | (b2042 & c2042);
  wire c_sub2043;
  assign c_sub2043 = (a2042 & b_inv2042) | (a2042 & c2042) | (b_inv2042 & c2042);
  wire s2043, sub2043, and2043, or2043;
  wire b_inv2043;
  assign b_inv2043 = ~b2043;
  assign s2043  = a2043 ^ b2043 ^ c2043;
  assign sub2043 = a2043 ^ b_inv2043 ^ c2043;
  assign and2043 = a2043 & b2043;
  assign or2043  = a2043 | b2043;
  assign c2044 = (a2043 & b2043) | (a2043 & c2043) | (b2043 & c2043);
  wire c_sub2044;
  assign c_sub2044 = (a2043 & b_inv2043) | (a2043 & c2043) | (b_inv2043 & c2043);
  wire s2044, sub2044, and2044, or2044;
  wire b_inv2044;
  assign b_inv2044 = ~b2044;
  assign s2044  = a2044 ^ b2044 ^ c2044;
  assign sub2044 = a2044 ^ b_inv2044 ^ c2044;
  assign and2044 = a2044 & b2044;
  assign or2044  = a2044 | b2044;
  assign c2045 = (a2044 & b2044) | (a2044 & c2044) | (b2044 & c2044);
  wire c_sub2045;
  assign c_sub2045 = (a2044 & b_inv2044) | (a2044 & c2044) | (b_inv2044 & c2044);
  wire s2045, sub2045, and2045, or2045;
  wire b_inv2045;
  assign b_inv2045 = ~b2045;
  assign s2045  = a2045 ^ b2045 ^ c2045;
  assign sub2045 = a2045 ^ b_inv2045 ^ c2045;
  assign and2045 = a2045 & b2045;
  assign or2045  = a2045 | b2045;
  assign c2046 = (a2045 & b2045) | (a2045 & c2045) | (b2045 & c2045);
  wire c_sub2046;
  assign c_sub2046 = (a2045 & b_inv2045) | (a2045 & c2045) | (b_inv2045 & c2045);
  wire s2046, sub2046, and2046, or2046;
  wire b_inv2046;
  assign b_inv2046 = ~b2046;
  assign s2046  = a2046 ^ b2046 ^ c2046;
  assign sub2046 = a2046 ^ b_inv2046 ^ c2046;
  assign and2046 = a2046 & b2046;
  assign or2046  = a2046 | b2046;
  assign c2047 = (a2046 & b2046) | (a2046 & c2046) | (b2046 & c2046);
  wire c_sub2047;
  assign c_sub2047 = (a2046 & b_inv2046) | (a2046 & c2046) | (b_inv2046 & c2046);
  wire s2047, sub2047, and2047, or2047;
  wire b_inv2047;
  assign b_inv2047 = ~b2047;
  assign s2047  = a2047 ^ b2047 ^ c2047;
  assign sub2047 = a2047 ^ b_inv2047 ^ c2047;
  assign and2047 = a2047 & b2047;
  assign or2047  = a2047 | b2047;
  assign c2048 = (a2047 & b2047) | (a2047 & c2047) | (b2047 & c2047);
  wire c_sub2048;
  assign c_sub2048 = (a2047 & b_inv2047) | (a2047 & c2047) | (b_inv2047 & c2047);
  assign y0 = (add_sel & s0) | (sub_sel & sub0) | (and_sel & and0) | (or_sel & or0);
  assign y1 = (add_sel & s1) | (sub_sel & sub1) | (and_sel & and1) | (or_sel & or1);
  assign y2 = (add_sel & s2) | (sub_sel & sub2) | (and_sel & and2) | (or_sel & or2);
  assign y3 = (add_sel & s3) | (sub_sel & sub3) | (and_sel & and3) | (or_sel & or3);
  assign y4 = (add_sel & s4) | (sub_sel & sub4) | (and_sel & and4) | (or_sel & or4);
  assign y5 = (add_sel & s5) | (sub_sel & sub5) | (and_sel & and5) | (or_sel & or5);
  assign y6 = (add_sel & s6) | (sub_sel & sub6) | (and_sel & and6) | (or_sel & or6);
  assign y7 = (add_sel & s7) | (sub_sel & sub7) | (and_sel & and7) | (or_sel & or7);
  assign y8 = (add_sel & s8) | (sub_sel & sub8) | (and_sel & and8) | (or_sel & or8);
  assign y9 = (add_sel & s9) | (sub_sel & sub9) | (and_sel & and9) | (or_sel & or9);
  assign y10 = (add_sel & s10) | (sub_sel & sub10) | (and_sel & and10) | (or_sel & or10);
  assign y11 = (add_sel & s11) | (sub_sel & sub11) | (and_sel & and11) | (or_sel & or11);
  assign y12 = (add_sel & s12) | (sub_sel & sub12) | (and_sel & and12) | (or_sel & or12);
  assign y13 = (add_sel & s13) | (sub_sel & sub13) | (and_sel & and13) | (or_sel & or13);
  assign y14 = (add_sel & s14) | (sub_sel & sub14) | (and_sel & and14) | (or_sel & or14);
  assign y15 = (add_sel & s15) | (sub_sel & sub15) | (and_sel & and15) | (or_sel & or15);
  assign y16 = (add_sel & s16) | (sub_sel & sub16) | (and_sel & and16) | (or_sel & or16);
  assign y17 = (add_sel & s17) | (sub_sel & sub17) | (and_sel & and17) | (or_sel & or17);
  assign y18 = (add_sel & s18) | (sub_sel & sub18) | (and_sel & and18) | (or_sel & or18);
  assign y19 = (add_sel & s19) | (sub_sel & sub19) | (and_sel & and19) | (or_sel & or19);
  assign y20 = (add_sel & s20) | (sub_sel & sub20) | (and_sel & and20) | (or_sel & or20);
  assign y21 = (add_sel & s21) | (sub_sel & sub21) | (and_sel & and21) | (or_sel & or21);
  assign y22 = (add_sel & s22) | (sub_sel & sub22) | (and_sel & and22) | (or_sel & or22);
  assign y23 = (add_sel & s23) | (sub_sel & sub23) | (and_sel & and23) | (or_sel & or23);
  assign y24 = (add_sel & s24) | (sub_sel & sub24) | (and_sel & and24) | (or_sel & or24);
  assign y25 = (add_sel & s25) | (sub_sel & sub25) | (and_sel & and25) | (or_sel & or25);
  assign y26 = (add_sel & s26) | (sub_sel & sub26) | (and_sel & and26) | (or_sel & or26);
  assign y27 = (add_sel & s27) | (sub_sel & sub27) | (and_sel & and27) | (or_sel & or27);
  assign y28 = (add_sel & s28) | (sub_sel & sub28) | (and_sel & and28) | (or_sel & or28);
  assign y29 = (add_sel & s29) | (sub_sel & sub29) | (and_sel & and29) | (or_sel & or29);
  assign y30 = (add_sel & s30) | (sub_sel & sub30) | (and_sel & and30) | (or_sel & or30);
  assign y31 = (add_sel & s31) | (sub_sel & sub31) | (and_sel & and31) | (or_sel & or31);
  assign y32 = (add_sel & s32) | (sub_sel & sub32) | (and_sel & and32) | (or_sel & or32);
  assign y33 = (add_sel & s33) | (sub_sel & sub33) | (and_sel & and33) | (or_sel & or33);
  assign y34 = (add_sel & s34) | (sub_sel & sub34) | (and_sel & and34) | (or_sel & or34);
  assign y35 = (add_sel & s35) | (sub_sel & sub35) | (and_sel & and35) | (or_sel & or35);
  assign y36 = (add_sel & s36) | (sub_sel & sub36) | (and_sel & and36) | (or_sel & or36);
  assign y37 = (add_sel & s37) | (sub_sel & sub37) | (and_sel & and37) | (or_sel & or37);
  assign y38 = (add_sel & s38) | (sub_sel & sub38) | (and_sel & and38) | (or_sel & or38);
  assign y39 = (add_sel & s39) | (sub_sel & sub39) | (and_sel & and39) | (or_sel & or39);
  assign y40 = (add_sel & s40) | (sub_sel & sub40) | (and_sel & and40) | (or_sel & or40);
  assign y41 = (add_sel & s41) | (sub_sel & sub41) | (and_sel & and41) | (or_sel & or41);
  assign y42 = (add_sel & s42) | (sub_sel & sub42) | (and_sel & and42) | (or_sel & or42);
  assign y43 = (add_sel & s43) | (sub_sel & sub43) | (and_sel & and43) | (or_sel & or43);
  assign y44 = (add_sel & s44) | (sub_sel & sub44) | (and_sel & and44) | (or_sel & or44);
  assign y45 = (add_sel & s45) | (sub_sel & sub45) | (and_sel & and45) | (or_sel & or45);
  assign y46 = (add_sel & s46) | (sub_sel & sub46) | (and_sel & and46) | (or_sel & or46);
  assign y47 = (add_sel & s47) | (sub_sel & sub47) | (and_sel & and47) | (or_sel & or47);
  assign y48 = (add_sel & s48) | (sub_sel & sub48) | (and_sel & and48) | (or_sel & or48);
  assign y49 = (add_sel & s49) | (sub_sel & sub49) | (and_sel & and49) | (or_sel & or49);
  assign y50 = (add_sel & s50) | (sub_sel & sub50) | (and_sel & and50) | (or_sel & or50);
  assign y51 = (add_sel & s51) | (sub_sel & sub51) | (and_sel & and51) | (or_sel & or51);
  assign y52 = (add_sel & s52) | (sub_sel & sub52) | (and_sel & and52) | (or_sel & or52);
  assign y53 = (add_sel & s53) | (sub_sel & sub53) | (and_sel & and53) | (or_sel & or53);
  assign y54 = (add_sel & s54) | (sub_sel & sub54) | (and_sel & and54) | (or_sel & or54);
  assign y55 = (add_sel & s55) | (sub_sel & sub55) | (and_sel & and55) | (or_sel & or55);
  assign y56 = (add_sel & s56) | (sub_sel & sub56) | (and_sel & and56) | (or_sel & or56);
  assign y57 = (add_sel & s57) | (sub_sel & sub57) | (and_sel & and57) | (or_sel & or57);
  assign y58 = (add_sel & s58) | (sub_sel & sub58) | (and_sel & and58) | (or_sel & or58);
  assign y59 = (add_sel & s59) | (sub_sel & sub59) | (and_sel & and59) | (or_sel & or59);
  assign y60 = (add_sel & s60) | (sub_sel & sub60) | (and_sel & and60) | (or_sel & or60);
  assign y61 = (add_sel & s61) | (sub_sel & sub61) | (and_sel & and61) | (or_sel & or61);
  assign y62 = (add_sel & s62) | (sub_sel & sub62) | (and_sel & and62) | (or_sel & or62);
  assign y63 = (add_sel & s63) | (sub_sel & sub63) | (and_sel & and63) | (or_sel & or63);
  assign y64 = (add_sel & s64) | (sub_sel & sub64) | (and_sel & and64) | (or_sel & or64);
  assign y65 = (add_sel & s65) | (sub_sel & sub65) | (and_sel & and65) | (or_sel & or65);
  assign y66 = (add_sel & s66) | (sub_sel & sub66) | (and_sel & and66) | (or_sel & or66);
  assign y67 = (add_sel & s67) | (sub_sel & sub67) | (and_sel & and67) | (or_sel & or67);
  assign y68 = (add_sel & s68) | (sub_sel & sub68) | (and_sel & and68) | (or_sel & or68);
  assign y69 = (add_sel & s69) | (sub_sel & sub69) | (and_sel & and69) | (or_sel & or69);
  assign y70 = (add_sel & s70) | (sub_sel & sub70) | (and_sel & and70) | (or_sel & or70);
  assign y71 = (add_sel & s71) | (sub_sel & sub71) | (and_sel & and71) | (or_sel & or71);
  assign y72 = (add_sel & s72) | (sub_sel & sub72) | (and_sel & and72) | (or_sel & or72);
  assign y73 = (add_sel & s73) | (sub_sel & sub73) | (and_sel & and73) | (or_sel & or73);
  assign y74 = (add_sel & s74) | (sub_sel & sub74) | (and_sel & and74) | (or_sel & or74);
  assign y75 = (add_sel & s75) | (sub_sel & sub75) | (and_sel & and75) | (or_sel & or75);
  assign y76 = (add_sel & s76) | (sub_sel & sub76) | (and_sel & and76) | (or_sel & or76);
  assign y77 = (add_sel & s77) | (sub_sel & sub77) | (and_sel & and77) | (or_sel & or77);
  assign y78 = (add_sel & s78) | (sub_sel & sub78) | (and_sel & and78) | (or_sel & or78);
  assign y79 = (add_sel & s79) | (sub_sel & sub79) | (and_sel & and79) | (or_sel & or79);
  assign y80 = (add_sel & s80) | (sub_sel & sub80) | (and_sel & and80) | (or_sel & or80);
  assign y81 = (add_sel & s81) | (sub_sel & sub81) | (and_sel & and81) | (or_sel & or81);
  assign y82 = (add_sel & s82) | (sub_sel & sub82) | (and_sel & and82) | (or_sel & or82);
  assign y83 = (add_sel & s83) | (sub_sel & sub83) | (and_sel & and83) | (or_sel & or83);
  assign y84 = (add_sel & s84) | (sub_sel & sub84) | (and_sel & and84) | (or_sel & or84);
  assign y85 = (add_sel & s85) | (sub_sel & sub85) | (and_sel & and85) | (or_sel & or85);
  assign y86 = (add_sel & s86) | (sub_sel & sub86) | (and_sel & and86) | (or_sel & or86);
  assign y87 = (add_sel & s87) | (sub_sel & sub87) | (and_sel & and87) | (or_sel & or87);
  assign y88 = (add_sel & s88) | (sub_sel & sub88) | (and_sel & and88) | (or_sel & or88);
  assign y89 = (add_sel & s89) | (sub_sel & sub89) | (and_sel & and89) | (or_sel & or89);
  assign y90 = (add_sel & s90) | (sub_sel & sub90) | (and_sel & and90) | (or_sel & or90);
  assign y91 = (add_sel & s91) | (sub_sel & sub91) | (and_sel & and91) | (or_sel & or91);
  assign y92 = (add_sel & s92) | (sub_sel & sub92) | (and_sel & and92) | (or_sel & or92);
  assign y93 = (add_sel & s93) | (sub_sel & sub93) | (and_sel & and93) | (or_sel & or93);
  assign y94 = (add_sel & s94) | (sub_sel & sub94) | (and_sel & and94) | (or_sel & or94);
  assign y95 = (add_sel & s95) | (sub_sel & sub95) | (and_sel & and95) | (or_sel & or95);
  assign y96 = (add_sel & s96) | (sub_sel & sub96) | (and_sel & and96) | (or_sel & or96);
  assign y97 = (add_sel & s97) | (sub_sel & sub97) | (and_sel & and97) | (or_sel & or97);
  assign y98 = (add_sel & s98) | (sub_sel & sub98) | (and_sel & and98) | (or_sel & or98);
  assign y99 = (add_sel & s99) | (sub_sel & sub99) | (and_sel & and99) | (or_sel & or99);
  assign y100 = (add_sel & s100) | (sub_sel & sub100) | (and_sel & and100) | (or_sel & or100);
  assign y101 = (add_sel & s101) | (sub_sel & sub101) | (and_sel & and101) | (or_sel & or101);
  assign y102 = (add_sel & s102) | (sub_sel & sub102) | (and_sel & and102) | (or_sel & or102);
  assign y103 = (add_sel & s103) | (sub_sel & sub103) | (and_sel & and103) | (or_sel & or103);
  assign y104 = (add_sel & s104) | (sub_sel & sub104) | (and_sel & and104) | (or_sel & or104);
  assign y105 = (add_sel & s105) | (sub_sel & sub105) | (and_sel & and105) | (or_sel & or105);
  assign y106 = (add_sel & s106) | (sub_sel & sub106) | (and_sel & and106) | (or_sel & or106);
  assign y107 = (add_sel & s107) | (sub_sel & sub107) | (and_sel & and107) | (or_sel & or107);
  assign y108 = (add_sel & s108) | (sub_sel & sub108) | (and_sel & and108) | (or_sel & or108);
  assign y109 = (add_sel & s109) | (sub_sel & sub109) | (and_sel & and109) | (or_sel & or109);
  assign y110 = (add_sel & s110) | (sub_sel & sub110) | (and_sel & and110) | (or_sel & or110);
  assign y111 = (add_sel & s111) | (sub_sel & sub111) | (and_sel & and111) | (or_sel & or111);
  assign y112 = (add_sel & s112) | (sub_sel & sub112) | (and_sel & and112) | (or_sel & or112);
  assign y113 = (add_sel & s113) | (sub_sel & sub113) | (and_sel & and113) | (or_sel & or113);
  assign y114 = (add_sel & s114) | (sub_sel & sub114) | (and_sel & and114) | (or_sel & or114);
  assign y115 = (add_sel & s115) | (sub_sel & sub115) | (and_sel & and115) | (or_sel & or115);
  assign y116 = (add_sel & s116) | (sub_sel & sub116) | (and_sel & and116) | (or_sel & or116);
  assign y117 = (add_sel & s117) | (sub_sel & sub117) | (and_sel & and117) | (or_sel & or117);
  assign y118 = (add_sel & s118) | (sub_sel & sub118) | (and_sel & and118) | (or_sel & or118);
  assign y119 = (add_sel & s119) | (sub_sel & sub119) | (and_sel & and119) | (or_sel & or119);
  assign y120 = (add_sel & s120) | (sub_sel & sub120) | (and_sel & and120) | (or_sel & or120);
  assign y121 = (add_sel & s121) | (sub_sel & sub121) | (and_sel & and121) | (or_sel & or121);
  assign y122 = (add_sel & s122) | (sub_sel & sub122) | (and_sel & and122) | (or_sel & or122);
  assign y123 = (add_sel & s123) | (sub_sel & sub123) | (and_sel & and123) | (or_sel & or123);
  assign y124 = (add_sel & s124) | (sub_sel & sub124) | (and_sel & and124) | (or_sel & or124);
  assign y125 = (add_sel & s125) | (sub_sel & sub125) | (and_sel & and125) | (or_sel & or125);
  assign y126 = (add_sel & s126) | (sub_sel & sub126) | (and_sel & and126) | (or_sel & or126);
  assign y127 = (add_sel & s127) | (sub_sel & sub127) | (and_sel & and127) | (or_sel & or127);
  assign y128 = (add_sel & s128) | (sub_sel & sub128) | (and_sel & and128) | (or_sel & or128);
  assign y129 = (add_sel & s129) | (sub_sel & sub129) | (and_sel & and129) | (or_sel & or129);
  assign y130 = (add_sel & s130) | (sub_sel & sub130) | (and_sel & and130) | (or_sel & or130);
  assign y131 = (add_sel & s131) | (sub_sel & sub131) | (and_sel & and131) | (or_sel & or131);
  assign y132 = (add_sel & s132) | (sub_sel & sub132) | (and_sel & and132) | (or_sel & or132);
  assign y133 = (add_sel & s133) | (sub_sel & sub133) | (and_sel & and133) | (or_sel & or133);
  assign y134 = (add_sel & s134) | (sub_sel & sub134) | (and_sel & and134) | (or_sel & or134);
  assign y135 = (add_sel & s135) | (sub_sel & sub135) | (and_sel & and135) | (or_sel & or135);
  assign y136 = (add_sel & s136) | (sub_sel & sub136) | (and_sel & and136) | (or_sel & or136);
  assign y137 = (add_sel & s137) | (sub_sel & sub137) | (and_sel & and137) | (or_sel & or137);
  assign y138 = (add_sel & s138) | (sub_sel & sub138) | (and_sel & and138) | (or_sel & or138);
  assign y139 = (add_sel & s139) | (sub_sel & sub139) | (and_sel & and139) | (or_sel & or139);
  assign y140 = (add_sel & s140) | (sub_sel & sub140) | (and_sel & and140) | (or_sel & or140);
  assign y141 = (add_sel & s141) | (sub_sel & sub141) | (and_sel & and141) | (or_sel & or141);
  assign y142 = (add_sel & s142) | (sub_sel & sub142) | (and_sel & and142) | (or_sel & or142);
  assign y143 = (add_sel & s143) | (sub_sel & sub143) | (and_sel & and143) | (or_sel & or143);
  assign y144 = (add_sel & s144) | (sub_sel & sub144) | (and_sel & and144) | (or_sel & or144);
  assign y145 = (add_sel & s145) | (sub_sel & sub145) | (and_sel & and145) | (or_sel & or145);
  assign y146 = (add_sel & s146) | (sub_sel & sub146) | (and_sel & and146) | (or_sel & or146);
  assign y147 = (add_sel & s147) | (sub_sel & sub147) | (and_sel & and147) | (or_sel & or147);
  assign y148 = (add_sel & s148) | (sub_sel & sub148) | (and_sel & and148) | (or_sel & or148);
  assign y149 = (add_sel & s149) | (sub_sel & sub149) | (and_sel & and149) | (or_sel & or149);
  assign y150 = (add_sel & s150) | (sub_sel & sub150) | (and_sel & and150) | (or_sel & or150);
  assign y151 = (add_sel & s151) | (sub_sel & sub151) | (and_sel & and151) | (or_sel & or151);
  assign y152 = (add_sel & s152) | (sub_sel & sub152) | (and_sel & and152) | (or_sel & or152);
  assign y153 = (add_sel & s153) | (sub_sel & sub153) | (and_sel & and153) | (or_sel & or153);
  assign y154 = (add_sel & s154) | (sub_sel & sub154) | (and_sel & and154) | (or_sel & or154);
  assign y155 = (add_sel & s155) | (sub_sel & sub155) | (and_sel & and155) | (or_sel & or155);
  assign y156 = (add_sel & s156) | (sub_sel & sub156) | (and_sel & and156) | (or_sel & or156);
  assign y157 = (add_sel & s157) | (sub_sel & sub157) | (and_sel & and157) | (or_sel & or157);
  assign y158 = (add_sel & s158) | (sub_sel & sub158) | (and_sel & and158) | (or_sel & or158);
  assign y159 = (add_sel & s159) | (sub_sel & sub159) | (and_sel & and159) | (or_sel & or159);
  assign y160 = (add_sel & s160) | (sub_sel & sub160) | (and_sel & and160) | (or_sel & or160);
  assign y161 = (add_sel & s161) | (sub_sel & sub161) | (and_sel & and161) | (or_sel & or161);
  assign y162 = (add_sel & s162) | (sub_sel & sub162) | (and_sel & and162) | (or_sel & or162);
  assign y163 = (add_sel & s163) | (sub_sel & sub163) | (and_sel & and163) | (or_sel & or163);
  assign y164 = (add_sel & s164) | (sub_sel & sub164) | (and_sel & and164) | (or_sel & or164);
  assign y165 = (add_sel & s165) | (sub_sel & sub165) | (and_sel & and165) | (or_sel & or165);
  assign y166 = (add_sel & s166) | (sub_sel & sub166) | (and_sel & and166) | (or_sel & or166);
  assign y167 = (add_sel & s167) | (sub_sel & sub167) | (and_sel & and167) | (or_sel & or167);
  assign y168 = (add_sel & s168) | (sub_sel & sub168) | (and_sel & and168) | (or_sel & or168);
  assign y169 = (add_sel & s169) | (sub_sel & sub169) | (and_sel & and169) | (or_sel & or169);
  assign y170 = (add_sel & s170) | (sub_sel & sub170) | (and_sel & and170) | (or_sel & or170);
  assign y171 = (add_sel & s171) | (sub_sel & sub171) | (and_sel & and171) | (or_sel & or171);
  assign y172 = (add_sel & s172) | (sub_sel & sub172) | (and_sel & and172) | (or_sel & or172);
  assign y173 = (add_sel & s173) | (sub_sel & sub173) | (and_sel & and173) | (or_sel & or173);
  assign y174 = (add_sel & s174) | (sub_sel & sub174) | (and_sel & and174) | (or_sel & or174);
  assign y175 = (add_sel & s175) | (sub_sel & sub175) | (and_sel & and175) | (or_sel & or175);
  assign y176 = (add_sel & s176) | (sub_sel & sub176) | (and_sel & and176) | (or_sel & or176);
  assign y177 = (add_sel & s177) | (sub_sel & sub177) | (and_sel & and177) | (or_sel & or177);
  assign y178 = (add_sel & s178) | (sub_sel & sub178) | (and_sel & and178) | (or_sel & or178);
  assign y179 = (add_sel & s179) | (sub_sel & sub179) | (and_sel & and179) | (or_sel & or179);
  assign y180 = (add_sel & s180) | (sub_sel & sub180) | (and_sel & and180) | (or_sel & or180);
  assign y181 = (add_sel & s181) | (sub_sel & sub181) | (and_sel & and181) | (or_sel & or181);
  assign y182 = (add_sel & s182) | (sub_sel & sub182) | (and_sel & and182) | (or_sel & or182);
  assign y183 = (add_sel & s183) | (sub_sel & sub183) | (and_sel & and183) | (or_sel & or183);
  assign y184 = (add_sel & s184) | (sub_sel & sub184) | (and_sel & and184) | (or_sel & or184);
  assign y185 = (add_sel & s185) | (sub_sel & sub185) | (and_sel & and185) | (or_sel & or185);
  assign y186 = (add_sel & s186) | (sub_sel & sub186) | (and_sel & and186) | (or_sel & or186);
  assign y187 = (add_sel & s187) | (sub_sel & sub187) | (and_sel & and187) | (or_sel & or187);
  assign y188 = (add_sel & s188) | (sub_sel & sub188) | (and_sel & and188) | (or_sel & or188);
  assign y189 = (add_sel & s189) | (sub_sel & sub189) | (and_sel & and189) | (or_sel & or189);
  assign y190 = (add_sel & s190) | (sub_sel & sub190) | (and_sel & and190) | (or_sel & or190);
  assign y191 = (add_sel & s191) | (sub_sel & sub191) | (and_sel & and191) | (or_sel & or191);
  assign y192 = (add_sel & s192) | (sub_sel & sub192) | (and_sel & and192) | (or_sel & or192);
  assign y193 = (add_sel & s193) | (sub_sel & sub193) | (and_sel & and193) | (or_sel & or193);
  assign y194 = (add_sel & s194) | (sub_sel & sub194) | (and_sel & and194) | (or_sel & or194);
  assign y195 = (add_sel & s195) | (sub_sel & sub195) | (and_sel & and195) | (or_sel & or195);
  assign y196 = (add_sel & s196) | (sub_sel & sub196) | (and_sel & and196) | (or_sel & or196);
  assign y197 = (add_sel & s197) | (sub_sel & sub197) | (and_sel & and197) | (or_sel & or197);
  assign y198 = (add_sel & s198) | (sub_sel & sub198) | (and_sel & and198) | (or_sel & or198);
  assign y199 = (add_sel & s199) | (sub_sel & sub199) | (and_sel & and199) | (or_sel & or199);
  assign y200 = (add_sel & s200) | (sub_sel & sub200) | (and_sel & and200) | (or_sel & or200);
  assign y201 = (add_sel & s201) | (sub_sel & sub201) | (and_sel & and201) | (or_sel & or201);
  assign y202 = (add_sel & s202) | (sub_sel & sub202) | (and_sel & and202) | (or_sel & or202);
  assign y203 = (add_sel & s203) | (sub_sel & sub203) | (and_sel & and203) | (or_sel & or203);
  assign y204 = (add_sel & s204) | (sub_sel & sub204) | (and_sel & and204) | (or_sel & or204);
  assign y205 = (add_sel & s205) | (sub_sel & sub205) | (and_sel & and205) | (or_sel & or205);
  assign y206 = (add_sel & s206) | (sub_sel & sub206) | (and_sel & and206) | (or_sel & or206);
  assign y207 = (add_sel & s207) | (sub_sel & sub207) | (and_sel & and207) | (or_sel & or207);
  assign y208 = (add_sel & s208) | (sub_sel & sub208) | (and_sel & and208) | (or_sel & or208);
  assign y209 = (add_sel & s209) | (sub_sel & sub209) | (and_sel & and209) | (or_sel & or209);
  assign y210 = (add_sel & s210) | (sub_sel & sub210) | (and_sel & and210) | (or_sel & or210);
  assign y211 = (add_sel & s211) | (sub_sel & sub211) | (and_sel & and211) | (or_sel & or211);
  assign y212 = (add_sel & s212) | (sub_sel & sub212) | (and_sel & and212) | (or_sel & or212);
  assign y213 = (add_sel & s213) | (sub_sel & sub213) | (and_sel & and213) | (or_sel & or213);
  assign y214 = (add_sel & s214) | (sub_sel & sub214) | (and_sel & and214) | (or_sel & or214);
  assign y215 = (add_sel & s215) | (sub_sel & sub215) | (and_sel & and215) | (or_sel & or215);
  assign y216 = (add_sel & s216) | (sub_sel & sub216) | (and_sel & and216) | (or_sel & or216);
  assign y217 = (add_sel & s217) | (sub_sel & sub217) | (and_sel & and217) | (or_sel & or217);
  assign y218 = (add_sel & s218) | (sub_sel & sub218) | (and_sel & and218) | (or_sel & or218);
  assign y219 = (add_sel & s219) | (sub_sel & sub219) | (and_sel & and219) | (or_sel & or219);
  assign y220 = (add_sel & s220) | (sub_sel & sub220) | (and_sel & and220) | (or_sel & or220);
  assign y221 = (add_sel & s221) | (sub_sel & sub221) | (and_sel & and221) | (or_sel & or221);
  assign y222 = (add_sel & s222) | (sub_sel & sub222) | (and_sel & and222) | (or_sel & or222);
  assign y223 = (add_sel & s223) | (sub_sel & sub223) | (and_sel & and223) | (or_sel & or223);
  assign y224 = (add_sel & s224) | (sub_sel & sub224) | (and_sel & and224) | (or_sel & or224);
  assign y225 = (add_sel & s225) | (sub_sel & sub225) | (and_sel & and225) | (or_sel & or225);
  assign y226 = (add_sel & s226) | (sub_sel & sub226) | (and_sel & and226) | (or_sel & or226);
  assign y227 = (add_sel & s227) | (sub_sel & sub227) | (and_sel & and227) | (or_sel & or227);
  assign y228 = (add_sel & s228) | (sub_sel & sub228) | (and_sel & and228) | (or_sel & or228);
  assign y229 = (add_sel & s229) | (sub_sel & sub229) | (and_sel & and229) | (or_sel & or229);
  assign y230 = (add_sel & s230) | (sub_sel & sub230) | (and_sel & and230) | (or_sel & or230);
  assign y231 = (add_sel & s231) | (sub_sel & sub231) | (and_sel & and231) | (or_sel & or231);
  assign y232 = (add_sel & s232) | (sub_sel & sub232) | (and_sel & and232) | (or_sel & or232);
  assign y233 = (add_sel & s233) | (sub_sel & sub233) | (and_sel & and233) | (or_sel & or233);
  assign y234 = (add_sel & s234) | (sub_sel & sub234) | (and_sel & and234) | (or_sel & or234);
  assign y235 = (add_sel & s235) | (sub_sel & sub235) | (and_sel & and235) | (or_sel & or235);
  assign y236 = (add_sel & s236) | (sub_sel & sub236) | (and_sel & and236) | (or_sel & or236);
  assign y237 = (add_sel & s237) | (sub_sel & sub237) | (and_sel & and237) | (or_sel & or237);
  assign y238 = (add_sel & s238) | (sub_sel & sub238) | (and_sel & and238) | (or_sel & or238);
  assign y239 = (add_sel & s239) | (sub_sel & sub239) | (and_sel & and239) | (or_sel & or239);
  assign y240 = (add_sel & s240) | (sub_sel & sub240) | (and_sel & and240) | (or_sel & or240);
  assign y241 = (add_sel & s241) | (sub_sel & sub241) | (and_sel & and241) | (or_sel & or241);
  assign y242 = (add_sel & s242) | (sub_sel & sub242) | (and_sel & and242) | (or_sel & or242);
  assign y243 = (add_sel & s243) | (sub_sel & sub243) | (and_sel & and243) | (or_sel & or243);
  assign y244 = (add_sel & s244) | (sub_sel & sub244) | (and_sel & and244) | (or_sel & or244);
  assign y245 = (add_sel & s245) | (sub_sel & sub245) | (and_sel & and245) | (or_sel & or245);
  assign y246 = (add_sel & s246) | (sub_sel & sub246) | (and_sel & and246) | (or_sel & or246);
  assign y247 = (add_sel & s247) | (sub_sel & sub247) | (and_sel & and247) | (or_sel & or247);
  assign y248 = (add_sel & s248) | (sub_sel & sub248) | (and_sel & and248) | (or_sel & or248);
  assign y249 = (add_sel & s249) | (sub_sel & sub249) | (and_sel & and249) | (or_sel & or249);
  assign y250 = (add_sel & s250) | (sub_sel & sub250) | (and_sel & and250) | (or_sel & or250);
  assign y251 = (add_sel & s251) | (sub_sel & sub251) | (and_sel & and251) | (or_sel & or251);
  assign y252 = (add_sel & s252) | (sub_sel & sub252) | (and_sel & and252) | (or_sel & or252);
  assign y253 = (add_sel & s253) | (sub_sel & sub253) | (and_sel & and253) | (or_sel & or253);
  assign y254 = (add_sel & s254) | (sub_sel & sub254) | (and_sel & and254) | (or_sel & or254);
  assign y255 = (add_sel & s255) | (sub_sel & sub255) | (and_sel & and255) | (or_sel & or255);
  assign y256 = (add_sel & s256) | (sub_sel & sub256) | (and_sel & and256) | (or_sel & or256);
  assign y257 = (add_sel & s257) | (sub_sel & sub257) | (and_sel & and257) | (or_sel & or257);
  assign y258 = (add_sel & s258) | (sub_sel & sub258) | (and_sel & and258) | (or_sel & or258);
  assign y259 = (add_sel & s259) | (sub_sel & sub259) | (and_sel & and259) | (or_sel & or259);
  assign y260 = (add_sel & s260) | (sub_sel & sub260) | (and_sel & and260) | (or_sel & or260);
  assign y261 = (add_sel & s261) | (sub_sel & sub261) | (and_sel & and261) | (or_sel & or261);
  assign y262 = (add_sel & s262) | (sub_sel & sub262) | (and_sel & and262) | (or_sel & or262);
  assign y263 = (add_sel & s263) | (sub_sel & sub263) | (and_sel & and263) | (or_sel & or263);
  assign y264 = (add_sel & s264) | (sub_sel & sub264) | (and_sel & and264) | (or_sel & or264);
  assign y265 = (add_sel & s265) | (sub_sel & sub265) | (and_sel & and265) | (or_sel & or265);
  assign y266 = (add_sel & s266) | (sub_sel & sub266) | (and_sel & and266) | (or_sel & or266);
  assign y267 = (add_sel & s267) | (sub_sel & sub267) | (and_sel & and267) | (or_sel & or267);
  assign y268 = (add_sel & s268) | (sub_sel & sub268) | (and_sel & and268) | (or_sel & or268);
  assign y269 = (add_sel & s269) | (sub_sel & sub269) | (and_sel & and269) | (or_sel & or269);
  assign y270 = (add_sel & s270) | (sub_sel & sub270) | (and_sel & and270) | (or_sel & or270);
  assign y271 = (add_sel & s271) | (sub_sel & sub271) | (and_sel & and271) | (or_sel & or271);
  assign y272 = (add_sel & s272) | (sub_sel & sub272) | (and_sel & and272) | (or_sel & or272);
  assign y273 = (add_sel & s273) | (sub_sel & sub273) | (and_sel & and273) | (or_sel & or273);
  assign y274 = (add_sel & s274) | (sub_sel & sub274) | (and_sel & and274) | (or_sel & or274);
  assign y275 = (add_sel & s275) | (sub_sel & sub275) | (and_sel & and275) | (or_sel & or275);
  assign y276 = (add_sel & s276) | (sub_sel & sub276) | (and_sel & and276) | (or_sel & or276);
  assign y277 = (add_sel & s277) | (sub_sel & sub277) | (and_sel & and277) | (or_sel & or277);
  assign y278 = (add_sel & s278) | (sub_sel & sub278) | (and_sel & and278) | (or_sel & or278);
  assign y279 = (add_sel & s279) | (sub_sel & sub279) | (and_sel & and279) | (or_sel & or279);
  assign y280 = (add_sel & s280) | (sub_sel & sub280) | (and_sel & and280) | (or_sel & or280);
  assign y281 = (add_sel & s281) | (sub_sel & sub281) | (and_sel & and281) | (or_sel & or281);
  assign y282 = (add_sel & s282) | (sub_sel & sub282) | (and_sel & and282) | (or_sel & or282);
  assign y283 = (add_sel & s283) | (sub_sel & sub283) | (and_sel & and283) | (or_sel & or283);
  assign y284 = (add_sel & s284) | (sub_sel & sub284) | (and_sel & and284) | (or_sel & or284);
  assign y285 = (add_sel & s285) | (sub_sel & sub285) | (and_sel & and285) | (or_sel & or285);
  assign y286 = (add_sel & s286) | (sub_sel & sub286) | (and_sel & and286) | (or_sel & or286);
  assign y287 = (add_sel & s287) | (sub_sel & sub287) | (and_sel & and287) | (or_sel & or287);
  assign y288 = (add_sel & s288) | (sub_sel & sub288) | (and_sel & and288) | (or_sel & or288);
  assign y289 = (add_sel & s289) | (sub_sel & sub289) | (and_sel & and289) | (or_sel & or289);
  assign y290 = (add_sel & s290) | (sub_sel & sub290) | (and_sel & and290) | (or_sel & or290);
  assign y291 = (add_sel & s291) | (sub_sel & sub291) | (and_sel & and291) | (or_sel & or291);
  assign y292 = (add_sel & s292) | (sub_sel & sub292) | (and_sel & and292) | (or_sel & or292);
  assign y293 = (add_sel & s293) | (sub_sel & sub293) | (and_sel & and293) | (or_sel & or293);
  assign y294 = (add_sel & s294) | (sub_sel & sub294) | (and_sel & and294) | (or_sel & or294);
  assign y295 = (add_sel & s295) | (sub_sel & sub295) | (and_sel & and295) | (or_sel & or295);
  assign y296 = (add_sel & s296) | (sub_sel & sub296) | (and_sel & and296) | (or_sel & or296);
  assign y297 = (add_sel & s297) | (sub_sel & sub297) | (and_sel & and297) | (or_sel & or297);
  assign y298 = (add_sel & s298) | (sub_sel & sub298) | (and_sel & and298) | (or_sel & or298);
  assign y299 = (add_sel & s299) | (sub_sel & sub299) | (and_sel & and299) | (or_sel & or299);
  assign y300 = (add_sel & s300) | (sub_sel & sub300) | (and_sel & and300) | (or_sel & or300);
  assign y301 = (add_sel & s301) | (sub_sel & sub301) | (and_sel & and301) | (or_sel & or301);
  assign y302 = (add_sel & s302) | (sub_sel & sub302) | (and_sel & and302) | (or_sel & or302);
  assign y303 = (add_sel & s303) | (sub_sel & sub303) | (and_sel & and303) | (or_sel & or303);
  assign y304 = (add_sel & s304) | (sub_sel & sub304) | (and_sel & and304) | (or_sel & or304);
  assign y305 = (add_sel & s305) | (sub_sel & sub305) | (and_sel & and305) | (or_sel & or305);
  assign y306 = (add_sel & s306) | (sub_sel & sub306) | (and_sel & and306) | (or_sel & or306);
  assign y307 = (add_sel & s307) | (sub_sel & sub307) | (and_sel & and307) | (or_sel & or307);
  assign y308 = (add_sel & s308) | (sub_sel & sub308) | (and_sel & and308) | (or_sel & or308);
  assign y309 = (add_sel & s309) | (sub_sel & sub309) | (and_sel & and309) | (or_sel & or309);
  assign y310 = (add_sel & s310) | (sub_sel & sub310) | (and_sel & and310) | (or_sel & or310);
  assign y311 = (add_sel & s311) | (sub_sel & sub311) | (and_sel & and311) | (or_sel & or311);
  assign y312 = (add_sel & s312) | (sub_sel & sub312) | (and_sel & and312) | (or_sel & or312);
  assign y313 = (add_sel & s313) | (sub_sel & sub313) | (and_sel & and313) | (or_sel & or313);
  assign y314 = (add_sel & s314) | (sub_sel & sub314) | (and_sel & and314) | (or_sel & or314);
  assign y315 = (add_sel & s315) | (sub_sel & sub315) | (and_sel & and315) | (or_sel & or315);
  assign y316 = (add_sel & s316) | (sub_sel & sub316) | (and_sel & and316) | (or_sel & or316);
  assign y317 = (add_sel & s317) | (sub_sel & sub317) | (and_sel & and317) | (or_sel & or317);
  assign y318 = (add_sel & s318) | (sub_sel & sub318) | (and_sel & and318) | (or_sel & or318);
  assign y319 = (add_sel & s319) | (sub_sel & sub319) | (and_sel & and319) | (or_sel & or319);
  assign y320 = (add_sel & s320) | (sub_sel & sub320) | (and_sel & and320) | (or_sel & or320);
  assign y321 = (add_sel & s321) | (sub_sel & sub321) | (and_sel & and321) | (or_sel & or321);
  assign y322 = (add_sel & s322) | (sub_sel & sub322) | (and_sel & and322) | (or_sel & or322);
  assign y323 = (add_sel & s323) | (sub_sel & sub323) | (and_sel & and323) | (or_sel & or323);
  assign y324 = (add_sel & s324) | (sub_sel & sub324) | (and_sel & and324) | (or_sel & or324);
  assign y325 = (add_sel & s325) | (sub_sel & sub325) | (and_sel & and325) | (or_sel & or325);
  assign y326 = (add_sel & s326) | (sub_sel & sub326) | (and_sel & and326) | (or_sel & or326);
  assign y327 = (add_sel & s327) | (sub_sel & sub327) | (and_sel & and327) | (or_sel & or327);
  assign y328 = (add_sel & s328) | (sub_sel & sub328) | (and_sel & and328) | (or_sel & or328);
  assign y329 = (add_sel & s329) | (sub_sel & sub329) | (and_sel & and329) | (or_sel & or329);
  assign y330 = (add_sel & s330) | (sub_sel & sub330) | (and_sel & and330) | (or_sel & or330);
  assign y331 = (add_sel & s331) | (sub_sel & sub331) | (and_sel & and331) | (or_sel & or331);
  assign y332 = (add_sel & s332) | (sub_sel & sub332) | (and_sel & and332) | (or_sel & or332);
  assign y333 = (add_sel & s333) | (sub_sel & sub333) | (and_sel & and333) | (or_sel & or333);
  assign y334 = (add_sel & s334) | (sub_sel & sub334) | (and_sel & and334) | (or_sel & or334);
  assign y335 = (add_sel & s335) | (sub_sel & sub335) | (and_sel & and335) | (or_sel & or335);
  assign y336 = (add_sel & s336) | (sub_sel & sub336) | (and_sel & and336) | (or_sel & or336);
  assign y337 = (add_sel & s337) | (sub_sel & sub337) | (and_sel & and337) | (or_sel & or337);
  assign y338 = (add_sel & s338) | (sub_sel & sub338) | (and_sel & and338) | (or_sel & or338);
  assign y339 = (add_sel & s339) | (sub_sel & sub339) | (and_sel & and339) | (or_sel & or339);
  assign y340 = (add_sel & s340) | (sub_sel & sub340) | (and_sel & and340) | (or_sel & or340);
  assign y341 = (add_sel & s341) | (sub_sel & sub341) | (and_sel & and341) | (or_sel & or341);
  assign y342 = (add_sel & s342) | (sub_sel & sub342) | (and_sel & and342) | (or_sel & or342);
  assign y343 = (add_sel & s343) | (sub_sel & sub343) | (and_sel & and343) | (or_sel & or343);
  assign y344 = (add_sel & s344) | (sub_sel & sub344) | (and_sel & and344) | (or_sel & or344);
  assign y345 = (add_sel & s345) | (sub_sel & sub345) | (and_sel & and345) | (or_sel & or345);
  assign y346 = (add_sel & s346) | (sub_sel & sub346) | (and_sel & and346) | (or_sel & or346);
  assign y347 = (add_sel & s347) | (sub_sel & sub347) | (and_sel & and347) | (or_sel & or347);
  assign y348 = (add_sel & s348) | (sub_sel & sub348) | (and_sel & and348) | (or_sel & or348);
  assign y349 = (add_sel & s349) | (sub_sel & sub349) | (and_sel & and349) | (or_sel & or349);
  assign y350 = (add_sel & s350) | (sub_sel & sub350) | (and_sel & and350) | (or_sel & or350);
  assign y351 = (add_sel & s351) | (sub_sel & sub351) | (and_sel & and351) | (or_sel & or351);
  assign y352 = (add_sel & s352) | (sub_sel & sub352) | (and_sel & and352) | (or_sel & or352);
  assign y353 = (add_sel & s353) | (sub_sel & sub353) | (and_sel & and353) | (or_sel & or353);
  assign y354 = (add_sel & s354) | (sub_sel & sub354) | (and_sel & and354) | (or_sel & or354);
  assign y355 = (add_sel & s355) | (sub_sel & sub355) | (and_sel & and355) | (or_sel & or355);
  assign y356 = (add_sel & s356) | (sub_sel & sub356) | (and_sel & and356) | (or_sel & or356);
  assign y357 = (add_sel & s357) | (sub_sel & sub357) | (and_sel & and357) | (or_sel & or357);
  assign y358 = (add_sel & s358) | (sub_sel & sub358) | (and_sel & and358) | (or_sel & or358);
  assign y359 = (add_sel & s359) | (sub_sel & sub359) | (and_sel & and359) | (or_sel & or359);
  assign y360 = (add_sel & s360) | (sub_sel & sub360) | (and_sel & and360) | (or_sel & or360);
  assign y361 = (add_sel & s361) | (sub_sel & sub361) | (and_sel & and361) | (or_sel & or361);
  assign y362 = (add_sel & s362) | (sub_sel & sub362) | (and_sel & and362) | (or_sel & or362);
  assign y363 = (add_sel & s363) | (sub_sel & sub363) | (and_sel & and363) | (or_sel & or363);
  assign y364 = (add_sel & s364) | (sub_sel & sub364) | (and_sel & and364) | (or_sel & or364);
  assign y365 = (add_sel & s365) | (sub_sel & sub365) | (and_sel & and365) | (or_sel & or365);
  assign y366 = (add_sel & s366) | (sub_sel & sub366) | (and_sel & and366) | (or_sel & or366);
  assign y367 = (add_sel & s367) | (sub_sel & sub367) | (and_sel & and367) | (or_sel & or367);
  assign y368 = (add_sel & s368) | (sub_sel & sub368) | (and_sel & and368) | (or_sel & or368);
  assign y369 = (add_sel & s369) | (sub_sel & sub369) | (and_sel & and369) | (or_sel & or369);
  assign y370 = (add_sel & s370) | (sub_sel & sub370) | (and_sel & and370) | (or_sel & or370);
  assign y371 = (add_sel & s371) | (sub_sel & sub371) | (and_sel & and371) | (or_sel & or371);
  assign y372 = (add_sel & s372) | (sub_sel & sub372) | (and_sel & and372) | (or_sel & or372);
  assign y373 = (add_sel & s373) | (sub_sel & sub373) | (and_sel & and373) | (or_sel & or373);
  assign y374 = (add_sel & s374) | (sub_sel & sub374) | (and_sel & and374) | (or_sel & or374);
  assign y375 = (add_sel & s375) | (sub_sel & sub375) | (and_sel & and375) | (or_sel & or375);
  assign y376 = (add_sel & s376) | (sub_sel & sub376) | (and_sel & and376) | (or_sel & or376);
  assign y377 = (add_sel & s377) | (sub_sel & sub377) | (and_sel & and377) | (or_sel & or377);
  assign y378 = (add_sel & s378) | (sub_sel & sub378) | (and_sel & and378) | (or_sel & or378);
  assign y379 = (add_sel & s379) | (sub_sel & sub379) | (and_sel & and379) | (or_sel & or379);
  assign y380 = (add_sel & s380) | (sub_sel & sub380) | (and_sel & and380) | (or_sel & or380);
  assign y381 = (add_sel & s381) | (sub_sel & sub381) | (and_sel & and381) | (or_sel & or381);
  assign y382 = (add_sel & s382) | (sub_sel & sub382) | (and_sel & and382) | (or_sel & or382);
  assign y383 = (add_sel & s383) | (sub_sel & sub383) | (and_sel & and383) | (or_sel & or383);
  assign y384 = (add_sel & s384) | (sub_sel & sub384) | (and_sel & and384) | (or_sel & or384);
  assign y385 = (add_sel & s385) | (sub_sel & sub385) | (and_sel & and385) | (or_sel & or385);
  assign y386 = (add_sel & s386) | (sub_sel & sub386) | (and_sel & and386) | (or_sel & or386);
  assign y387 = (add_sel & s387) | (sub_sel & sub387) | (and_sel & and387) | (or_sel & or387);
  assign y388 = (add_sel & s388) | (sub_sel & sub388) | (and_sel & and388) | (or_sel & or388);
  assign y389 = (add_sel & s389) | (sub_sel & sub389) | (and_sel & and389) | (or_sel & or389);
  assign y390 = (add_sel & s390) | (sub_sel & sub390) | (and_sel & and390) | (or_sel & or390);
  assign y391 = (add_sel & s391) | (sub_sel & sub391) | (and_sel & and391) | (or_sel & or391);
  assign y392 = (add_sel & s392) | (sub_sel & sub392) | (and_sel & and392) | (or_sel & or392);
  assign y393 = (add_sel & s393) | (sub_sel & sub393) | (and_sel & and393) | (or_sel & or393);
  assign y394 = (add_sel & s394) | (sub_sel & sub394) | (and_sel & and394) | (or_sel & or394);
  assign y395 = (add_sel & s395) | (sub_sel & sub395) | (and_sel & and395) | (or_sel & or395);
  assign y396 = (add_sel & s396) | (sub_sel & sub396) | (and_sel & and396) | (or_sel & or396);
  assign y397 = (add_sel & s397) | (sub_sel & sub397) | (and_sel & and397) | (or_sel & or397);
  assign y398 = (add_sel & s398) | (sub_sel & sub398) | (and_sel & and398) | (or_sel & or398);
  assign y399 = (add_sel & s399) | (sub_sel & sub399) | (and_sel & and399) | (or_sel & or399);
  assign y400 = (add_sel & s400) | (sub_sel & sub400) | (and_sel & and400) | (or_sel & or400);
  assign y401 = (add_sel & s401) | (sub_sel & sub401) | (and_sel & and401) | (or_sel & or401);
  assign y402 = (add_sel & s402) | (sub_sel & sub402) | (and_sel & and402) | (or_sel & or402);
  assign y403 = (add_sel & s403) | (sub_sel & sub403) | (and_sel & and403) | (or_sel & or403);
  assign y404 = (add_sel & s404) | (sub_sel & sub404) | (and_sel & and404) | (or_sel & or404);
  assign y405 = (add_sel & s405) | (sub_sel & sub405) | (and_sel & and405) | (or_sel & or405);
  assign y406 = (add_sel & s406) | (sub_sel & sub406) | (and_sel & and406) | (or_sel & or406);
  assign y407 = (add_sel & s407) | (sub_sel & sub407) | (and_sel & and407) | (or_sel & or407);
  assign y408 = (add_sel & s408) | (sub_sel & sub408) | (and_sel & and408) | (or_sel & or408);
  assign y409 = (add_sel & s409) | (sub_sel & sub409) | (and_sel & and409) | (or_sel & or409);
  assign y410 = (add_sel & s410) | (sub_sel & sub410) | (and_sel & and410) | (or_sel & or410);
  assign y411 = (add_sel & s411) | (sub_sel & sub411) | (and_sel & and411) | (or_sel & or411);
  assign y412 = (add_sel & s412) | (sub_sel & sub412) | (and_sel & and412) | (or_sel & or412);
  assign y413 = (add_sel & s413) | (sub_sel & sub413) | (and_sel & and413) | (or_sel & or413);
  assign y414 = (add_sel & s414) | (sub_sel & sub414) | (and_sel & and414) | (or_sel & or414);
  assign y415 = (add_sel & s415) | (sub_sel & sub415) | (and_sel & and415) | (or_sel & or415);
  assign y416 = (add_sel & s416) | (sub_sel & sub416) | (and_sel & and416) | (or_sel & or416);
  assign y417 = (add_sel & s417) | (sub_sel & sub417) | (and_sel & and417) | (or_sel & or417);
  assign y418 = (add_sel & s418) | (sub_sel & sub418) | (and_sel & and418) | (or_sel & or418);
  assign y419 = (add_sel & s419) | (sub_sel & sub419) | (and_sel & and419) | (or_sel & or419);
  assign y420 = (add_sel & s420) | (sub_sel & sub420) | (and_sel & and420) | (or_sel & or420);
  assign y421 = (add_sel & s421) | (sub_sel & sub421) | (and_sel & and421) | (or_sel & or421);
  assign y422 = (add_sel & s422) | (sub_sel & sub422) | (and_sel & and422) | (or_sel & or422);
  assign y423 = (add_sel & s423) | (sub_sel & sub423) | (and_sel & and423) | (or_sel & or423);
  assign y424 = (add_sel & s424) | (sub_sel & sub424) | (and_sel & and424) | (or_sel & or424);
  assign y425 = (add_sel & s425) | (sub_sel & sub425) | (and_sel & and425) | (or_sel & or425);
  assign y426 = (add_sel & s426) | (sub_sel & sub426) | (and_sel & and426) | (or_sel & or426);
  assign y427 = (add_sel & s427) | (sub_sel & sub427) | (and_sel & and427) | (or_sel & or427);
  assign y428 = (add_sel & s428) | (sub_sel & sub428) | (and_sel & and428) | (or_sel & or428);
  assign y429 = (add_sel & s429) | (sub_sel & sub429) | (and_sel & and429) | (or_sel & or429);
  assign y430 = (add_sel & s430) | (sub_sel & sub430) | (and_sel & and430) | (or_sel & or430);
  assign y431 = (add_sel & s431) | (sub_sel & sub431) | (and_sel & and431) | (or_sel & or431);
  assign y432 = (add_sel & s432) | (sub_sel & sub432) | (and_sel & and432) | (or_sel & or432);
  assign y433 = (add_sel & s433) | (sub_sel & sub433) | (and_sel & and433) | (or_sel & or433);
  assign y434 = (add_sel & s434) | (sub_sel & sub434) | (and_sel & and434) | (or_sel & or434);
  assign y435 = (add_sel & s435) | (sub_sel & sub435) | (and_sel & and435) | (or_sel & or435);
  assign y436 = (add_sel & s436) | (sub_sel & sub436) | (and_sel & and436) | (or_sel & or436);
  assign y437 = (add_sel & s437) | (sub_sel & sub437) | (and_sel & and437) | (or_sel & or437);
  assign y438 = (add_sel & s438) | (sub_sel & sub438) | (and_sel & and438) | (or_sel & or438);
  assign y439 = (add_sel & s439) | (sub_sel & sub439) | (and_sel & and439) | (or_sel & or439);
  assign y440 = (add_sel & s440) | (sub_sel & sub440) | (and_sel & and440) | (or_sel & or440);
  assign y441 = (add_sel & s441) | (sub_sel & sub441) | (and_sel & and441) | (or_sel & or441);
  assign y442 = (add_sel & s442) | (sub_sel & sub442) | (and_sel & and442) | (or_sel & or442);
  assign y443 = (add_sel & s443) | (sub_sel & sub443) | (and_sel & and443) | (or_sel & or443);
  assign y444 = (add_sel & s444) | (sub_sel & sub444) | (and_sel & and444) | (or_sel & or444);
  assign y445 = (add_sel & s445) | (sub_sel & sub445) | (and_sel & and445) | (or_sel & or445);
  assign y446 = (add_sel & s446) | (sub_sel & sub446) | (and_sel & and446) | (or_sel & or446);
  assign y447 = (add_sel & s447) | (sub_sel & sub447) | (and_sel & and447) | (or_sel & or447);
  assign y448 = (add_sel & s448) | (sub_sel & sub448) | (and_sel & and448) | (or_sel & or448);
  assign y449 = (add_sel & s449) | (sub_sel & sub449) | (and_sel & and449) | (or_sel & or449);
  assign y450 = (add_sel & s450) | (sub_sel & sub450) | (and_sel & and450) | (or_sel & or450);
  assign y451 = (add_sel & s451) | (sub_sel & sub451) | (and_sel & and451) | (or_sel & or451);
  assign y452 = (add_sel & s452) | (sub_sel & sub452) | (and_sel & and452) | (or_sel & or452);
  assign y453 = (add_sel & s453) | (sub_sel & sub453) | (and_sel & and453) | (or_sel & or453);
  assign y454 = (add_sel & s454) | (sub_sel & sub454) | (and_sel & and454) | (or_sel & or454);
  assign y455 = (add_sel & s455) | (sub_sel & sub455) | (and_sel & and455) | (or_sel & or455);
  assign y456 = (add_sel & s456) | (sub_sel & sub456) | (and_sel & and456) | (or_sel & or456);
  assign y457 = (add_sel & s457) | (sub_sel & sub457) | (and_sel & and457) | (or_sel & or457);
  assign y458 = (add_sel & s458) | (sub_sel & sub458) | (and_sel & and458) | (or_sel & or458);
  assign y459 = (add_sel & s459) | (sub_sel & sub459) | (and_sel & and459) | (or_sel & or459);
  assign y460 = (add_sel & s460) | (sub_sel & sub460) | (and_sel & and460) | (or_sel & or460);
  assign y461 = (add_sel & s461) | (sub_sel & sub461) | (and_sel & and461) | (or_sel & or461);
  assign y462 = (add_sel & s462) | (sub_sel & sub462) | (and_sel & and462) | (or_sel & or462);
  assign y463 = (add_sel & s463) | (sub_sel & sub463) | (and_sel & and463) | (or_sel & or463);
  assign y464 = (add_sel & s464) | (sub_sel & sub464) | (and_sel & and464) | (or_sel & or464);
  assign y465 = (add_sel & s465) | (sub_sel & sub465) | (and_sel & and465) | (or_sel & or465);
  assign y466 = (add_sel & s466) | (sub_sel & sub466) | (and_sel & and466) | (or_sel & or466);
  assign y467 = (add_sel & s467) | (sub_sel & sub467) | (and_sel & and467) | (or_sel & or467);
  assign y468 = (add_sel & s468) | (sub_sel & sub468) | (and_sel & and468) | (or_sel & or468);
  assign y469 = (add_sel & s469) | (sub_sel & sub469) | (and_sel & and469) | (or_sel & or469);
  assign y470 = (add_sel & s470) | (sub_sel & sub470) | (and_sel & and470) | (or_sel & or470);
  assign y471 = (add_sel & s471) | (sub_sel & sub471) | (and_sel & and471) | (or_sel & or471);
  assign y472 = (add_sel & s472) | (sub_sel & sub472) | (and_sel & and472) | (or_sel & or472);
  assign y473 = (add_sel & s473) | (sub_sel & sub473) | (and_sel & and473) | (or_sel & or473);
  assign y474 = (add_sel & s474) | (sub_sel & sub474) | (and_sel & and474) | (or_sel & or474);
  assign y475 = (add_sel & s475) | (sub_sel & sub475) | (and_sel & and475) | (or_sel & or475);
  assign y476 = (add_sel & s476) | (sub_sel & sub476) | (and_sel & and476) | (or_sel & or476);
  assign y477 = (add_sel & s477) | (sub_sel & sub477) | (and_sel & and477) | (or_sel & or477);
  assign y478 = (add_sel & s478) | (sub_sel & sub478) | (and_sel & and478) | (or_sel & or478);
  assign y479 = (add_sel & s479) | (sub_sel & sub479) | (and_sel & and479) | (or_sel & or479);
  assign y480 = (add_sel & s480) | (sub_sel & sub480) | (and_sel & and480) | (or_sel & or480);
  assign y481 = (add_sel & s481) | (sub_sel & sub481) | (and_sel & and481) | (or_sel & or481);
  assign y482 = (add_sel & s482) | (sub_sel & sub482) | (and_sel & and482) | (or_sel & or482);
  assign y483 = (add_sel & s483) | (sub_sel & sub483) | (and_sel & and483) | (or_sel & or483);
  assign y484 = (add_sel & s484) | (sub_sel & sub484) | (and_sel & and484) | (or_sel & or484);
  assign y485 = (add_sel & s485) | (sub_sel & sub485) | (and_sel & and485) | (or_sel & or485);
  assign y486 = (add_sel & s486) | (sub_sel & sub486) | (and_sel & and486) | (or_sel & or486);
  assign y487 = (add_sel & s487) | (sub_sel & sub487) | (and_sel & and487) | (or_sel & or487);
  assign y488 = (add_sel & s488) | (sub_sel & sub488) | (and_sel & and488) | (or_sel & or488);
  assign y489 = (add_sel & s489) | (sub_sel & sub489) | (and_sel & and489) | (or_sel & or489);
  assign y490 = (add_sel & s490) | (sub_sel & sub490) | (and_sel & and490) | (or_sel & or490);
  assign y491 = (add_sel & s491) | (sub_sel & sub491) | (and_sel & and491) | (or_sel & or491);
  assign y492 = (add_sel & s492) | (sub_sel & sub492) | (and_sel & and492) | (or_sel & or492);
  assign y493 = (add_sel & s493) | (sub_sel & sub493) | (and_sel & and493) | (or_sel & or493);
  assign y494 = (add_sel & s494) | (sub_sel & sub494) | (and_sel & and494) | (or_sel & or494);
  assign y495 = (add_sel & s495) | (sub_sel & sub495) | (and_sel & and495) | (or_sel & or495);
  assign y496 = (add_sel & s496) | (sub_sel & sub496) | (and_sel & and496) | (or_sel & or496);
  assign y497 = (add_sel & s497) | (sub_sel & sub497) | (and_sel & and497) | (or_sel & or497);
  assign y498 = (add_sel & s498) | (sub_sel & sub498) | (and_sel & and498) | (or_sel & or498);
  assign y499 = (add_sel & s499) | (sub_sel & sub499) | (and_sel & and499) | (or_sel & or499);
  assign y500 = (add_sel & s500) | (sub_sel & sub500) | (and_sel & and500) | (or_sel & or500);
  assign y501 = (add_sel & s501) | (sub_sel & sub501) | (and_sel & and501) | (or_sel & or501);
  assign y502 = (add_sel & s502) | (sub_sel & sub502) | (and_sel & and502) | (or_sel & or502);
  assign y503 = (add_sel & s503) | (sub_sel & sub503) | (and_sel & and503) | (or_sel & or503);
  assign y504 = (add_sel & s504) | (sub_sel & sub504) | (and_sel & and504) | (or_sel & or504);
  assign y505 = (add_sel & s505) | (sub_sel & sub505) | (and_sel & and505) | (or_sel & or505);
  assign y506 = (add_sel & s506) | (sub_sel & sub506) | (and_sel & and506) | (or_sel & or506);
  assign y507 = (add_sel & s507) | (sub_sel & sub507) | (and_sel & and507) | (or_sel & or507);
  assign y508 = (add_sel & s508) | (sub_sel & sub508) | (and_sel & and508) | (or_sel & or508);
  assign y509 = (add_sel & s509) | (sub_sel & sub509) | (and_sel & and509) | (or_sel & or509);
  assign y510 = (add_sel & s510) | (sub_sel & sub510) | (and_sel & and510) | (or_sel & or510);
  assign y511 = (add_sel & s511) | (sub_sel & sub511) | (and_sel & and511) | (or_sel & or511);
  assign y512 = (add_sel & s512) | (sub_sel & sub512) | (and_sel & and512) | (or_sel & or512);
  assign y513 = (add_sel & s513) | (sub_sel & sub513) | (and_sel & and513) | (or_sel & or513);
  assign y514 = (add_sel & s514) | (sub_sel & sub514) | (and_sel & and514) | (or_sel & or514);
  assign y515 = (add_sel & s515) | (sub_sel & sub515) | (and_sel & and515) | (or_sel & or515);
  assign y516 = (add_sel & s516) | (sub_sel & sub516) | (and_sel & and516) | (or_sel & or516);
  assign y517 = (add_sel & s517) | (sub_sel & sub517) | (and_sel & and517) | (or_sel & or517);
  assign y518 = (add_sel & s518) | (sub_sel & sub518) | (and_sel & and518) | (or_sel & or518);
  assign y519 = (add_sel & s519) | (sub_sel & sub519) | (and_sel & and519) | (or_sel & or519);
  assign y520 = (add_sel & s520) | (sub_sel & sub520) | (and_sel & and520) | (or_sel & or520);
  assign y521 = (add_sel & s521) | (sub_sel & sub521) | (and_sel & and521) | (or_sel & or521);
  assign y522 = (add_sel & s522) | (sub_sel & sub522) | (and_sel & and522) | (or_sel & or522);
  assign y523 = (add_sel & s523) | (sub_sel & sub523) | (and_sel & and523) | (or_sel & or523);
  assign y524 = (add_sel & s524) | (sub_sel & sub524) | (and_sel & and524) | (or_sel & or524);
  assign y525 = (add_sel & s525) | (sub_sel & sub525) | (and_sel & and525) | (or_sel & or525);
  assign y526 = (add_sel & s526) | (sub_sel & sub526) | (and_sel & and526) | (or_sel & or526);
  assign y527 = (add_sel & s527) | (sub_sel & sub527) | (and_sel & and527) | (or_sel & or527);
  assign y528 = (add_sel & s528) | (sub_sel & sub528) | (and_sel & and528) | (or_sel & or528);
  assign y529 = (add_sel & s529) | (sub_sel & sub529) | (and_sel & and529) | (or_sel & or529);
  assign y530 = (add_sel & s530) | (sub_sel & sub530) | (and_sel & and530) | (or_sel & or530);
  assign y531 = (add_sel & s531) | (sub_sel & sub531) | (and_sel & and531) | (or_sel & or531);
  assign y532 = (add_sel & s532) | (sub_sel & sub532) | (and_sel & and532) | (or_sel & or532);
  assign y533 = (add_sel & s533) | (sub_sel & sub533) | (and_sel & and533) | (or_sel & or533);
  assign y534 = (add_sel & s534) | (sub_sel & sub534) | (and_sel & and534) | (or_sel & or534);
  assign y535 = (add_sel & s535) | (sub_sel & sub535) | (and_sel & and535) | (or_sel & or535);
  assign y536 = (add_sel & s536) | (sub_sel & sub536) | (and_sel & and536) | (or_sel & or536);
  assign y537 = (add_sel & s537) | (sub_sel & sub537) | (and_sel & and537) | (or_sel & or537);
  assign y538 = (add_sel & s538) | (sub_sel & sub538) | (and_sel & and538) | (or_sel & or538);
  assign y539 = (add_sel & s539) | (sub_sel & sub539) | (and_sel & and539) | (or_sel & or539);
  assign y540 = (add_sel & s540) | (sub_sel & sub540) | (and_sel & and540) | (or_sel & or540);
  assign y541 = (add_sel & s541) | (sub_sel & sub541) | (and_sel & and541) | (or_sel & or541);
  assign y542 = (add_sel & s542) | (sub_sel & sub542) | (and_sel & and542) | (or_sel & or542);
  assign y543 = (add_sel & s543) | (sub_sel & sub543) | (and_sel & and543) | (or_sel & or543);
  assign y544 = (add_sel & s544) | (sub_sel & sub544) | (and_sel & and544) | (or_sel & or544);
  assign y545 = (add_sel & s545) | (sub_sel & sub545) | (and_sel & and545) | (or_sel & or545);
  assign y546 = (add_sel & s546) | (sub_sel & sub546) | (and_sel & and546) | (or_sel & or546);
  assign y547 = (add_sel & s547) | (sub_sel & sub547) | (and_sel & and547) | (or_sel & or547);
  assign y548 = (add_sel & s548) | (sub_sel & sub548) | (and_sel & and548) | (or_sel & or548);
  assign y549 = (add_sel & s549) | (sub_sel & sub549) | (and_sel & and549) | (or_sel & or549);
  assign y550 = (add_sel & s550) | (sub_sel & sub550) | (and_sel & and550) | (or_sel & or550);
  assign y551 = (add_sel & s551) | (sub_sel & sub551) | (and_sel & and551) | (or_sel & or551);
  assign y552 = (add_sel & s552) | (sub_sel & sub552) | (and_sel & and552) | (or_sel & or552);
  assign y553 = (add_sel & s553) | (sub_sel & sub553) | (and_sel & and553) | (or_sel & or553);
  assign y554 = (add_sel & s554) | (sub_sel & sub554) | (and_sel & and554) | (or_sel & or554);
  assign y555 = (add_sel & s555) | (sub_sel & sub555) | (and_sel & and555) | (or_sel & or555);
  assign y556 = (add_sel & s556) | (sub_sel & sub556) | (and_sel & and556) | (or_sel & or556);
  assign y557 = (add_sel & s557) | (sub_sel & sub557) | (and_sel & and557) | (or_sel & or557);
  assign y558 = (add_sel & s558) | (sub_sel & sub558) | (and_sel & and558) | (or_sel & or558);
  assign y559 = (add_sel & s559) | (sub_sel & sub559) | (and_sel & and559) | (or_sel & or559);
  assign y560 = (add_sel & s560) | (sub_sel & sub560) | (and_sel & and560) | (or_sel & or560);
  assign y561 = (add_sel & s561) | (sub_sel & sub561) | (and_sel & and561) | (or_sel & or561);
  assign y562 = (add_sel & s562) | (sub_sel & sub562) | (and_sel & and562) | (or_sel & or562);
  assign y563 = (add_sel & s563) | (sub_sel & sub563) | (and_sel & and563) | (or_sel & or563);
  assign y564 = (add_sel & s564) | (sub_sel & sub564) | (and_sel & and564) | (or_sel & or564);
  assign y565 = (add_sel & s565) | (sub_sel & sub565) | (and_sel & and565) | (or_sel & or565);
  assign y566 = (add_sel & s566) | (sub_sel & sub566) | (and_sel & and566) | (or_sel & or566);
  assign y567 = (add_sel & s567) | (sub_sel & sub567) | (and_sel & and567) | (or_sel & or567);
  assign y568 = (add_sel & s568) | (sub_sel & sub568) | (and_sel & and568) | (or_sel & or568);
  assign y569 = (add_sel & s569) | (sub_sel & sub569) | (and_sel & and569) | (or_sel & or569);
  assign y570 = (add_sel & s570) | (sub_sel & sub570) | (and_sel & and570) | (or_sel & or570);
  assign y571 = (add_sel & s571) | (sub_sel & sub571) | (and_sel & and571) | (or_sel & or571);
  assign y572 = (add_sel & s572) | (sub_sel & sub572) | (and_sel & and572) | (or_sel & or572);
  assign y573 = (add_sel & s573) | (sub_sel & sub573) | (and_sel & and573) | (or_sel & or573);
  assign y574 = (add_sel & s574) | (sub_sel & sub574) | (and_sel & and574) | (or_sel & or574);
  assign y575 = (add_sel & s575) | (sub_sel & sub575) | (and_sel & and575) | (or_sel & or575);
  assign y576 = (add_sel & s576) | (sub_sel & sub576) | (and_sel & and576) | (or_sel & or576);
  assign y577 = (add_sel & s577) | (sub_sel & sub577) | (and_sel & and577) | (or_sel & or577);
  assign y578 = (add_sel & s578) | (sub_sel & sub578) | (and_sel & and578) | (or_sel & or578);
  assign y579 = (add_sel & s579) | (sub_sel & sub579) | (and_sel & and579) | (or_sel & or579);
  assign y580 = (add_sel & s580) | (sub_sel & sub580) | (and_sel & and580) | (or_sel & or580);
  assign y581 = (add_sel & s581) | (sub_sel & sub581) | (and_sel & and581) | (or_sel & or581);
  assign y582 = (add_sel & s582) | (sub_sel & sub582) | (and_sel & and582) | (or_sel & or582);
  assign y583 = (add_sel & s583) | (sub_sel & sub583) | (and_sel & and583) | (or_sel & or583);
  assign y584 = (add_sel & s584) | (sub_sel & sub584) | (and_sel & and584) | (or_sel & or584);
  assign y585 = (add_sel & s585) | (sub_sel & sub585) | (and_sel & and585) | (or_sel & or585);
  assign y586 = (add_sel & s586) | (sub_sel & sub586) | (and_sel & and586) | (or_sel & or586);
  assign y587 = (add_sel & s587) | (sub_sel & sub587) | (and_sel & and587) | (or_sel & or587);
  assign y588 = (add_sel & s588) | (sub_sel & sub588) | (and_sel & and588) | (or_sel & or588);
  assign y589 = (add_sel & s589) | (sub_sel & sub589) | (and_sel & and589) | (or_sel & or589);
  assign y590 = (add_sel & s590) | (sub_sel & sub590) | (and_sel & and590) | (or_sel & or590);
  assign y591 = (add_sel & s591) | (sub_sel & sub591) | (and_sel & and591) | (or_sel & or591);
  assign y592 = (add_sel & s592) | (sub_sel & sub592) | (and_sel & and592) | (or_sel & or592);
  assign y593 = (add_sel & s593) | (sub_sel & sub593) | (and_sel & and593) | (or_sel & or593);
  assign y594 = (add_sel & s594) | (sub_sel & sub594) | (and_sel & and594) | (or_sel & or594);
  assign y595 = (add_sel & s595) | (sub_sel & sub595) | (and_sel & and595) | (or_sel & or595);
  assign y596 = (add_sel & s596) | (sub_sel & sub596) | (and_sel & and596) | (or_sel & or596);
  assign y597 = (add_sel & s597) | (sub_sel & sub597) | (and_sel & and597) | (or_sel & or597);
  assign y598 = (add_sel & s598) | (sub_sel & sub598) | (and_sel & and598) | (or_sel & or598);
  assign y599 = (add_sel & s599) | (sub_sel & sub599) | (and_sel & and599) | (or_sel & or599);
  assign y600 = (add_sel & s600) | (sub_sel & sub600) | (and_sel & and600) | (or_sel & or600);
  assign y601 = (add_sel & s601) | (sub_sel & sub601) | (and_sel & and601) | (or_sel & or601);
  assign y602 = (add_sel & s602) | (sub_sel & sub602) | (and_sel & and602) | (or_sel & or602);
  assign y603 = (add_sel & s603) | (sub_sel & sub603) | (and_sel & and603) | (or_sel & or603);
  assign y604 = (add_sel & s604) | (sub_sel & sub604) | (and_sel & and604) | (or_sel & or604);
  assign y605 = (add_sel & s605) | (sub_sel & sub605) | (and_sel & and605) | (or_sel & or605);
  assign y606 = (add_sel & s606) | (sub_sel & sub606) | (and_sel & and606) | (or_sel & or606);
  assign y607 = (add_sel & s607) | (sub_sel & sub607) | (and_sel & and607) | (or_sel & or607);
  assign y608 = (add_sel & s608) | (sub_sel & sub608) | (and_sel & and608) | (or_sel & or608);
  assign y609 = (add_sel & s609) | (sub_sel & sub609) | (and_sel & and609) | (or_sel & or609);
  assign y610 = (add_sel & s610) | (sub_sel & sub610) | (and_sel & and610) | (or_sel & or610);
  assign y611 = (add_sel & s611) | (sub_sel & sub611) | (and_sel & and611) | (or_sel & or611);
  assign y612 = (add_sel & s612) | (sub_sel & sub612) | (and_sel & and612) | (or_sel & or612);
  assign y613 = (add_sel & s613) | (sub_sel & sub613) | (and_sel & and613) | (or_sel & or613);
  assign y614 = (add_sel & s614) | (sub_sel & sub614) | (and_sel & and614) | (or_sel & or614);
  assign y615 = (add_sel & s615) | (sub_sel & sub615) | (and_sel & and615) | (or_sel & or615);
  assign y616 = (add_sel & s616) | (sub_sel & sub616) | (and_sel & and616) | (or_sel & or616);
  assign y617 = (add_sel & s617) | (sub_sel & sub617) | (and_sel & and617) | (or_sel & or617);
  assign y618 = (add_sel & s618) | (sub_sel & sub618) | (and_sel & and618) | (or_sel & or618);
  assign y619 = (add_sel & s619) | (sub_sel & sub619) | (and_sel & and619) | (or_sel & or619);
  assign y620 = (add_sel & s620) | (sub_sel & sub620) | (and_sel & and620) | (or_sel & or620);
  assign y621 = (add_sel & s621) | (sub_sel & sub621) | (and_sel & and621) | (or_sel & or621);
  assign y622 = (add_sel & s622) | (sub_sel & sub622) | (and_sel & and622) | (or_sel & or622);
  assign y623 = (add_sel & s623) | (sub_sel & sub623) | (and_sel & and623) | (or_sel & or623);
  assign y624 = (add_sel & s624) | (sub_sel & sub624) | (and_sel & and624) | (or_sel & or624);
  assign y625 = (add_sel & s625) | (sub_sel & sub625) | (and_sel & and625) | (or_sel & or625);
  assign y626 = (add_sel & s626) | (sub_sel & sub626) | (and_sel & and626) | (or_sel & or626);
  assign y627 = (add_sel & s627) | (sub_sel & sub627) | (and_sel & and627) | (or_sel & or627);
  assign y628 = (add_sel & s628) | (sub_sel & sub628) | (and_sel & and628) | (or_sel & or628);
  assign y629 = (add_sel & s629) | (sub_sel & sub629) | (and_sel & and629) | (or_sel & or629);
  assign y630 = (add_sel & s630) | (sub_sel & sub630) | (and_sel & and630) | (or_sel & or630);
  assign y631 = (add_sel & s631) | (sub_sel & sub631) | (and_sel & and631) | (or_sel & or631);
  assign y632 = (add_sel & s632) | (sub_sel & sub632) | (and_sel & and632) | (or_sel & or632);
  assign y633 = (add_sel & s633) | (sub_sel & sub633) | (and_sel & and633) | (or_sel & or633);
  assign y634 = (add_sel & s634) | (sub_sel & sub634) | (and_sel & and634) | (or_sel & or634);
  assign y635 = (add_sel & s635) | (sub_sel & sub635) | (and_sel & and635) | (or_sel & or635);
  assign y636 = (add_sel & s636) | (sub_sel & sub636) | (and_sel & and636) | (or_sel & or636);
  assign y637 = (add_sel & s637) | (sub_sel & sub637) | (and_sel & and637) | (or_sel & or637);
  assign y638 = (add_sel & s638) | (sub_sel & sub638) | (and_sel & and638) | (or_sel & or638);
  assign y639 = (add_sel & s639) | (sub_sel & sub639) | (and_sel & and639) | (or_sel & or639);
  assign y640 = (add_sel & s640) | (sub_sel & sub640) | (and_sel & and640) | (or_sel & or640);
  assign y641 = (add_sel & s641) | (sub_sel & sub641) | (and_sel & and641) | (or_sel & or641);
  assign y642 = (add_sel & s642) | (sub_sel & sub642) | (and_sel & and642) | (or_sel & or642);
  assign y643 = (add_sel & s643) | (sub_sel & sub643) | (and_sel & and643) | (or_sel & or643);
  assign y644 = (add_sel & s644) | (sub_sel & sub644) | (and_sel & and644) | (or_sel & or644);
  assign y645 = (add_sel & s645) | (sub_sel & sub645) | (and_sel & and645) | (or_sel & or645);
  assign y646 = (add_sel & s646) | (sub_sel & sub646) | (and_sel & and646) | (or_sel & or646);
  assign y647 = (add_sel & s647) | (sub_sel & sub647) | (and_sel & and647) | (or_sel & or647);
  assign y648 = (add_sel & s648) | (sub_sel & sub648) | (and_sel & and648) | (or_sel & or648);
  assign y649 = (add_sel & s649) | (sub_sel & sub649) | (and_sel & and649) | (or_sel & or649);
  assign y650 = (add_sel & s650) | (sub_sel & sub650) | (and_sel & and650) | (or_sel & or650);
  assign y651 = (add_sel & s651) | (sub_sel & sub651) | (and_sel & and651) | (or_sel & or651);
  assign y652 = (add_sel & s652) | (sub_sel & sub652) | (and_sel & and652) | (or_sel & or652);
  assign y653 = (add_sel & s653) | (sub_sel & sub653) | (and_sel & and653) | (or_sel & or653);
  assign y654 = (add_sel & s654) | (sub_sel & sub654) | (and_sel & and654) | (or_sel & or654);
  assign y655 = (add_sel & s655) | (sub_sel & sub655) | (and_sel & and655) | (or_sel & or655);
  assign y656 = (add_sel & s656) | (sub_sel & sub656) | (and_sel & and656) | (or_sel & or656);
  assign y657 = (add_sel & s657) | (sub_sel & sub657) | (and_sel & and657) | (or_sel & or657);
  assign y658 = (add_sel & s658) | (sub_sel & sub658) | (and_sel & and658) | (or_sel & or658);
  assign y659 = (add_sel & s659) | (sub_sel & sub659) | (and_sel & and659) | (or_sel & or659);
  assign y660 = (add_sel & s660) | (sub_sel & sub660) | (and_sel & and660) | (or_sel & or660);
  assign y661 = (add_sel & s661) | (sub_sel & sub661) | (and_sel & and661) | (or_sel & or661);
  assign y662 = (add_sel & s662) | (sub_sel & sub662) | (and_sel & and662) | (or_sel & or662);
  assign y663 = (add_sel & s663) | (sub_sel & sub663) | (and_sel & and663) | (or_sel & or663);
  assign y664 = (add_sel & s664) | (sub_sel & sub664) | (and_sel & and664) | (or_sel & or664);
  assign y665 = (add_sel & s665) | (sub_sel & sub665) | (and_sel & and665) | (or_sel & or665);
  assign y666 = (add_sel & s666) | (sub_sel & sub666) | (and_sel & and666) | (or_sel & or666);
  assign y667 = (add_sel & s667) | (sub_sel & sub667) | (and_sel & and667) | (or_sel & or667);
  assign y668 = (add_sel & s668) | (sub_sel & sub668) | (and_sel & and668) | (or_sel & or668);
  assign y669 = (add_sel & s669) | (sub_sel & sub669) | (and_sel & and669) | (or_sel & or669);
  assign y670 = (add_sel & s670) | (sub_sel & sub670) | (and_sel & and670) | (or_sel & or670);
  assign y671 = (add_sel & s671) | (sub_sel & sub671) | (and_sel & and671) | (or_sel & or671);
  assign y672 = (add_sel & s672) | (sub_sel & sub672) | (and_sel & and672) | (or_sel & or672);
  assign y673 = (add_sel & s673) | (sub_sel & sub673) | (and_sel & and673) | (or_sel & or673);
  assign y674 = (add_sel & s674) | (sub_sel & sub674) | (and_sel & and674) | (or_sel & or674);
  assign y675 = (add_sel & s675) | (sub_sel & sub675) | (and_sel & and675) | (or_sel & or675);
  assign y676 = (add_sel & s676) | (sub_sel & sub676) | (and_sel & and676) | (or_sel & or676);
  assign y677 = (add_sel & s677) | (sub_sel & sub677) | (and_sel & and677) | (or_sel & or677);
  assign y678 = (add_sel & s678) | (sub_sel & sub678) | (and_sel & and678) | (or_sel & or678);
  assign y679 = (add_sel & s679) | (sub_sel & sub679) | (and_sel & and679) | (or_sel & or679);
  assign y680 = (add_sel & s680) | (sub_sel & sub680) | (and_sel & and680) | (or_sel & or680);
  assign y681 = (add_sel & s681) | (sub_sel & sub681) | (and_sel & and681) | (or_sel & or681);
  assign y682 = (add_sel & s682) | (sub_sel & sub682) | (and_sel & and682) | (or_sel & or682);
  assign y683 = (add_sel & s683) | (sub_sel & sub683) | (and_sel & and683) | (or_sel & or683);
  assign y684 = (add_sel & s684) | (sub_sel & sub684) | (and_sel & and684) | (or_sel & or684);
  assign y685 = (add_sel & s685) | (sub_sel & sub685) | (and_sel & and685) | (or_sel & or685);
  assign y686 = (add_sel & s686) | (sub_sel & sub686) | (and_sel & and686) | (or_sel & or686);
  assign y687 = (add_sel & s687) | (sub_sel & sub687) | (and_sel & and687) | (or_sel & or687);
  assign y688 = (add_sel & s688) | (sub_sel & sub688) | (and_sel & and688) | (or_sel & or688);
  assign y689 = (add_sel & s689) | (sub_sel & sub689) | (and_sel & and689) | (or_sel & or689);
  assign y690 = (add_sel & s690) | (sub_sel & sub690) | (and_sel & and690) | (or_sel & or690);
  assign y691 = (add_sel & s691) | (sub_sel & sub691) | (and_sel & and691) | (or_sel & or691);
  assign y692 = (add_sel & s692) | (sub_sel & sub692) | (and_sel & and692) | (or_sel & or692);
  assign y693 = (add_sel & s693) | (sub_sel & sub693) | (and_sel & and693) | (or_sel & or693);
  assign y694 = (add_sel & s694) | (sub_sel & sub694) | (and_sel & and694) | (or_sel & or694);
  assign y695 = (add_sel & s695) | (sub_sel & sub695) | (and_sel & and695) | (or_sel & or695);
  assign y696 = (add_sel & s696) | (sub_sel & sub696) | (and_sel & and696) | (or_sel & or696);
  assign y697 = (add_sel & s697) | (sub_sel & sub697) | (and_sel & and697) | (or_sel & or697);
  assign y698 = (add_sel & s698) | (sub_sel & sub698) | (and_sel & and698) | (or_sel & or698);
  assign y699 = (add_sel & s699) | (sub_sel & sub699) | (and_sel & and699) | (or_sel & or699);
  assign y700 = (add_sel & s700) | (sub_sel & sub700) | (and_sel & and700) | (or_sel & or700);
  assign y701 = (add_sel & s701) | (sub_sel & sub701) | (and_sel & and701) | (or_sel & or701);
  assign y702 = (add_sel & s702) | (sub_sel & sub702) | (and_sel & and702) | (or_sel & or702);
  assign y703 = (add_sel & s703) | (sub_sel & sub703) | (and_sel & and703) | (or_sel & or703);
  assign y704 = (add_sel & s704) | (sub_sel & sub704) | (and_sel & and704) | (or_sel & or704);
  assign y705 = (add_sel & s705) | (sub_sel & sub705) | (and_sel & and705) | (or_sel & or705);
  assign y706 = (add_sel & s706) | (sub_sel & sub706) | (and_sel & and706) | (or_sel & or706);
  assign y707 = (add_sel & s707) | (sub_sel & sub707) | (and_sel & and707) | (or_sel & or707);
  assign y708 = (add_sel & s708) | (sub_sel & sub708) | (and_sel & and708) | (or_sel & or708);
  assign y709 = (add_sel & s709) | (sub_sel & sub709) | (and_sel & and709) | (or_sel & or709);
  assign y710 = (add_sel & s710) | (sub_sel & sub710) | (and_sel & and710) | (or_sel & or710);
  assign y711 = (add_sel & s711) | (sub_sel & sub711) | (and_sel & and711) | (or_sel & or711);
  assign y712 = (add_sel & s712) | (sub_sel & sub712) | (and_sel & and712) | (or_sel & or712);
  assign y713 = (add_sel & s713) | (sub_sel & sub713) | (and_sel & and713) | (or_sel & or713);
  assign y714 = (add_sel & s714) | (sub_sel & sub714) | (and_sel & and714) | (or_sel & or714);
  assign y715 = (add_sel & s715) | (sub_sel & sub715) | (and_sel & and715) | (or_sel & or715);
  assign y716 = (add_sel & s716) | (sub_sel & sub716) | (and_sel & and716) | (or_sel & or716);
  assign y717 = (add_sel & s717) | (sub_sel & sub717) | (and_sel & and717) | (or_sel & or717);
  assign y718 = (add_sel & s718) | (sub_sel & sub718) | (and_sel & and718) | (or_sel & or718);
  assign y719 = (add_sel & s719) | (sub_sel & sub719) | (and_sel & and719) | (or_sel & or719);
  assign y720 = (add_sel & s720) | (sub_sel & sub720) | (and_sel & and720) | (or_sel & or720);
  assign y721 = (add_sel & s721) | (sub_sel & sub721) | (and_sel & and721) | (or_sel & or721);
  assign y722 = (add_sel & s722) | (sub_sel & sub722) | (and_sel & and722) | (or_sel & or722);
  assign y723 = (add_sel & s723) | (sub_sel & sub723) | (and_sel & and723) | (or_sel & or723);
  assign y724 = (add_sel & s724) | (sub_sel & sub724) | (and_sel & and724) | (or_sel & or724);
  assign y725 = (add_sel & s725) | (sub_sel & sub725) | (and_sel & and725) | (or_sel & or725);
  assign y726 = (add_sel & s726) | (sub_sel & sub726) | (and_sel & and726) | (or_sel & or726);
  assign y727 = (add_sel & s727) | (sub_sel & sub727) | (and_sel & and727) | (or_sel & or727);
  assign y728 = (add_sel & s728) | (sub_sel & sub728) | (and_sel & and728) | (or_sel & or728);
  assign y729 = (add_sel & s729) | (sub_sel & sub729) | (and_sel & and729) | (or_sel & or729);
  assign y730 = (add_sel & s730) | (sub_sel & sub730) | (and_sel & and730) | (or_sel & or730);
  assign y731 = (add_sel & s731) | (sub_sel & sub731) | (and_sel & and731) | (or_sel & or731);
  assign y732 = (add_sel & s732) | (sub_sel & sub732) | (and_sel & and732) | (or_sel & or732);
  assign y733 = (add_sel & s733) | (sub_sel & sub733) | (and_sel & and733) | (or_sel & or733);
  assign y734 = (add_sel & s734) | (sub_sel & sub734) | (and_sel & and734) | (or_sel & or734);
  assign y735 = (add_sel & s735) | (sub_sel & sub735) | (and_sel & and735) | (or_sel & or735);
  assign y736 = (add_sel & s736) | (sub_sel & sub736) | (and_sel & and736) | (or_sel & or736);
  assign y737 = (add_sel & s737) | (sub_sel & sub737) | (and_sel & and737) | (or_sel & or737);
  assign y738 = (add_sel & s738) | (sub_sel & sub738) | (and_sel & and738) | (or_sel & or738);
  assign y739 = (add_sel & s739) | (sub_sel & sub739) | (and_sel & and739) | (or_sel & or739);
  assign y740 = (add_sel & s740) | (sub_sel & sub740) | (and_sel & and740) | (or_sel & or740);
  assign y741 = (add_sel & s741) | (sub_sel & sub741) | (and_sel & and741) | (or_sel & or741);
  assign y742 = (add_sel & s742) | (sub_sel & sub742) | (and_sel & and742) | (or_sel & or742);
  assign y743 = (add_sel & s743) | (sub_sel & sub743) | (and_sel & and743) | (or_sel & or743);
  assign y744 = (add_sel & s744) | (sub_sel & sub744) | (and_sel & and744) | (or_sel & or744);
  assign y745 = (add_sel & s745) | (sub_sel & sub745) | (and_sel & and745) | (or_sel & or745);
  assign y746 = (add_sel & s746) | (sub_sel & sub746) | (and_sel & and746) | (or_sel & or746);
  assign y747 = (add_sel & s747) | (sub_sel & sub747) | (and_sel & and747) | (or_sel & or747);
  assign y748 = (add_sel & s748) | (sub_sel & sub748) | (and_sel & and748) | (or_sel & or748);
  assign y749 = (add_sel & s749) | (sub_sel & sub749) | (and_sel & and749) | (or_sel & or749);
  assign y750 = (add_sel & s750) | (sub_sel & sub750) | (and_sel & and750) | (or_sel & or750);
  assign y751 = (add_sel & s751) | (sub_sel & sub751) | (and_sel & and751) | (or_sel & or751);
  assign y752 = (add_sel & s752) | (sub_sel & sub752) | (and_sel & and752) | (or_sel & or752);
  assign y753 = (add_sel & s753) | (sub_sel & sub753) | (and_sel & and753) | (or_sel & or753);
  assign y754 = (add_sel & s754) | (sub_sel & sub754) | (and_sel & and754) | (or_sel & or754);
  assign y755 = (add_sel & s755) | (sub_sel & sub755) | (and_sel & and755) | (or_sel & or755);
  assign y756 = (add_sel & s756) | (sub_sel & sub756) | (and_sel & and756) | (or_sel & or756);
  assign y757 = (add_sel & s757) | (sub_sel & sub757) | (and_sel & and757) | (or_sel & or757);
  assign y758 = (add_sel & s758) | (sub_sel & sub758) | (and_sel & and758) | (or_sel & or758);
  assign y759 = (add_sel & s759) | (sub_sel & sub759) | (and_sel & and759) | (or_sel & or759);
  assign y760 = (add_sel & s760) | (sub_sel & sub760) | (and_sel & and760) | (or_sel & or760);
  assign y761 = (add_sel & s761) | (sub_sel & sub761) | (and_sel & and761) | (or_sel & or761);
  assign y762 = (add_sel & s762) | (sub_sel & sub762) | (and_sel & and762) | (or_sel & or762);
  assign y763 = (add_sel & s763) | (sub_sel & sub763) | (and_sel & and763) | (or_sel & or763);
  assign y764 = (add_sel & s764) | (sub_sel & sub764) | (and_sel & and764) | (or_sel & or764);
  assign y765 = (add_sel & s765) | (sub_sel & sub765) | (and_sel & and765) | (or_sel & or765);
  assign y766 = (add_sel & s766) | (sub_sel & sub766) | (and_sel & and766) | (or_sel & or766);
  assign y767 = (add_sel & s767) | (sub_sel & sub767) | (and_sel & and767) | (or_sel & or767);
  assign y768 = (add_sel & s768) | (sub_sel & sub768) | (and_sel & and768) | (or_sel & or768);
  assign y769 = (add_sel & s769) | (sub_sel & sub769) | (and_sel & and769) | (or_sel & or769);
  assign y770 = (add_sel & s770) | (sub_sel & sub770) | (and_sel & and770) | (or_sel & or770);
  assign y771 = (add_sel & s771) | (sub_sel & sub771) | (and_sel & and771) | (or_sel & or771);
  assign y772 = (add_sel & s772) | (sub_sel & sub772) | (and_sel & and772) | (or_sel & or772);
  assign y773 = (add_sel & s773) | (sub_sel & sub773) | (and_sel & and773) | (or_sel & or773);
  assign y774 = (add_sel & s774) | (sub_sel & sub774) | (and_sel & and774) | (or_sel & or774);
  assign y775 = (add_sel & s775) | (sub_sel & sub775) | (and_sel & and775) | (or_sel & or775);
  assign y776 = (add_sel & s776) | (sub_sel & sub776) | (and_sel & and776) | (or_sel & or776);
  assign y777 = (add_sel & s777) | (sub_sel & sub777) | (and_sel & and777) | (or_sel & or777);
  assign y778 = (add_sel & s778) | (sub_sel & sub778) | (and_sel & and778) | (or_sel & or778);
  assign y779 = (add_sel & s779) | (sub_sel & sub779) | (and_sel & and779) | (or_sel & or779);
  assign y780 = (add_sel & s780) | (sub_sel & sub780) | (and_sel & and780) | (or_sel & or780);
  assign y781 = (add_sel & s781) | (sub_sel & sub781) | (and_sel & and781) | (or_sel & or781);
  assign y782 = (add_sel & s782) | (sub_sel & sub782) | (and_sel & and782) | (or_sel & or782);
  assign y783 = (add_sel & s783) | (sub_sel & sub783) | (and_sel & and783) | (or_sel & or783);
  assign y784 = (add_sel & s784) | (sub_sel & sub784) | (and_sel & and784) | (or_sel & or784);
  assign y785 = (add_sel & s785) | (sub_sel & sub785) | (and_sel & and785) | (or_sel & or785);
  assign y786 = (add_sel & s786) | (sub_sel & sub786) | (and_sel & and786) | (or_sel & or786);
  assign y787 = (add_sel & s787) | (sub_sel & sub787) | (and_sel & and787) | (or_sel & or787);
  assign y788 = (add_sel & s788) | (sub_sel & sub788) | (and_sel & and788) | (or_sel & or788);
  assign y789 = (add_sel & s789) | (sub_sel & sub789) | (and_sel & and789) | (or_sel & or789);
  assign y790 = (add_sel & s790) | (sub_sel & sub790) | (and_sel & and790) | (or_sel & or790);
  assign y791 = (add_sel & s791) | (sub_sel & sub791) | (and_sel & and791) | (or_sel & or791);
  assign y792 = (add_sel & s792) | (sub_sel & sub792) | (and_sel & and792) | (or_sel & or792);
  assign y793 = (add_sel & s793) | (sub_sel & sub793) | (and_sel & and793) | (or_sel & or793);
  assign y794 = (add_sel & s794) | (sub_sel & sub794) | (and_sel & and794) | (or_sel & or794);
  assign y795 = (add_sel & s795) | (sub_sel & sub795) | (and_sel & and795) | (or_sel & or795);
  assign y796 = (add_sel & s796) | (sub_sel & sub796) | (and_sel & and796) | (or_sel & or796);
  assign y797 = (add_sel & s797) | (sub_sel & sub797) | (and_sel & and797) | (or_sel & or797);
  assign y798 = (add_sel & s798) | (sub_sel & sub798) | (and_sel & and798) | (or_sel & or798);
  assign y799 = (add_sel & s799) | (sub_sel & sub799) | (and_sel & and799) | (or_sel & or799);
  assign y800 = (add_sel & s800) | (sub_sel & sub800) | (and_sel & and800) | (or_sel & or800);
  assign y801 = (add_sel & s801) | (sub_sel & sub801) | (and_sel & and801) | (or_sel & or801);
  assign y802 = (add_sel & s802) | (sub_sel & sub802) | (and_sel & and802) | (or_sel & or802);
  assign y803 = (add_sel & s803) | (sub_sel & sub803) | (and_sel & and803) | (or_sel & or803);
  assign y804 = (add_sel & s804) | (sub_sel & sub804) | (and_sel & and804) | (or_sel & or804);
  assign y805 = (add_sel & s805) | (sub_sel & sub805) | (and_sel & and805) | (or_sel & or805);
  assign y806 = (add_sel & s806) | (sub_sel & sub806) | (and_sel & and806) | (or_sel & or806);
  assign y807 = (add_sel & s807) | (sub_sel & sub807) | (and_sel & and807) | (or_sel & or807);
  assign y808 = (add_sel & s808) | (sub_sel & sub808) | (and_sel & and808) | (or_sel & or808);
  assign y809 = (add_sel & s809) | (sub_sel & sub809) | (and_sel & and809) | (or_sel & or809);
  assign y810 = (add_sel & s810) | (sub_sel & sub810) | (and_sel & and810) | (or_sel & or810);
  assign y811 = (add_sel & s811) | (sub_sel & sub811) | (and_sel & and811) | (or_sel & or811);
  assign y812 = (add_sel & s812) | (sub_sel & sub812) | (and_sel & and812) | (or_sel & or812);
  assign y813 = (add_sel & s813) | (sub_sel & sub813) | (and_sel & and813) | (or_sel & or813);
  assign y814 = (add_sel & s814) | (sub_sel & sub814) | (and_sel & and814) | (or_sel & or814);
  assign y815 = (add_sel & s815) | (sub_sel & sub815) | (and_sel & and815) | (or_sel & or815);
  assign y816 = (add_sel & s816) | (sub_sel & sub816) | (and_sel & and816) | (or_sel & or816);
  assign y817 = (add_sel & s817) | (sub_sel & sub817) | (and_sel & and817) | (or_sel & or817);
  assign y818 = (add_sel & s818) | (sub_sel & sub818) | (and_sel & and818) | (or_sel & or818);
  assign y819 = (add_sel & s819) | (sub_sel & sub819) | (and_sel & and819) | (or_sel & or819);
  assign y820 = (add_sel & s820) | (sub_sel & sub820) | (and_sel & and820) | (or_sel & or820);
  assign y821 = (add_sel & s821) | (sub_sel & sub821) | (and_sel & and821) | (or_sel & or821);
  assign y822 = (add_sel & s822) | (sub_sel & sub822) | (and_sel & and822) | (or_sel & or822);
  assign y823 = (add_sel & s823) | (sub_sel & sub823) | (and_sel & and823) | (or_sel & or823);
  assign y824 = (add_sel & s824) | (sub_sel & sub824) | (and_sel & and824) | (or_sel & or824);
  assign y825 = (add_sel & s825) | (sub_sel & sub825) | (and_sel & and825) | (or_sel & or825);
  assign y826 = (add_sel & s826) | (sub_sel & sub826) | (and_sel & and826) | (or_sel & or826);
  assign y827 = (add_sel & s827) | (sub_sel & sub827) | (and_sel & and827) | (or_sel & or827);
  assign y828 = (add_sel & s828) | (sub_sel & sub828) | (and_sel & and828) | (or_sel & or828);
  assign y829 = (add_sel & s829) | (sub_sel & sub829) | (and_sel & and829) | (or_sel & or829);
  assign y830 = (add_sel & s830) | (sub_sel & sub830) | (and_sel & and830) | (or_sel & or830);
  assign y831 = (add_sel & s831) | (sub_sel & sub831) | (and_sel & and831) | (or_sel & or831);
  assign y832 = (add_sel & s832) | (sub_sel & sub832) | (and_sel & and832) | (or_sel & or832);
  assign y833 = (add_sel & s833) | (sub_sel & sub833) | (and_sel & and833) | (or_sel & or833);
  assign y834 = (add_sel & s834) | (sub_sel & sub834) | (and_sel & and834) | (or_sel & or834);
  assign y835 = (add_sel & s835) | (sub_sel & sub835) | (and_sel & and835) | (or_sel & or835);
  assign y836 = (add_sel & s836) | (sub_sel & sub836) | (and_sel & and836) | (or_sel & or836);
  assign y837 = (add_sel & s837) | (sub_sel & sub837) | (and_sel & and837) | (or_sel & or837);
  assign y838 = (add_sel & s838) | (sub_sel & sub838) | (and_sel & and838) | (or_sel & or838);
  assign y839 = (add_sel & s839) | (sub_sel & sub839) | (and_sel & and839) | (or_sel & or839);
  assign y840 = (add_sel & s840) | (sub_sel & sub840) | (and_sel & and840) | (or_sel & or840);
  assign y841 = (add_sel & s841) | (sub_sel & sub841) | (and_sel & and841) | (or_sel & or841);
  assign y842 = (add_sel & s842) | (sub_sel & sub842) | (and_sel & and842) | (or_sel & or842);
  assign y843 = (add_sel & s843) | (sub_sel & sub843) | (and_sel & and843) | (or_sel & or843);
  assign y844 = (add_sel & s844) | (sub_sel & sub844) | (and_sel & and844) | (or_sel & or844);
  assign y845 = (add_sel & s845) | (sub_sel & sub845) | (and_sel & and845) | (or_sel & or845);
  assign y846 = (add_sel & s846) | (sub_sel & sub846) | (and_sel & and846) | (or_sel & or846);
  assign y847 = (add_sel & s847) | (sub_sel & sub847) | (and_sel & and847) | (or_sel & or847);
  assign y848 = (add_sel & s848) | (sub_sel & sub848) | (and_sel & and848) | (or_sel & or848);
  assign y849 = (add_sel & s849) | (sub_sel & sub849) | (and_sel & and849) | (or_sel & or849);
  assign y850 = (add_sel & s850) | (sub_sel & sub850) | (and_sel & and850) | (or_sel & or850);
  assign y851 = (add_sel & s851) | (sub_sel & sub851) | (and_sel & and851) | (or_sel & or851);
  assign y852 = (add_sel & s852) | (sub_sel & sub852) | (and_sel & and852) | (or_sel & or852);
  assign y853 = (add_sel & s853) | (sub_sel & sub853) | (and_sel & and853) | (or_sel & or853);
  assign y854 = (add_sel & s854) | (sub_sel & sub854) | (and_sel & and854) | (or_sel & or854);
  assign y855 = (add_sel & s855) | (sub_sel & sub855) | (and_sel & and855) | (or_sel & or855);
  assign y856 = (add_sel & s856) | (sub_sel & sub856) | (and_sel & and856) | (or_sel & or856);
  assign y857 = (add_sel & s857) | (sub_sel & sub857) | (and_sel & and857) | (or_sel & or857);
  assign y858 = (add_sel & s858) | (sub_sel & sub858) | (and_sel & and858) | (or_sel & or858);
  assign y859 = (add_sel & s859) | (sub_sel & sub859) | (and_sel & and859) | (or_sel & or859);
  assign y860 = (add_sel & s860) | (sub_sel & sub860) | (and_sel & and860) | (or_sel & or860);
  assign y861 = (add_sel & s861) | (sub_sel & sub861) | (and_sel & and861) | (or_sel & or861);
  assign y862 = (add_sel & s862) | (sub_sel & sub862) | (and_sel & and862) | (or_sel & or862);
  assign y863 = (add_sel & s863) | (sub_sel & sub863) | (and_sel & and863) | (or_sel & or863);
  assign y864 = (add_sel & s864) | (sub_sel & sub864) | (and_sel & and864) | (or_sel & or864);
  assign y865 = (add_sel & s865) | (sub_sel & sub865) | (and_sel & and865) | (or_sel & or865);
  assign y866 = (add_sel & s866) | (sub_sel & sub866) | (and_sel & and866) | (or_sel & or866);
  assign y867 = (add_sel & s867) | (sub_sel & sub867) | (and_sel & and867) | (or_sel & or867);
  assign y868 = (add_sel & s868) | (sub_sel & sub868) | (and_sel & and868) | (or_sel & or868);
  assign y869 = (add_sel & s869) | (sub_sel & sub869) | (and_sel & and869) | (or_sel & or869);
  assign y870 = (add_sel & s870) | (sub_sel & sub870) | (and_sel & and870) | (or_sel & or870);
  assign y871 = (add_sel & s871) | (sub_sel & sub871) | (and_sel & and871) | (or_sel & or871);
  assign y872 = (add_sel & s872) | (sub_sel & sub872) | (and_sel & and872) | (or_sel & or872);
  assign y873 = (add_sel & s873) | (sub_sel & sub873) | (and_sel & and873) | (or_sel & or873);
  assign y874 = (add_sel & s874) | (sub_sel & sub874) | (and_sel & and874) | (or_sel & or874);
  assign y875 = (add_sel & s875) | (sub_sel & sub875) | (and_sel & and875) | (or_sel & or875);
  assign y876 = (add_sel & s876) | (sub_sel & sub876) | (and_sel & and876) | (or_sel & or876);
  assign y877 = (add_sel & s877) | (sub_sel & sub877) | (and_sel & and877) | (or_sel & or877);
  assign y878 = (add_sel & s878) | (sub_sel & sub878) | (and_sel & and878) | (or_sel & or878);
  assign y879 = (add_sel & s879) | (sub_sel & sub879) | (and_sel & and879) | (or_sel & or879);
  assign y880 = (add_sel & s880) | (sub_sel & sub880) | (and_sel & and880) | (or_sel & or880);
  assign y881 = (add_sel & s881) | (sub_sel & sub881) | (and_sel & and881) | (or_sel & or881);
  assign y882 = (add_sel & s882) | (sub_sel & sub882) | (and_sel & and882) | (or_sel & or882);
  assign y883 = (add_sel & s883) | (sub_sel & sub883) | (and_sel & and883) | (or_sel & or883);
  assign y884 = (add_sel & s884) | (sub_sel & sub884) | (and_sel & and884) | (or_sel & or884);
  assign y885 = (add_sel & s885) | (sub_sel & sub885) | (and_sel & and885) | (or_sel & or885);
  assign y886 = (add_sel & s886) | (sub_sel & sub886) | (and_sel & and886) | (or_sel & or886);
  assign y887 = (add_sel & s887) | (sub_sel & sub887) | (and_sel & and887) | (or_sel & or887);
  assign y888 = (add_sel & s888) | (sub_sel & sub888) | (and_sel & and888) | (or_sel & or888);
  assign y889 = (add_sel & s889) | (sub_sel & sub889) | (and_sel & and889) | (or_sel & or889);
  assign y890 = (add_sel & s890) | (sub_sel & sub890) | (and_sel & and890) | (or_sel & or890);
  assign y891 = (add_sel & s891) | (sub_sel & sub891) | (and_sel & and891) | (or_sel & or891);
  assign y892 = (add_sel & s892) | (sub_sel & sub892) | (and_sel & and892) | (or_sel & or892);
  assign y893 = (add_sel & s893) | (sub_sel & sub893) | (and_sel & and893) | (or_sel & or893);
  assign y894 = (add_sel & s894) | (sub_sel & sub894) | (and_sel & and894) | (or_sel & or894);
  assign y895 = (add_sel & s895) | (sub_sel & sub895) | (and_sel & and895) | (or_sel & or895);
  assign y896 = (add_sel & s896) | (sub_sel & sub896) | (and_sel & and896) | (or_sel & or896);
  assign y897 = (add_sel & s897) | (sub_sel & sub897) | (and_sel & and897) | (or_sel & or897);
  assign y898 = (add_sel & s898) | (sub_sel & sub898) | (and_sel & and898) | (or_sel & or898);
  assign y899 = (add_sel & s899) | (sub_sel & sub899) | (and_sel & and899) | (or_sel & or899);
  assign y900 = (add_sel & s900) | (sub_sel & sub900) | (and_sel & and900) | (or_sel & or900);
  assign y901 = (add_sel & s901) | (sub_sel & sub901) | (and_sel & and901) | (or_sel & or901);
  assign y902 = (add_sel & s902) | (sub_sel & sub902) | (and_sel & and902) | (or_sel & or902);
  assign y903 = (add_sel & s903) | (sub_sel & sub903) | (and_sel & and903) | (or_sel & or903);
  assign y904 = (add_sel & s904) | (sub_sel & sub904) | (and_sel & and904) | (or_sel & or904);
  assign y905 = (add_sel & s905) | (sub_sel & sub905) | (and_sel & and905) | (or_sel & or905);
  assign y906 = (add_sel & s906) | (sub_sel & sub906) | (and_sel & and906) | (or_sel & or906);
  assign y907 = (add_sel & s907) | (sub_sel & sub907) | (and_sel & and907) | (or_sel & or907);
  assign y908 = (add_sel & s908) | (sub_sel & sub908) | (and_sel & and908) | (or_sel & or908);
  assign y909 = (add_sel & s909) | (sub_sel & sub909) | (and_sel & and909) | (or_sel & or909);
  assign y910 = (add_sel & s910) | (sub_sel & sub910) | (and_sel & and910) | (or_sel & or910);
  assign y911 = (add_sel & s911) | (sub_sel & sub911) | (and_sel & and911) | (or_sel & or911);
  assign y912 = (add_sel & s912) | (sub_sel & sub912) | (and_sel & and912) | (or_sel & or912);
  assign y913 = (add_sel & s913) | (sub_sel & sub913) | (and_sel & and913) | (or_sel & or913);
  assign y914 = (add_sel & s914) | (sub_sel & sub914) | (and_sel & and914) | (or_sel & or914);
  assign y915 = (add_sel & s915) | (sub_sel & sub915) | (and_sel & and915) | (or_sel & or915);
  assign y916 = (add_sel & s916) | (sub_sel & sub916) | (and_sel & and916) | (or_sel & or916);
  assign y917 = (add_sel & s917) | (sub_sel & sub917) | (and_sel & and917) | (or_sel & or917);
  assign y918 = (add_sel & s918) | (sub_sel & sub918) | (and_sel & and918) | (or_sel & or918);
  assign y919 = (add_sel & s919) | (sub_sel & sub919) | (and_sel & and919) | (or_sel & or919);
  assign y920 = (add_sel & s920) | (sub_sel & sub920) | (and_sel & and920) | (or_sel & or920);
  assign y921 = (add_sel & s921) | (sub_sel & sub921) | (and_sel & and921) | (or_sel & or921);
  assign y922 = (add_sel & s922) | (sub_sel & sub922) | (and_sel & and922) | (or_sel & or922);
  assign y923 = (add_sel & s923) | (sub_sel & sub923) | (and_sel & and923) | (or_sel & or923);
  assign y924 = (add_sel & s924) | (sub_sel & sub924) | (and_sel & and924) | (or_sel & or924);
  assign y925 = (add_sel & s925) | (sub_sel & sub925) | (and_sel & and925) | (or_sel & or925);
  assign y926 = (add_sel & s926) | (sub_sel & sub926) | (and_sel & and926) | (or_sel & or926);
  assign y927 = (add_sel & s927) | (sub_sel & sub927) | (and_sel & and927) | (or_sel & or927);
  assign y928 = (add_sel & s928) | (sub_sel & sub928) | (and_sel & and928) | (or_sel & or928);
  assign y929 = (add_sel & s929) | (sub_sel & sub929) | (and_sel & and929) | (or_sel & or929);
  assign y930 = (add_sel & s930) | (sub_sel & sub930) | (and_sel & and930) | (or_sel & or930);
  assign y931 = (add_sel & s931) | (sub_sel & sub931) | (and_sel & and931) | (or_sel & or931);
  assign y932 = (add_sel & s932) | (sub_sel & sub932) | (and_sel & and932) | (or_sel & or932);
  assign y933 = (add_sel & s933) | (sub_sel & sub933) | (and_sel & and933) | (or_sel & or933);
  assign y934 = (add_sel & s934) | (sub_sel & sub934) | (and_sel & and934) | (or_sel & or934);
  assign y935 = (add_sel & s935) | (sub_sel & sub935) | (and_sel & and935) | (or_sel & or935);
  assign y936 = (add_sel & s936) | (sub_sel & sub936) | (and_sel & and936) | (or_sel & or936);
  assign y937 = (add_sel & s937) | (sub_sel & sub937) | (and_sel & and937) | (or_sel & or937);
  assign y938 = (add_sel & s938) | (sub_sel & sub938) | (and_sel & and938) | (or_sel & or938);
  assign y939 = (add_sel & s939) | (sub_sel & sub939) | (and_sel & and939) | (or_sel & or939);
  assign y940 = (add_sel & s940) | (sub_sel & sub940) | (and_sel & and940) | (or_sel & or940);
  assign y941 = (add_sel & s941) | (sub_sel & sub941) | (and_sel & and941) | (or_sel & or941);
  assign y942 = (add_sel & s942) | (sub_sel & sub942) | (and_sel & and942) | (or_sel & or942);
  assign y943 = (add_sel & s943) | (sub_sel & sub943) | (and_sel & and943) | (or_sel & or943);
  assign y944 = (add_sel & s944) | (sub_sel & sub944) | (and_sel & and944) | (or_sel & or944);
  assign y945 = (add_sel & s945) | (sub_sel & sub945) | (and_sel & and945) | (or_sel & or945);
  assign y946 = (add_sel & s946) | (sub_sel & sub946) | (and_sel & and946) | (or_sel & or946);
  assign y947 = (add_sel & s947) | (sub_sel & sub947) | (and_sel & and947) | (or_sel & or947);
  assign y948 = (add_sel & s948) | (sub_sel & sub948) | (and_sel & and948) | (or_sel & or948);
  assign y949 = (add_sel & s949) | (sub_sel & sub949) | (and_sel & and949) | (or_sel & or949);
  assign y950 = (add_sel & s950) | (sub_sel & sub950) | (and_sel & and950) | (or_sel & or950);
  assign y951 = (add_sel & s951) | (sub_sel & sub951) | (and_sel & and951) | (or_sel & or951);
  assign y952 = (add_sel & s952) | (sub_sel & sub952) | (and_sel & and952) | (or_sel & or952);
  assign y953 = (add_sel & s953) | (sub_sel & sub953) | (and_sel & and953) | (or_sel & or953);
  assign y954 = (add_sel & s954) | (sub_sel & sub954) | (and_sel & and954) | (or_sel & or954);
  assign y955 = (add_sel & s955) | (sub_sel & sub955) | (and_sel & and955) | (or_sel & or955);
  assign y956 = (add_sel & s956) | (sub_sel & sub956) | (and_sel & and956) | (or_sel & or956);
  assign y957 = (add_sel & s957) | (sub_sel & sub957) | (and_sel & and957) | (or_sel & or957);
  assign y958 = (add_sel & s958) | (sub_sel & sub958) | (and_sel & and958) | (or_sel & or958);
  assign y959 = (add_sel & s959) | (sub_sel & sub959) | (and_sel & and959) | (or_sel & or959);
  assign y960 = (add_sel & s960) | (sub_sel & sub960) | (and_sel & and960) | (or_sel & or960);
  assign y961 = (add_sel & s961) | (sub_sel & sub961) | (and_sel & and961) | (or_sel & or961);
  assign y962 = (add_sel & s962) | (sub_sel & sub962) | (and_sel & and962) | (or_sel & or962);
  assign y963 = (add_sel & s963) | (sub_sel & sub963) | (and_sel & and963) | (or_sel & or963);
  assign y964 = (add_sel & s964) | (sub_sel & sub964) | (and_sel & and964) | (or_sel & or964);
  assign y965 = (add_sel & s965) | (sub_sel & sub965) | (and_sel & and965) | (or_sel & or965);
  assign y966 = (add_sel & s966) | (sub_sel & sub966) | (and_sel & and966) | (or_sel & or966);
  assign y967 = (add_sel & s967) | (sub_sel & sub967) | (and_sel & and967) | (or_sel & or967);
  assign y968 = (add_sel & s968) | (sub_sel & sub968) | (and_sel & and968) | (or_sel & or968);
  assign y969 = (add_sel & s969) | (sub_sel & sub969) | (and_sel & and969) | (or_sel & or969);
  assign y970 = (add_sel & s970) | (sub_sel & sub970) | (and_sel & and970) | (or_sel & or970);
  assign y971 = (add_sel & s971) | (sub_sel & sub971) | (and_sel & and971) | (or_sel & or971);
  assign y972 = (add_sel & s972) | (sub_sel & sub972) | (and_sel & and972) | (or_sel & or972);
  assign y973 = (add_sel & s973) | (sub_sel & sub973) | (and_sel & and973) | (or_sel & or973);
  assign y974 = (add_sel & s974) | (sub_sel & sub974) | (and_sel & and974) | (or_sel & or974);
  assign y975 = (add_sel & s975) | (sub_sel & sub975) | (and_sel & and975) | (or_sel & or975);
  assign y976 = (add_sel & s976) | (sub_sel & sub976) | (and_sel & and976) | (or_sel & or976);
  assign y977 = (add_sel & s977) | (sub_sel & sub977) | (and_sel & and977) | (or_sel & or977);
  assign y978 = (add_sel & s978) | (sub_sel & sub978) | (and_sel & and978) | (or_sel & or978);
  assign y979 = (add_sel & s979) | (sub_sel & sub979) | (and_sel & and979) | (or_sel & or979);
  assign y980 = (add_sel & s980) | (sub_sel & sub980) | (and_sel & and980) | (or_sel & or980);
  assign y981 = (add_sel & s981) | (sub_sel & sub981) | (and_sel & and981) | (or_sel & or981);
  assign y982 = (add_sel & s982) | (sub_sel & sub982) | (and_sel & and982) | (or_sel & or982);
  assign y983 = (add_sel & s983) | (sub_sel & sub983) | (and_sel & and983) | (or_sel & or983);
  assign y984 = (add_sel & s984) | (sub_sel & sub984) | (and_sel & and984) | (or_sel & or984);
  assign y985 = (add_sel & s985) | (sub_sel & sub985) | (and_sel & and985) | (or_sel & or985);
  assign y986 = (add_sel & s986) | (sub_sel & sub986) | (and_sel & and986) | (or_sel & or986);
  assign y987 = (add_sel & s987) | (sub_sel & sub987) | (and_sel & and987) | (or_sel & or987);
  assign y988 = (add_sel & s988) | (sub_sel & sub988) | (and_sel & and988) | (or_sel & or988);
  assign y989 = (add_sel & s989) | (sub_sel & sub989) | (and_sel & and989) | (or_sel & or989);
  assign y990 = (add_sel & s990) | (sub_sel & sub990) | (and_sel & and990) | (or_sel & or990);
  assign y991 = (add_sel & s991) | (sub_sel & sub991) | (and_sel & and991) | (or_sel & or991);
  assign y992 = (add_sel & s992) | (sub_sel & sub992) | (and_sel & and992) | (or_sel & or992);
  assign y993 = (add_sel & s993) | (sub_sel & sub993) | (and_sel & and993) | (or_sel & or993);
  assign y994 = (add_sel & s994) | (sub_sel & sub994) | (and_sel & and994) | (or_sel & or994);
  assign y995 = (add_sel & s995) | (sub_sel & sub995) | (and_sel & and995) | (or_sel & or995);
  assign y996 = (add_sel & s996) | (sub_sel & sub996) | (and_sel & and996) | (or_sel & or996);
  assign y997 = (add_sel & s997) | (sub_sel & sub997) | (and_sel & and997) | (or_sel & or997);
  assign y998 = (add_sel & s998) | (sub_sel & sub998) | (and_sel & and998) | (or_sel & or998);
  assign y999 = (add_sel & s999) | (sub_sel & sub999) | (and_sel & and999) | (or_sel & or999);
  assign y1000 = (add_sel & s1000) | (sub_sel & sub1000) | (and_sel & and1000) | (or_sel & or1000);
  assign y1001 = (add_sel & s1001) | (sub_sel & sub1001) | (and_sel & and1001) | (or_sel & or1001);
  assign y1002 = (add_sel & s1002) | (sub_sel & sub1002) | (and_sel & and1002) | (or_sel & or1002);
  assign y1003 = (add_sel & s1003) | (sub_sel & sub1003) | (and_sel & and1003) | (or_sel & or1003);
  assign y1004 = (add_sel & s1004) | (sub_sel & sub1004) | (and_sel & and1004) | (or_sel & or1004);
  assign y1005 = (add_sel & s1005) | (sub_sel & sub1005) | (and_sel & and1005) | (or_sel & or1005);
  assign y1006 = (add_sel & s1006) | (sub_sel & sub1006) | (and_sel & and1006) | (or_sel & or1006);
  assign y1007 = (add_sel & s1007) | (sub_sel & sub1007) | (and_sel & and1007) | (or_sel & or1007);
  assign y1008 = (add_sel & s1008) | (sub_sel & sub1008) | (and_sel & and1008) | (or_sel & or1008);
  assign y1009 = (add_sel & s1009) | (sub_sel & sub1009) | (and_sel & and1009) | (or_sel & or1009);
  assign y1010 = (add_sel & s1010) | (sub_sel & sub1010) | (and_sel & and1010) | (or_sel & or1010);
  assign y1011 = (add_sel & s1011) | (sub_sel & sub1011) | (and_sel & and1011) | (or_sel & or1011);
  assign y1012 = (add_sel & s1012) | (sub_sel & sub1012) | (and_sel & and1012) | (or_sel & or1012);
  assign y1013 = (add_sel & s1013) | (sub_sel & sub1013) | (and_sel & and1013) | (or_sel & or1013);
  assign y1014 = (add_sel & s1014) | (sub_sel & sub1014) | (and_sel & and1014) | (or_sel & or1014);
  assign y1015 = (add_sel & s1015) | (sub_sel & sub1015) | (and_sel & and1015) | (or_sel & or1015);
  assign y1016 = (add_sel & s1016) | (sub_sel & sub1016) | (and_sel & and1016) | (or_sel & or1016);
  assign y1017 = (add_sel & s1017) | (sub_sel & sub1017) | (and_sel & and1017) | (or_sel & or1017);
  assign y1018 = (add_sel & s1018) | (sub_sel & sub1018) | (and_sel & and1018) | (or_sel & or1018);
  assign y1019 = (add_sel & s1019) | (sub_sel & sub1019) | (and_sel & and1019) | (or_sel & or1019);
  assign y1020 = (add_sel & s1020) | (sub_sel & sub1020) | (and_sel & and1020) | (or_sel & or1020);
  assign y1021 = (add_sel & s1021) | (sub_sel & sub1021) | (and_sel & and1021) | (or_sel & or1021);
  assign y1022 = (add_sel & s1022) | (sub_sel & sub1022) | (and_sel & and1022) | (or_sel & or1022);
  assign y1023 = (add_sel & s1023) | (sub_sel & sub1023) | (and_sel & and1023) | (or_sel & or1023);
  assign y1024 = (add_sel & s1024) | (sub_sel & sub1024) | (and_sel & and1024) | (or_sel & or1024);
  assign y1025 = (add_sel & s1025) | (sub_sel & sub1025) | (and_sel & and1025) | (or_sel & or1025);
  assign y1026 = (add_sel & s1026) | (sub_sel & sub1026) | (and_sel & and1026) | (or_sel & or1026);
  assign y1027 = (add_sel & s1027) | (sub_sel & sub1027) | (and_sel & and1027) | (or_sel & or1027);
  assign y1028 = (add_sel & s1028) | (sub_sel & sub1028) | (and_sel & and1028) | (or_sel & or1028);
  assign y1029 = (add_sel & s1029) | (sub_sel & sub1029) | (and_sel & and1029) | (or_sel & or1029);
  assign y1030 = (add_sel & s1030) | (sub_sel & sub1030) | (and_sel & and1030) | (or_sel & or1030);
  assign y1031 = (add_sel & s1031) | (sub_sel & sub1031) | (and_sel & and1031) | (or_sel & or1031);
  assign y1032 = (add_sel & s1032) | (sub_sel & sub1032) | (and_sel & and1032) | (or_sel & or1032);
  assign y1033 = (add_sel & s1033) | (sub_sel & sub1033) | (and_sel & and1033) | (or_sel & or1033);
  assign y1034 = (add_sel & s1034) | (sub_sel & sub1034) | (and_sel & and1034) | (or_sel & or1034);
  assign y1035 = (add_sel & s1035) | (sub_sel & sub1035) | (and_sel & and1035) | (or_sel & or1035);
  assign y1036 = (add_sel & s1036) | (sub_sel & sub1036) | (and_sel & and1036) | (or_sel & or1036);
  assign y1037 = (add_sel & s1037) | (sub_sel & sub1037) | (and_sel & and1037) | (or_sel & or1037);
  assign y1038 = (add_sel & s1038) | (sub_sel & sub1038) | (and_sel & and1038) | (or_sel & or1038);
  assign y1039 = (add_sel & s1039) | (sub_sel & sub1039) | (and_sel & and1039) | (or_sel & or1039);
  assign y1040 = (add_sel & s1040) | (sub_sel & sub1040) | (and_sel & and1040) | (or_sel & or1040);
  assign y1041 = (add_sel & s1041) | (sub_sel & sub1041) | (and_sel & and1041) | (or_sel & or1041);
  assign y1042 = (add_sel & s1042) | (sub_sel & sub1042) | (and_sel & and1042) | (or_sel & or1042);
  assign y1043 = (add_sel & s1043) | (sub_sel & sub1043) | (and_sel & and1043) | (or_sel & or1043);
  assign y1044 = (add_sel & s1044) | (sub_sel & sub1044) | (and_sel & and1044) | (or_sel & or1044);
  assign y1045 = (add_sel & s1045) | (sub_sel & sub1045) | (and_sel & and1045) | (or_sel & or1045);
  assign y1046 = (add_sel & s1046) | (sub_sel & sub1046) | (and_sel & and1046) | (or_sel & or1046);
  assign y1047 = (add_sel & s1047) | (sub_sel & sub1047) | (and_sel & and1047) | (or_sel & or1047);
  assign y1048 = (add_sel & s1048) | (sub_sel & sub1048) | (and_sel & and1048) | (or_sel & or1048);
  assign y1049 = (add_sel & s1049) | (sub_sel & sub1049) | (and_sel & and1049) | (or_sel & or1049);
  assign y1050 = (add_sel & s1050) | (sub_sel & sub1050) | (and_sel & and1050) | (or_sel & or1050);
  assign y1051 = (add_sel & s1051) | (sub_sel & sub1051) | (and_sel & and1051) | (or_sel & or1051);
  assign y1052 = (add_sel & s1052) | (sub_sel & sub1052) | (and_sel & and1052) | (or_sel & or1052);
  assign y1053 = (add_sel & s1053) | (sub_sel & sub1053) | (and_sel & and1053) | (or_sel & or1053);
  assign y1054 = (add_sel & s1054) | (sub_sel & sub1054) | (and_sel & and1054) | (or_sel & or1054);
  assign y1055 = (add_sel & s1055) | (sub_sel & sub1055) | (and_sel & and1055) | (or_sel & or1055);
  assign y1056 = (add_sel & s1056) | (sub_sel & sub1056) | (and_sel & and1056) | (or_sel & or1056);
  assign y1057 = (add_sel & s1057) | (sub_sel & sub1057) | (and_sel & and1057) | (or_sel & or1057);
  assign y1058 = (add_sel & s1058) | (sub_sel & sub1058) | (and_sel & and1058) | (or_sel & or1058);
  assign y1059 = (add_sel & s1059) | (sub_sel & sub1059) | (and_sel & and1059) | (or_sel & or1059);
  assign y1060 = (add_sel & s1060) | (sub_sel & sub1060) | (and_sel & and1060) | (or_sel & or1060);
  assign y1061 = (add_sel & s1061) | (sub_sel & sub1061) | (and_sel & and1061) | (or_sel & or1061);
  assign y1062 = (add_sel & s1062) | (sub_sel & sub1062) | (and_sel & and1062) | (or_sel & or1062);
  assign y1063 = (add_sel & s1063) | (sub_sel & sub1063) | (and_sel & and1063) | (or_sel & or1063);
  assign y1064 = (add_sel & s1064) | (sub_sel & sub1064) | (and_sel & and1064) | (or_sel & or1064);
  assign y1065 = (add_sel & s1065) | (sub_sel & sub1065) | (and_sel & and1065) | (or_sel & or1065);
  assign y1066 = (add_sel & s1066) | (sub_sel & sub1066) | (and_sel & and1066) | (or_sel & or1066);
  assign y1067 = (add_sel & s1067) | (sub_sel & sub1067) | (and_sel & and1067) | (or_sel & or1067);
  assign y1068 = (add_sel & s1068) | (sub_sel & sub1068) | (and_sel & and1068) | (or_sel & or1068);
  assign y1069 = (add_sel & s1069) | (sub_sel & sub1069) | (and_sel & and1069) | (or_sel & or1069);
  assign y1070 = (add_sel & s1070) | (sub_sel & sub1070) | (and_sel & and1070) | (or_sel & or1070);
  assign y1071 = (add_sel & s1071) | (sub_sel & sub1071) | (and_sel & and1071) | (or_sel & or1071);
  assign y1072 = (add_sel & s1072) | (sub_sel & sub1072) | (and_sel & and1072) | (or_sel & or1072);
  assign y1073 = (add_sel & s1073) | (sub_sel & sub1073) | (and_sel & and1073) | (or_sel & or1073);
  assign y1074 = (add_sel & s1074) | (sub_sel & sub1074) | (and_sel & and1074) | (or_sel & or1074);
  assign y1075 = (add_sel & s1075) | (sub_sel & sub1075) | (and_sel & and1075) | (or_sel & or1075);
  assign y1076 = (add_sel & s1076) | (sub_sel & sub1076) | (and_sel & and1076) | (or_sel & or1076);
  assign y1077 = (add_sel & s1077) | (sub_sel & sub1077) | (and_sel & and1077) | (or_sel & or1077);
  assign y1078 = (add_sel & s1078) | (sub_sel & sub1078) | (and_sel & and1078) | (or_sel & or1078);
  assign y1079 = (add_sel & s1079) | (sub_sel & sub1079) | (and_sel & and1079) | (or_sel & or1079);
  assign y1080 = (add_sel & s1080) | (sub_sel & sub1080) | (and_sel & and1080) | (or_sel & or1080);
  assign y1081 = (add_sel & s1081) | (sub_sel & sub1081) | (and_sel & and1081) | (or_sel & or1081);
  assign y1082 = (add_sel & s1082) | (sub_sel & sub1082) | (and_sel & and1082) | (or_sel & or1082);
  assign y1083 = (add_sel & s1083) | (sub_sel & sub1083) | (and_sel & and1083) | (or_sel & or1083);
  assign y1084 = (add_sel & s1084) | (sub_sel & sub1084) | (and_sel & and1084) | (or_sel & or1084);
  assign y1085 = (add_sel & s1085) | (sub_sel & sub1085) | (and_sel & and1085) | (or_sel & or1085);
  assign y1086 = (add_sel & s1086) | (sub_sel & sub1086) | (and_sel & and1086) | (or_sel & or1086);
  assign y1087 = (add_sel & s1087) | (sub_sel & sub1087) | (and_sel & and1087) | (or_sel & or1087);
  assign y1088 = (add_sel & s1088) | (sub_sel & sub1088) | (and_sel & and1088) | (or_sel & or1088);
  assign y1089 = (add_sel & s1089) | (sub_sel & sub1089) | (and_sel & and1089) | (or_sel & or1089);
  assign y1090 = (add_sel & s1090) | (sub_sel & sub1090) | (and_sel & and1090) | (or_sel & or1090);
  assign y1091 = (add_sel & s1091) | (sub_sel & sub1091) | (and_sel & and1091) | (or_sel & or1091);
  assign y1092 = (add_sel & s1092) | (sub_sel & sub1092) | (and_sel & and1092) | (or_sel & or1092);
  assign y1093 = (add_sel & s1093) | (sub_sel & sub1093) | (and_sel & and1093) | (or_sel & or1093);
  assign y1094 = (add_sel & s1094) | (sub_sel & sub1094) | (and_sel & and1094) | (or_sel & or1094);
  assign y1095 = (add_sel & s1095) | (sub_sel & sub1095) | (and_sel & and1095) | (or_sel & or1095);
  assign y1096 = (add_sel & s1096) | (sub_sel & sub1096) | (and_sel & and1096) | (or_sel & or1096);
  assign y1097 = (add_sel & s1097) | (sub_sel & sub1097) | (and_sel & and1097) | (or_sel & or1097);
  assign y1098 = (add_sel & s1098) | (sub_sel & sub1098) | (and_sel & and1098) | (or_sel & or1098);
  assign y1099 = (add_sel & s1099) | (sub_sel & sub1099) | (and_sel & and1099) | (or_sel & or1099);
  assign y1100 = (add_sel & s1100) | (sub_sel & sub1100) | (and_sel & and1100) | (or_sel & or1100);
  assign y1101 = (add_sel & s1101) | (sub_sel & sub1101) | (and_sel & and1101) | (or_sel & or1101);
  assign y1102 = (add_sel & s1102) | (sub_sel & sub1102) | (and_sel & and1102) | (or_sel & or1102);
  assign y1103 = (add_sel & s1103) | (sub_sel & sub1103) | (and_sel & and1103) | (or_sel & or1103);
  assign y1104 = (add_sel & s1104) | (sub_sel & sub1104) | (and_sel & and1104) | (or_sel & or1104);
  assign y1105 = (add_sel & s1105) | (sub_sel & sub1105) | (and_sel & and1105) | (or_sel & or1105);
  assign y1106 = (add_sel & s1106) | (sub_sel & sub1106) | (and_sel & and1106) | (or_sel & or1106);
  assign y1107 = (add_sel & s1107) | (sub_sel & sub1107) | (and_sel & and1107) | (or_sel & or1107);
  assign y1108 = (add_sel & s1108) | (sub_sel & sub1108) | (and_sel & and1108) | (or_sel & or1108);
  assign y1109 = (add_sel & s1109) | (sub_sel & sub1109) | (and_sel & and1109) | (or_sel & or1109);
  assign y1110 = (add_sel & s1110) | (sub_sel & sub1110) | (and_sel & and1110) | (or_sel & or1110);
  assign y1111 = (add_sel & s1111) | (sub_sel & sub1111) | (and_sel & and1111) | (or_sel & or1111);
  assign y1112 = (add_sel & s1112) | (sub_sel & sub1112) | (and_sel & and1112) | (or_sel & or1112);
  assign y1113 = (add_sel & s1113) | (sub_sel & sub1113) | (and_sel & and1113) | (or_sel & or1113);
  assign y1114 = (add_sel & s1114) | (sub_sel & sub1114) | (and_sel & and1114) | (or_sel & or1114);
  assign y1115 = (add_sel & s1115) | (sub_sel & sub1115) | (and_sel & and1115) | (or_sel & or1115);
  assign y1116 = (add_sel & s1116) | (sub_sel & sub1116) | (and_sel & and1116) | (or_sel & or1116);
  assign y1117 = (add_sel & s1117) | (sub_sel & sub1117) | (and_sel & and1117) | (or_sel & or1117);
  assign y1118 = (add_sel & s1118) | (sub_sel & sub1118) | (and_sel & and1118) | (or_sel & or1118);
  assign y1119 = (add_sel & s1119) | (sub_sel & sub1119) | (and_sel & and1119) | (or_sel & or1119);
  assign y1120 = (add_sel & s1120) | (sub_sel & sub1120) | (and_sel & and1120) | (or_sel & or1120);
  assign y1121 = (add_sel & s1121) | (sub_sel & sub1121) | (and_sel & and1121) | (or_sel & or1121);
  assign y1122 = (add_sel & s1122) | (sub_sel & sub1122) | (and_sel & and1122) | (or_sel & or1122);
  assign y1123 = (add_sel & s1123) | (sub_sel & sub1123) | (and_sel & and1123) | (or_sel & or1123);
  assign y1124 = (add_sel & s1124) | (sub_sel & sub1124) | (and_sel & and1124) | (or_sel & or1124);
  assign y1125 = (add_sel & s1125) | (sub_sel & sub1125) | (and_sel & and1125) | (or_sel & or1125);
  assign y1126 = (add_sel & s1126) | (sub_sel & sub1126) | (and_sel & and1126) | (or_sel & or1126);
  assign y1127 = (add_sel & s1127) | (sub_sel & sub1127) | (and_sel & and1127) | (or_sel & or1127);
  assign y1128 = (add_sel & s1128) | (sub_sel & sub1128) | (and_sel & and1128) | (or_sel & or1128);
  assign y1129 = (add_sel & s1129) | (sub_sel & sub1129) | (and_sel & and1129) | (or_sel & or1129);
  assign y1130 = (add_sel & s1130) | (sub_sel & sub1130) | (and_sel & and1130) | (or_sel & or1130);
  assign y1131 = (add_sel & s1131) | (sub_sel & sub1131) | (and_sel & and1131) | (or_sel & or1131);
  assign y1132 = (add_sel & s1132) | (sub_sel & sub1132) | (and_sel & and1132) | (or_sel & or1132);
  assign y1133 = (add_sel & s1133) | (sub_sel & sub1133) | (and_sel & and1133) | (or_sel & or1133);
  assign y1134 = (add_sel & s1134) | (sub_sel & sub1134) | (and_sel & and1134) | (or_sel & or1134);
  assign y1135 = (add_sel & s1135) | (sub_sel & sub1135) | (and_sel & and1135) | (or_sel & or1135);
  assign y1136 = (add_sel & s1136) | (sub_sel & sub1136) | (and_sel & and1136) | (or_sel & or1136);
  assign y1137 = (add_sel & s1137) | (sub_sel & sub1137) | (and_sel & and1137) | (or_sel & or1137);
  assign y1138 = (add_sel & s1138) | (sub_sel & sub1138) | (and_sel & and1138) | (or_sel & or1138);
  assign y1139 = (add_sel & s1139) | (sub_sel & sub1139) | (and_sel & and1139) | (or_sel & or1139);
  assign y1140 = (add_sel & s1140) | (sub_sel & sub1140) | (and_sel & and1140) | (or_sel & or1140);
  assign y1141 = (add_sel & s1141) | (sub_sel & sub1141) | (and_sel & and1141) | (or_sel & or1141);
  assign y1142 = (add_sel & s1142) | (sub_sel & sub1142) | (and_sel & and1142) | (or_sel & or1142);
  assign y1143 = (add_sel & s1143) | (sub_sel & sub1143) | (and_sel & and1143) | (or_sel & or1143);
  assign y1144 = (add_sel & s1144) | (sub_sel & sub1144) | (and_sel & and1144) | (or_sel & or1144);
  assign y1145 = (add_sel & s1145) | (sub_sel & sub1145) | (and_sel & and1145) | (or_sel & or1145);
  assign y1146 = (add_sel & s1146) | (sub_sel & sub1146) | (and_sel & and1146) | (or_sel & or1146);
  assign y1147 = (add_sel & s1147) | (sub_sel & sub1147) | (and_sel & and1147) | (or_sel & or1147);
  assign y1148 = (add_sel & s1148) | (sub_sel & sub1148) | (and_sel & and1148) | (or_sel & or1148);
  assign y1149 = (add_sel & s1149) | (sub_sel & sub1149) | (and_sel & and1149) | (or_sel & or1149);
  assign y1150 = (add_sel & s1150) | (sub_sel & sub1150) | (and_sel & and1150) | (or_sel & or1150);
  assign y1151 = (add_sel & s1151) | (sub_sel & sub1151) | (and_sel & and1151) | (or_sel & or1151);
  assign y1152 = (add_sel & s1152) | (sub_sel & sub1152) | (and_sel & and1152) | (or_sel & or1152);
  assign y1153 = (add_sel & s1153) | (sub_sel & sub1153) | (and_sel & and1153) | (or_sel & or1153);
  assign y1154 = (add_sel & s1154) | (sub_sel & sub1154) | (and_sel & and1154) | (or_sel & or1154);
  assign y1155 = (add_sel & s1155) | (sub_sel & sub1155) | (and_sel & and1155) | (or_sel & or1155);
  assign y1156 = (add_sel & s1156) | (sub_sel & sub1156) | (and_sel & and1156) | (or_sel & or1156);
  assign y1157 = (add_sel & s1157) | (sub_sel & sub1157) | (and_sel & and1157) | (or_sel & or1157);
  assign y1158 = (add_sel & s1158) | (sub_sel & sub1158) | (and_sel & and1158) | (or_sel & or1158);
  assign y1159 = (add_sel & s1159) | (sub_sel & sub1159) | (and_sel & and1159) | (or_sel & or1159);
  assign y1160 = (add_sel & s1160) | (sub_sel & sub1160) | (and_sel & and1160) | (or_sel & or1160);
  assign y1161 = (add_sel & s1161) | (sub_sel & sub1161) | (and_sel & and1161) | (or_sel & or1161);
  assign y1162 = (add_sel & s1162) | (sub_sel & sub1162) | (and_sel & and1162) | (or_sel & or1162);
  assign y1163 = (add_sel & s1163) | (sub_sel & sub1163) | (and_sel & and1163) | (or_sel & or1163);
  assign y1164 = (add_sel & s1164) | (sub_sel & sub1164) | (and_sel & and1164) | (or_sel & or1164);
  assign y1165 = (add_sel & s1165) | (sub_sel & sub1165) | (and_sel & and1165) | (or_sel & or1165);
  assign y1166 = (add_sel & s1166) | (sub_sel & sub1166) | (and_sel & and1166) | (or_sel & or1166);
  assign y1167 = (add_sel & s1167) | (sub_sel & sub1167) | (and_sel & and1167) | (or_sel & or1167);
  assign y1168 = (add_sel & s1168) | (sub_sel & sub1168) | (and_sel & and1168) | (or_sel & or1168);
  assign y1169 = (add_sel & s1169) | (sub_sel & sub1169) | (and_sel & and1169) | (or_sel & or1169);
  assign y1170 = (add_sel & s1170) | (sub_sel & sub1170) | (and_sel & and1170) | (or_sel & or1170);
  assign y1171 = (add_sel & s1171) | (sub_sel & sub1171) | (and_sel & and1171) | (or_sel & or1171);
  assign y1172 = (add_sel & s1172) | (sub_sel & sub1172) | (and_sel & and1172) | (or_sel & or1172);
  assign y1173 = (add_sel & s1173) | (sub_sel & sub1173) | (and_sel & and1173) | (or_sel & or1173);
  assign y1174 = (add_sel & s1174) | (sub_sel & sub1174) | (and_sel & and1174) | (or_sel & or1174);
  assign y1175 = (add_sel & s1175) | (sub_sel & sub1175) | (and_sel & and1175) | (or_sel & or1175);
  assign y1176 = (add_sel & s1176) | (sub_sel & sub1176) | (and_sel & and1176) | (or_sel & or1176);
  assign y1177 = (add_sel & s1177) | (sub_sel & sub1177) | (and_sel & and1177) | (or_sel & or1177);
  assign y1178 = (add_sel & s1178) | (sub_sel & sub1178) | (and_sel & and1178) | (or_sel & or1178);
  assign y1179 = (add_sel & s1179) | (sub_sel & sub1179) | (and_sel & and1179) | (or_sel & or1179);
  assign y1180 = (add_sel & s1180) | (sub_sel & sub1180) | (and_sel & and1180) | (or_sel & or1180);
  assign y1181 = (add_sel & s1181) | (sub_sel & sub1181) | (and_sel & and1181) | (or_sel & or1181);
  assign y1182 = (add_sel & s1182) | (sub_sel & sub1182) | (and_sel & and1182) | (or_sel & or1182);
  assign y1183 = (add_sel & s1183) | (sub_sel & sub1183) | (and_sel & and1183) | (or_sel & or1183);
  assign y1184 = (add_sel & s1184) | (sub_sel & sub1184) | (and_sel & and1184) | (or_sel & or1184);
  assign y1185 = (add_sel & s1185) | (sub_sel & sub1185) | (and_sel & and1185) | (or_sel & or1185);
  assign y1186 = (add_sel & s1186) | (sub_sel & sub1186) | (and_sel & and1186) | (or_sel & or1186);
  assign y1187 = (add_sel & s1187) | (sub_sel & sub1187) | (and_sel & and1187) | (or_sel & or1187);
  assign y1188 = (add_sel & s1188) | (sub_sel & sub1188) | (and_sel & and1188) | (or_sel & or1188);
  assign y1189 = (add_sel & s1189) | (sub_sel & sub1189) | (and_sel & and1189) | (or_sel & or1189);
  assign y1190 = (add_sel & s1190) | (sub_sel & sub1190) | (and_sel & and1190) | (or_sel & or1190);
  assign y1191 = (add_sel & s1191) | (sub_sel & sub1191) | (and_sel & and1191) | (or_sel & or1191);
  assign y1192 = (add_sel & s1192) | (sub_sel & sub1192) | (and_sel & and1192) | (or_sel & or1192);
  assign y1193 = (add_sel & s1193) | (sub_sel & sub1193) | (and_sel & and1193) | (or_sel & or1193);
  assign y1194 = (add_sel & s1194) | (sub_sel & sub1194) | (and_sel & and1194) | (or_sel & or1194);
  assign y1195 = (add_sel & s1195) | (sub_sel & sub1195) | (and_sel & and1195) | (or_sel & or1195);
  assign y1196 = (add_sel & s1196) | (sub_sel & sub1196) | (and_sel & and1196) | (or_sel & or1196);
  assign y1197 = (add_sel & s1197) | (sub_sel & sub1197) | (and_sel & and1197) | (or_sel & or1197);
  assign y1198 = (add_sel & s1198) | (sub_sel & sub1198) | (and_sel & and1198) | (or_sel & or1198);
  assign y1199 = (add_sel & s1199) | (sub_sel & sub1199) | (and_sel & and1199) | (or_sel & or1199);
  assign y1200 = (add_sel & s1200) | (sub_sel & sub1200) | (and_sel & and1200) | (or_sel & or1200);
  assign y1201 = (add_sel & s1201) | (sub_sel & sub1201) | (and_sel & and1201) | (or_sel & or1201);
  assign y1202 = (add_sel & s1202) | (sub_sel & sub1202) | (and_sel & and1202) | (or_sel & or1202);
  assign y1203 = (add_sel & s1203) | (sub_sel & sub1203) | (and_sel & and1203) | (or_sel & or1203);
  assign y1204 = (add_sel & s1204) | (sub_sel & sub1204) | (and_sel & and1204) | (or_sel & or1204);
  assign y1205 = (add_sel & s1205) | (sub_sel & sub1205) | (and_sel & and1205) | (or_sel & or1205);
  assign y1206 = (add_sel & s1206) | (sub_sel & sub1206) | (and_sel & and1206) | (or_sel & or1206);
  assign y1207 = (add_sel & s1207) | (sub_sel & sub1207) | (and_sel & and1207) | (or_sel & or1207);
  assign y1208 = (add_sel & s1208) | (sub_sel & sub1208) | (and_sel & and1208) | (or_sel & or1208);
  assign y1209 = (add_sel & s1209) | (sub_sel & sub1209) | (and_sel & and1209) | (or_sel & or1209);
  assign y1210 = (add_sel & s1210) | (sub_sel & sub1210) | (and_sel & and1210) | (or_sel & or1210);
  assign y1211 = (add_sel & s1211) | (sub_sel & sub1211) | (and_sel & and1211) | (or_sel & or1211);
  assign y1212 = (add_sel & s1212) | (sub_sel & sub1212) | (and_sel & and1212) | (or_sel & or1212);
  assign y1213 = (add_sel & s1213) | (sub_sel & sub1213) | (and_sel & and1213) | (or_sel & or1213);
  assign y1214 = (add_sel & s1214) | (sub_sel & sub1214) | (and_sel & and1214) | (or_sel & or1214);
  assign y1215 = (add_sel & s1215) | (sub_sel & sub1215) | (and_sel & and1215) | (or_sel & or1215);
  assign y1216 = (add_sel & s1216) | (sub_sel & sub1216) | (and_sel & and1216) | (or_sel & or1216);
  assign y1217 = (add_sel & s1217) | (sub_sel & sub1217) | (and_sel & and1217) | (or_sel & or1217);
  assign y1218 = (add_sel & s1218) | (sub_sel & sub1218) | (and_sel & and1218) | (or_sel & or1218);
  assign y1219 = (add_sel & s1219) | (sub_sel & sub1219) | (and_sel & and1219) | (or_sel & or1219);
  assign y1220 = (add_sel & s1220) | (sub_sel & sub1220) | (and_sel & and1220) | (or_sel & or1220);
  assign y1221 = (add_sel & s1221) | (sub_sel & sub1221) | (and_sel & and1221) | (or_sel & or1221);
  assign y1222 = (add_sel & s1222) | (sub_sel & sub1222) | (and_sel & and1222) | (or_sel & or1222);
  assign y1223 = (add_sel & s1223) | (sub_sel & sub1223) | (and_sel & and1223) | (or_sel & or1223);
  assign y1224 = (add_sel & s1224) | (sub_sel & sub1224) | (and_sel & and1224) | (or_sel & or1224);
  assign y1225 = (add_sel & s1225) | (sub_sel & sub1225) | (and_sel & and1225) | (or_sel & or1225);
  assign y1226 = (add_sel & s1226) | (sub_sel & sub1226) | (and_sel & and1226) | (or_sel & or1226);
  assign y1227 = (add_sel & s1227) | (sub_sel & sub1227) | (and_sel & and1227) | (or_sel & or1227);
  assign y1228 = (add_sel & s1228) | (sub_sel & sub1228) | (and_sel & and1228) | (or_sel & or1228);
  assign y1229 = (add_sel & s1229) | (sub_sel & sub1229) | (and_sel & and1229) | (or_sel & or1229);
  assign y1230 = (add_sel & s1230) | (sub_sel & sub1230) | (and_sel & and1230) | (or_sel & or1230);
  assign y1231 = (add_sel & s1231) | (sub_sel & sub1231) | (and_sel & and1231) | (or_sel & or1231);
  assign y1232 = (add_sel & s1232) | (sub_sel & sub1232) | (and_sel & and1232) | (or_sel & or1232);
  assign y1233 = (add_sel & s1233) | (sub_sel & sub1233) | (and_sel & and1233) | (or_sel & or1233);
  assign y1234 = (add_sel & s1234) | (sub_sel & sub1234) | (and_sel & and1234) | (or_sel & or1234);
  assign y1235 = (add_sel & s1235) | (sub_sel & sub1235) | (and_sel & and1235) | (or_sel & or1235);
  assign y1236 = (add_sel & s1236) | (sub_sel & sub1236) | (and_sel & and1236) | (or_sel & or1236);
  assign y1237 = (add_sel & s1237) | (sub_sel & sub1237) | (and_sel & and1237) | (or_sel & or1237);
  assign y1238 = (add_sel & s1238) | (sub_sel & sub1238) | (and_sel & and1238) | (or_sel & or1238);
  assign y1239 = (add_sel & s1239) | (sub_sel & sub1239) | (and_sel & and1239) | (or_sel & or1239);
  assign y1240 = (add_sel & s1240) | (sub_sel & sub1240) | (and_sel & and1240) | (or_sel & or1240);
  assign y1241 = (add_sel & s1241) | (sub_sel & sub1241) | (and_sel & and1241) | (or_sel & or1241);
  assign y1242 = (add_sel & s1242) | (sub_sel & sub1242) | (and_sel & and1242) | (or_sel & or1242);
  assign y1243 = (add_sel & s1243) | (sub_sel & sub1243) | (and_sel & and1243) | (or_sel & or1243);
  assign y1244 = (add_sel & s1244) | (sub_sel & sub1244) | (and_sel & and1244) | (or_sel & or1244);
  assign y1245 = (add_sel & s1245) | (sub_sel & sub1245) | (and_sel & and1245) | (or_sel & or1245);
  assign y1246 = (add_sel & s1246) | (sub_sel & sub1246) | (and_sel & and1246) | (or_sel & or1246);
  assign y1247 = (add_sel & s1247) | (sub_sel & sub1247) | (and_sel & and1247) | (or_sel & or1247);
  assign y1248 = (add_sel & s1248) | (sub_sel & sub1248) | (and_sel & and1248) | (or_sel & or1248);
  assign y1249 = (add_sel & s1249) | (sub_sel & sub1249) | (and_sel & and1249) | (or_sel & or1249);
  assign y1250 = (add_sel & s1250) | (sub_sel & sub1250) | (and_sel & and1250) | (or_sel & or1250);
  assign y1251 = (add_sel & s1251) | (sub_sel & sub1251) | (and_sel & and1251) | (or_sel & or1251);
  assign y1252 = (add_sel & s1252) | (sub_sel & sub1252) | (and_sel & and1252) | (or_sel & or1252);
  assign y1253 = (add_sel & s1253) | (sub_sel & sub1253) | (and_sel & and1253) | (or_sel & or1253);
  assign y1254 = (add_sel & s1254) | (sub_sel & sub1254) | (and_sel & and1254) | (or_sel & or1254);
  assign y1255 = (add_sel & s1255) | (sub_sel & sub1255) | (and_sel & and1255) | (or_sel & or1255);
  assign y1256 = (add_sel & s1256) | (sub_sel & sub1256) | (and_sel & and1256) | (or_sel & or1256);
  assign y1257 = (add_sel & s1257) | (sub_sel & sub1257) | (and_sel & and1257) | (or_sel & or1257);
  assign y1258 = (add_sel & s1258) | (sub_sel & sub1258) | (and_sel & and1258) | (or_sel & or1258);
  assign y1259 = (add_sel & s1259) | (sub_sel & sub1259) | (and_sel & and1259) | (or_sel & or1259);
  assign y1260 = (add_sel & s1260) | (sub_sel & sub1260) | (and_sel & and1260) | (or_sel & or1260);
  assign y1261 = (add_sel & s1261) | (sub_sel & sub1261) | (and_sel & and1261) | (or_sel & or1261);
  assign y1262 = (add_sel & s1262) | (sub_sel & sub1262) | (and_sel & and1262) | (or_sel & or1262);
  assign y1263 = (add_sel & s1263) | (sub_sel & sub1263) | (and_sel & and1263) | (or_sel & or1263);
  assign y1264 = (add_sel & s1264) | (sub_sel & sub1264) | (and_sel & and1264) | (or_sel & or1264);
  assign y1265 = (add_sel & s1265) | (sub_sel & sub1265) | (and_sel & and1265) | (or_sel & or1265);
  assign y1266 = (add_sel & s1266) | (sub_sel & sub1266) | (and_sel & and1266) | (or_sel & or1266);
  assign y1267 = (add_sel & s1267) | (sub_sel & sub1267) | (and_sel & and1267) | (or_sel & or1267);
  assign y1268 = (add_sel & s1268) | (sub_sel & sub1268) | (and_sel & and1268) | (or_sel & or1268);
  assign y1269 = (add_sel & s1269) | (sub_sel & sub1269) | (and_sel & and1269) | (or_sel & or1269);
  assign y1270 = (add_sel & s1270) | (sub_sel & sub1270) | (and_sel & and1270) | (or_sel & or1270);
  assign y1271 = (add_sel & s1271) | (sub_sel & sub1271) | (and_sel & and1271) | (or_sel & or1271);
  assign y1272 = (add_sel & s1272) | (sub_sel & sub1272) | (and_sel & and1272) | (or_sel & or1272);
  assign y1273 = (add_sel & s1273) | (sub_sel & sub1273) | (and_sel & and1273) | (or_sel & or1273);
  assign y1274 = (add_sel & s1274) | (sub_sel & sub1274) | (and_sel & and1274) | (or_sel & or1274);
  assign y1275 = (add_sel & s1275) | (sub_sel & sub1275) | (and_sel & and1275) | (or_sel & or1275);
  assign y1276 = (add_sel & s1276) | (sub_sel & sub1276) | (and_sel & and1276) | (or_sel & or1276);
  assign y1277 = (add_sel & s1277) | (sub_sel & sub1277) | (and_sel & and1277) | (or_sel & or1277);
  assign y1278 = (add_sel & s1278) | (sub_sel & sub1278) | (and_sel & and1278) | (or_sel & or1278);
  assign y1279 = (add_sel & s1279) | (sub_sel & sub1279) | (and_sel & and1279) | (or_sel & or1279);
  assign y1280 = (add_sel & s1280) | (sub_sel & sub1280) | (and_sel & and1280) | (or_sel & or1280);
  assign y1281 = (add_sel & s1281) | (sub_sel & sub1281) | (and_sel & and1281) | (or_sel & or1281);
  assign y1282 = (add_sel & s1282) | (sub_sel & sub1282) | (and_sel & and1282) | (or_sel & or1282);
  assign y1283 = (add_sel & s1283) | (sub_sel & sub1283) | (and_sel & and1283) | (or_sel & or1283);
  assign y1284 = (add_sel & s1284) | (sub_sel & sub1284) | (and_sel & and1284) | (or_sel & or1284);
  assign y1285 = (add_sel & s1285) | (sub_sel & sub1285) | (and_sel & and1285) | (or_sel & or1285);
  assign y1286 = (add_sel & s1286) | (sub_sel & sub1286) | (and_sel & and1286) | (or_sel & or1286);
  assign y1287 = (add_sel & s1287) | (sub_sel & sub1287) | (and_sel & and1287) | (or_sel & or1287);
  assign y1288 = (add_sel & s1288) | (sub_sel & sub1288) | (and_sel & and1288) | (or_sel & or1288);
  assign y1289 = (add_sel & s1289) | (sub_sel & sub1289) | (and_sel & and1289) | (or_sel & or1289);
  assign y1290 = (add_sel & s1290) | (sub_sel & sub1290) | (and_sel & and1290) | (or_sel & or1290);
  assign y1291 = (add_sel & s1291) | (sub_sel & sub1291) | (and_sel & and1291) | (or_sel & or1291);
  assign y1292 = (add_sel & s1292) | (sub_sel & sub1292) | (and_sel & and1292) | (or_sel & or1292);
  assign y1293 = (add_sel & s1293) | (sub_sel & sub1293) | (and_sel & and1293) | (or_sel & or1293);
  assign y1294 = (add_sel & s1294) | (sub_sel & sub1294) | (and_sel & and1294) | (or_sel & or1294);
  assign y1295 = (add_sel & s1295) | (sub_sel & sub1295) | (and_sel & and1295) | (or_sel & or1295);
  assign y1296 = (add_sel & s1296) | (sub_sel & sub1296) | (and_sel & and1296) | (or_sel & or1296);
  assign y1297 = (add_sel & s1297) | (sub_sel & sub1297) | (and_sel & and1297) | (or_sel & or1297);
  assign y1298 = (add_sel & s1298) | (sub_sel & sub1298) | (and_sel & and1298) | (or_sel & or1298);
  assign y1299 = (add_sel & s1299) | (sub_sel & sub1299) | (and_sel & and1299) | (or_sel & or1299);
  assign y1300 = (add_sel & s1300) | (sub_sel & sub1300) | (and_sel & and1300) | (or_sel & or1300);
  assign y1301 = (add_sel & s1301) | (sub_sel & sub1301) | (and_sel & and1301) | (or_sel & or1301);
  assign y1302 = (add_sel & s1302) | (sub_sel & sub1302) | (and_sel & and1302) | (or_sel & or1302);
  assign y1303 = (add_sel & s1303) | (sub_sel & sub1303) | (and_sel & and1303) | (or_sel & or1303);
  assign y1304 = (add_sel & s1304) | (sub_sel & sub1304) | (and_sel & and1304) | (or_sel & or1304);
  assign y1305 = (add_sel & s1305) | (sub_sel & sub1305) | (and_sel & and1305) | (or_sel & or1305);
  assign y1306 = (add_sel & s1306) | (sub_sel & sub1306) | (and_sel & and1306) | (or_sel & or1306);
  assign y1307 = (add_sel & s1307) | (sub_sel & sub1307) | (and_sel & and1307) | (or_sel & or1307);
  assign y1308 = (add_sel & s1308) | (sub_sel & sub1308) | (and_sel & and1308) | (or_sel & or1308);
  assign y1309 = (add_sel & s1309) | (sub_sel & sub1309) | (and_sel & and1309) | (or_sel & or1309);
  assign y1310 = (add_sel & s1310) | (sub_sel & sub1310) | (and_sel & and1310) | (or_sel & or1310);
  assign y1311 = (add_sel & s1311) | (sub_sel & sub1311) | (and_sel & and1311) | (or_sel & or1311);
  assign y1312 = (add_sel & s1312) | (sub_sel & sub1312) | (and_sel & and1312) | (or_sel & or1312);
  assign y1313 = (add_sel & s1313) | (sub_sel & sub1313) | (and_sel & and1313) | (or_sel & or1313);
  assign y1314 = (add_sel & s1314) | (sub_sel & sub1314) | (and_sel & and1314) | (or_sel & or1314);
  assign y1315 = (add_sel & s1315) | (sub_sel & sub1315) | (and_sel & and1315) | (or_sel & or1315);
  assign y1316 = (add_sel & s1316) | (sub_sel & sub1316) | (and_sel & and1316) | (or_sel & or1316);
  assign y1317 = (add_sel & s1317) | (sub_sel & sub1317) | (and_sel & and1317) | (or_sel & or1317);
  assign y1318 = (add_sel & s1318) | (sub_sel & sub1318) | (and_sel & and1318) | (or_sel & or1318);
  assign y1319 = (add_sel & s1319) | (sub_sel & sub1319) | (and_sel & and1319) | (or_sel & or1319);
  assign y1320 = (add_sel & s1320) | (sub_sel & sub1320) | (and_sel & and1320) | (or_sel & or1320);
  assign y1321 = (add_sel & s1321) | (sub_sel & sub1321) | (and_sel & and1321) | (or_sel & or1321);
  assign y1322 = (add_sel & s1322) | (sub_sel & sub1322) | (and_sel & and1322) | (or_sel & or1322);
  assign y1323 = (add_sel & s1323) | (sub_sel & sub1323) | (and_sel & and1323) | (or_sel & or1323);
  assign y1324 = (add_sel & s1324) | (sub_sel & sub1324) | (and_sel & and1324) | (or_sel & or1324);
  assign y1325 = (add_sel & s1325) | (sub_sel & sub1325) | (and_sel & and1325) | (or_sel & or1325);
  assign y1326 = (add_sel & s1326) | (sub_sel & sub1326) | (and_sel & and1326) | (or_sel & or1326);
  assign y1327 = (add_sel & s1327) | (sub_sel & sub1327) | (and_sel & and1327) | (or_sel & or1327);
  assign y1328 = (add_sel & s1328) | (sub_sel & sub1328) | (and_sel & and1328) | (or_sel & or1328);
  assign y1329 = (add_sel & s1329) | (sub_sel & sub1329) | (and_sel & and1329) | (or_sel & or1329);
  assign y1330 = (add_sel & s1330) | (sub_sel & sub1330) | (and_sel & and1330) | (or_sel & or1330);
  assign y1331 = (add_sel & s1331) | (sub_sel & sub1331) | (and_sel & and1331) | (or_sel & or1331);
  assign y1332 = (add_sel & s1332) | (sub_sel & sub1332) | (and_sel & and1332) | (or_sel & or1332);
  assign y1333 = (add_sel & s1333) | (sub_sel & sub1333) | (and_sel & and1333) | (or_sel & or1333);
  assign y1334 = (add_sel & s1334) | (sub_sel & sub1334) | (and_sel & and1334) | (or_sel & or1334);
  assign y1335 = (add_sel & s1335) | (sub_sel & sub1335) | (and_sel & and1335) | (or_sel & or1335);
  assign y1336 = (add_sel & s1336) | (sub_sel & sub1336) | (and_sel & and1336) | (or_sel & or1336);
  assign y1337 = (add_sel & s1337) | (sub_sel & sub1337) | (and_sel & and1337) | (or_sel & or1337);
  assign y1338 = (add_sel & s1338) | (sub_sel & sub1338) | (and_sel & and1338) | (or_sel & or1338);
  assign y1339 = (add_sel & s1339) | (sub_sel & sub1339) | (and_sel & and1339) | (or_sel & or1339);
  assign y1340 = (add_sel & s1340) | (sub_sel & sub1340) | (and_sel & and1340) | (or_sel & or1340);
  assign y1341 = (add_sel & s1341) | (sub_sel & sub1341) | (and_sel & and1341) | (or_sel & or1341);
  assign y1342 = (add_sel & s1342) | (sub_sel & sub1342) | (and_sel & and1342) | (or_sel & or1342);
  assign y1343 = (add_sel & s1343) | (sub_sel & sub1343) | (and_sel & and1343) | (or_sel & or1343);
  assign y1344 = (add_sel & s1344) | (sub_sel & sub1344) | (and_sel & and1344) | (or_sel & or1344);
  assign y1345 = (add_sel & s1345) | (sub_sel & sub1345) | (and_sel & and1345) | (or_sel & or1345);
  assign y1346 = (add_sel & s1346) | (sub_sel & sub1346) | (and_sel & and1346) | (or_sel & or1346);
  assign y1347 = (add_sel & s1347) | (sub_sel & sub1347) | (and_sel & and1347) | (or_sel & or1347);
  assign y1348 = (add_sel & s1348) | (sub_sel & sub1348) | (and_sel & and1348) | (or_sel & or1348);
  assign y1349 = (add_sel & s1349) | (sub_sel & sub1349) | (and_sel & and1349) | (or_sel & or1349);
  assign y1350 = (add_sel & s1350) | (sub_sel & sub1350) | (and_sel & and1350) | (or_sel & or1350);
  assign y1351 = (add_sel & s1351) | (sub_sel & sub1351) | (and_sel & and1351) | (or_sel & or1351);
  assign y1352 = (add_sel & s1352) | (sub_sel & sub1352) | (and_sel & and1352) | (or_sel & or1352);
  assign y1353 = (add_sel & s1353) | (sub_sel & sub1353) | (and_sel & and1353) | (or_sel & or1353);
  assign y1354 = (add_sel & s1354) | (sub_sel & sub1354) | (and_sel & and1354) | (or_sel & or1354);
  assign y1355 = (add_sel & s1355) | (sub_sel & sub1355) | (and_sel & and1355) | (or_sel & or1355);
  assign y1356 = (add_sel & s1356) | (sub_sel & sub1356) | (and_sel & and1356) | (or_sel & or1356);
  assign y1357 = (add_sel & s1357) | (sub_sel & sub1357) | (and_sel & and1357) | (or_sel & or1357);
  assign y1358 = (add_sel & s1358) | (sub_sel & sub1358) | (and_sel & and1358) | (or_sel & or1358);
  assign y1359 = (add_sel & s1359) | (sub_sel & sub1359) | (and_sel & and1359) | (or_sel & or1359);
  assign y1360 = (add_sel & s1360) | (sub_sel & sub1360) | (and_sel & and1360) | (or_sel & or1360);
  assign y1361 = (add_sel & s1361) | (sub_sel & sub1361) | (and_sel & and1361) | (or_sel & or1361);
  assign y1362 = (add_sel & s1362) | (sub_sel & sub1362) | (and_sel & and1362) | (or_sel & or1362);
  assign y1363 = (add_sel & s1363) | (sub_sel & sub1363) | (and_sel & and1363) | (or_sel & or1363);
  assign y1364 = (add_sel & s1364) | (sub_sel & sub1364) | (and_sel & and1364) | (or_sel & or1364);
  assign y1365 = (add_sel & s1365) | (sub_sel & sub1365) | (and_sel & and1365) | (or_sel & or1365);
  assign y1366 = (add_sel & s1366) | (sub_sel & sub1366) | (and_sel & and1366) | (or_sel & or1366);
  assign y1367 = (add_sel & s1367) | (sub_sel & sub1367) | (and_sel & and1367) | (or_sel & or1367);
  assign y1368 = (add_sel & s1368) | (sub_sel & sub1368) | (and_sel & and1368) | (or_sel & or1368);
  assign y1369 = (add_sel & s1369) | (sub_sel & sub1369) | (and_sel & and1369) | (or_sel & or1369);
  assign y1370 = (add_sel & s1370) | (sub_sel & sub1370) | (and_sel & and1370) | (or_sel & or1370);
  assign y1371 = (add_sel & s1371) | (sub_sel & sub1371) | (and_sel & and1371) | (or_sel & or1371);
  assign y1372 = (add_sel & s1372) | (sub_sel & sub1372) | (and_sel & and1372) | (or_sel & or1372);
  assign y1373 = (add_sel & s1373) | (sub_sel & sub1373) | (and_sel & and1373) | (or_sel & or1373);
  assign y1374 = (add_sel & s1374) | (sub_sel & sub1374) | (and_sel & and1374) | (or_sel & or1374);
  assign y1375 = (add_sel & s1375) | (sub_sel & sub1375) | (and_sel & and1375) | (or_sel & or1375);
  assign y1376 = (add_sel & s1376) | (sub_sel & sub1376) | (and_sel & and1376) | (or_sel & or1376);
  assign y1377 = (add_sel & s1377) | (sub_sel & sub1377) | (and_sel & and1377) | (or_sel & or1377);
  assign y1378 = (add_sel & s1378) | (sub_sel & sub1378) | (and_sel & and1378) | (or_sel & or1378);
  assign y1379 = (add_sel & s1379) | (sub_sel & sub1379) | (and_sel & and1379) | (or_sel & or1379);
  assign y1380 = (add_sel & s1380) | (sub_sel & sub1380) | (and_sel & and1380) | (or_sel & or1380);
  assign y1381 = (add_sel & s1381) | (sub_sel & sub1381) | (and_sel & and1381) | (or_sel & or1381);
  assign y1382 = (add_sel & s1382) | (sub_sel & sub1382) | (and_sel & and1382) | (or_sel & or1382);
  assign y1383 = (add_sel & s1383) | (sub_sel & sub1383) | (and_sel & and1383) | (or_sel & or1383);
  assign y1384 = (add_sel & s1384) | (sub_sel & sub1384) | (and_sel & and1384) | (or_sel & or1384);
  assign y1385 = (add_sel & s1385) | (sub_sel & sub1385) | (and_sel & and1385) | (or_sel & or1385);
  assign y1386 = (add_sel & s1386) | (sub_sel & sub1386) | (and_sel & and1386) | (or_sel & or1386);
  assign y1387 = (add_sel & s1387) | (sub_sel & sub1387) | (and_sel & and1387) | (or_sel & or1387);
  assign y1388 = (add_sel & s1388) | (sub_sel & sub1388) | (and_sel & and1388) | (or_sel & or1388);
  assign y1389 = (add_sel & s1389) | (sub_sel & sub1389) | (and_sel & and1389) | (or_sel & or1389);
  assign y1390 = (add_sel & s1390) | (sub_sel & sub1390) | (and_sel & and1390) | (or_sel & or1390);
  assign y1391 = (add_sel & s1391) | (sub_sel & sub1391) | (and_sel & and1391) | (or_sel & or1391);
  assign y1392 = (add_sel & s1392) | (sub_sel & sub1392) | (and_sel & and1392) | (or_sel & or1392);
  assign y1393 = (add_sel & s1393) | (sub_sel & sub1393) | (and_sel & and1393) | (or_sel & or1393);
  assign y1394 = (add_sel & s1394) | (sub_sel & sub1394) | (and_sel & and1394) | (or_sel & or1394);
  assign y1395 = (add_sel & s1395) | (sub_sel & sub1395) | (and_sel & and1395) | (or_sel & or1395);
  assign y1396 = (add_sel & s1396) | (sub_sel & sub1396) | (and_sel & and1396) | (or_sel & or1396);
  assign y1397 = (add_sel & s1397) | (sub_sel & sub1397) | (and_sel & and1397) | (or_sel & or1397);
  assign y1398 = (add_sel & s1398) | (sub_sel & sub1398) | (and_sel & and1398) | (or_sel & or1398);
  assign y1399 = (add_sel & s1399) | (sub_sel & sub1399) | (and_sel & and1399) | (or_sel & or1399);
  assign y1400 = (add_sel & s1400) | (sub_sel & sub1400) | (and_sel & and1400) | (or_sel & or1400);
  assign y1401 = (add_sel & s1401) | (sub_sel & sub1401) | (and_sel & and1401) | (or_sel & or1401);
  assign y1402 = (add_sel & s1402) | (sub_sel & sub1402) | (and_sel & and1402) | (or_sel & or1402);
  assign y1403 = (add_sel & s1403) | (sub_sel & sub1403) | (and_sel & and1403) | (or_sel & or1403);
  assign y1404 = (add_sel & s1404) | (sub_sel & sub1404) | (and_sel & and1404) | (or_sel & or1404);
  assign y1405 = (add_sel & s1405) | (sub_sel & sub1405) | (and_sel & and1405) | (or_sel & or1405);
  assign y1406 = (add_sel & s1406) | (sub_sel & sub1406) | (and_sel & and1406) | (or_sel & or1406);
  assign y1407 = (add_sel & s1407) | (sub_sel & sub1407) | (and_sel & and1407) | (or_sel & or1407);
  assign y1408 = (add_sel & s1408) | (sub_sel & sub1408) | (and_sel & and1408) | (or_sel & or1408);
  assign y1409 = (add_sel & s1409) | (sub_sel & sub1409) | (and_sel & and1409) | (or_sel & or1409);
  assign y1410 = (add_sel & s1410) | (sub_sel & sub1410) | (and_sel & and1410) | (or_sel & or1410);
  assign y1411 = (add_sel & s1411) | (sub_sel & sub1411) | (and_sel & and1411) | (or_sel & or1411);
  assign y1412 = (add_sel & s1412) | (sub_sel & sub1412) | (and_sel & and1412) | (or_sel & or1412);
  assign y1413 = (add_sel & s1413) | (sub_sel & sub1413) | (and_sel & and1413) | (or_sel & or1413);
  assign y1414 = (add_sel & s1414) | (sub_sel & sub1414) | (and_sel & and1414) | (or_sel & or1414);
  assign y1415 = (add_sel & s1415) | (sub_sel & sub1415) | (and_sel & and1415) | (or_sel & or1415);
  assign y1416 = (add_sel & s1416) | (sub_sel & sub1416) | (and_sel & and1416) | (or_sel & or1416);
  assign y1417 = (add_sel & s1417) | (sub_sel & sub1417) | (and_sel & and1417) | (or_sel & or1417);
  assign y1418 = (add_sel & s1418) | (sub_sel & sub1418) | (and_sel & and1418) | (or_sel & or1418);
  assign y1419 = (add_sel & s1419) | (sub_sel & sub1419) | (and_sel & and1419) | (or_sel & or1419);
  assign y1420 = (add_sel & s1420) | (sub_sel & sub1420) | (and_sel & and1420) | (or_sel & or1420);
  assign y1421 = (add_sel & s1421) | (sub_sel & sub1421) | (and_sel & and1421) | (or_sel & or1421);
  assign y1422 = (add_sel & s1422) | (sub_sel & sub1422) | (and_sel & and1422) | (or_sel & or1422);
  assign y1423 = (add_sel & s1423) | (sub_sel & sub1423) | (and_sel & and1423) | (or_sel & or1423);
  assign y1424 = (add_sel & s1424) | (sub_sel & sub1424) | (and_sel & and1424) | (or_sel & or1424);
  assign y1425 = (add_sel & s1425) | (sub_sel & sub1425) | (and_sel & and1425) | (or_sel & or1425);
  assign y1426 = (add_sel & s1426) | (sub_sel & sub1426) | (and_sel & and1426) | (or_sel & or1426);
  assign y1427 = (add_sel & s1427) | (sub_sel & sub1427) | (and_sel & and1427) | (or_sel & or1427);
  assign y1428 = (add_sel & s1428) | (sub_sel & sub1428) | (and_sel & and1428) | (or_sel & or1428);
  assign y1429 = (add_sel & s1429) | (sub_sel & sub1429) | (and_sel & and1429) | (or_sel & or1429);
  assign y1430 = (add_sel & s1430) | (sub_sel & sub1430) | (and_sel & and1430) | (or_sel & or1430);
  assign y1431 = (add_sel & s1431) | (sub_sel & sub1431) | (and_sel & and1431) | (or_sel & or1431);
  assign y1432 = (add_sel & s1432) | (sub_sel & sub1432) | (and_sel & and1432) | (or_sel & or1432);
  assign y1433 = (add_sel & s1433) | (sub_sel & sub1433) | (and_sel & and1433) | (or_sel & or1433);
  assign y1434 = (add_sel & s1434) | (sub_sel & sub1434) | (and_sel & and1434) | (or_sel & or1434);
  assign y1435 = (add_sel & s1435) | (sub_sel & sub1435) | (and_sel & and1435) | (or_sel & or1435);
  assign y1436 = (add_sel & s1436) | (sub_sel & sub1436) | (and_sel & and1436) | (or_sel & or1436);
  assign y1437 = (add_sel & s1437) | (sub_sel & sub1437) | (and_sel & and1437) | (or_sel & or1437);
  assign y1438 = (add_sel & s1438) | (sub_sel & sub1438) | (and_sel & and1438) | (or_sel & or1438);
  assign y1439 = (add_sel & s1439) | (sub_sel & sub1439) | (and_sel & and1439) | (or_sel & or1439);
  assign y1440 = (add_sel & s1440) | (sub_sel & sub1440) | (and_sel & and1440) | (or_sel & or1440);
  assign y1441 = (add_sel & s1441) | (sub_sel & sub1441) | (and_sel & and1441) | (or_sel & or1441);
  assign y1442 = (add_sel & s1442) | (sub_sel & sub1442) | (and_sel & and1442) | (or_sel & or1442);
  assign y1443 = (add_sel & s1443) | (sub_sel & sub1443) | (and_sel & and1443) | (or_sel & or1443);
  assign y1444 = (add_sel & s1444) | (sub_sel & sub1444) | (and_sel & and1444) | (or_sel & or1444);
  assign y1445 = (add_sel & s1445) | (sub_sel & sub1445) | (and_sel & and1445) | (or_sel & or1445);
  assign y1446 = (add_sel & s1446) | (sub_sel & sub1446) | (and_sel & and1446) | (or_sel & or1446);
  assign y1447 = (add_sel & s1447) | (sub_sel & sub1447) | (and_sel & and1447) | (or_sel & or1447);
  assign y1448 = (add_sel & s1448) | (sub_sel & sub1448) | (and_sel & and1448) | (or_sel & or1448);
  assign y1449 = (add_sel & s1449) | (sub_sel & sub1449) | (and_sel & and1449) | (or_sel & or1449);
  assign y1450 = (add_sel & s1450) | (sub_sel & sub1450) | (and_sel & and1450) | (or_sel & or1450);
  assign y1451 = (add_sel & s1451) | (sub_sel & sub1451) | (and_sel & and1451) | (or_sel & or1451);
  assign y1452 = (add_sel & s1452) | (sub_sel & sub1452) | (and_sel & and1452) | (or_sel & or1452);
  assign y1453 = (add_sel & s1453) | (sub_sel & sub1453) | (and_sel & and1453) | (or_sel & or1453);
  assign y1454 = (add_sel & s1454) | (sub_sel & sub1454) | (and_sel & and1454) | (or_sel & or1454);
  assign y1455 = (add_sel & s1455) | (sub_sel & sub1455) | (and_sel & and1455) | (or_sel & or1455);
  assign y1456 = (add_sel & s1456) | (sub_sel & sub1456) | (and_sel & and1456) | (or_sel & or1456);
  assign y1457 = (add_sel & s1457) | (sub_sel & sub1457) | (and_sel & and1457) | (or_sel & or1457);
  assign y1458 = (add_sel & s1458) | (sub_sel & sub1458) | (and_sel & and1458) | (or_sel & or1458);
  assign y1459 = (add_sel & s1459) | (sub_sel & sub1459) | (and_sel & and1459) | (or_sel & or1459);
  assign y1460 = (add_sel & s1460) | (sub_sel & sub1460) | (and_sel & and1460) | (or_sel & or1460);
  assign y1461 = (add_sel & s1461) | (sub_sel & sub1461) | (and_sel & and1461) | (or_sel & or1461);
  assign y1462 = (add_sel & s1462) | (sub_sel & sub1462) | (and_sel & and1462) | (or_sel & or1462);
  assign y1463 = (add_sel & s1463) | (sub_sel & sub1463) | (and_sel & and1463) | (or_sel & or1463);
  assign y1464 = (add_sel & s1464) | (sub_sel & sub1464) | (and_sel & and1464) | (or_sel & or1464);
  assign y1465 = (add_sel & s1465) | (sub_sel & sub1465) | (and_sel & and1465) | (or_sel & or1465);
  assign y1466 = (add_sel & s1466) | (sub_sel & sub1466) | (and_sel & and1466) | (or_sel & or1466);
  assign y1467 = (add_sel & s1467) | (sub_sel & sub1467) | (and_sel & and1467) | (or_sel & or1467);
  assign y1468 = (add_sel & s1468) | (sub_sel & sub1468) | (and_sel & and1468) | (or_sel & or1468);
  assign y1469 = (add_sel & s1469) | (sub_sel & sub1469) | (and_sel & and1469) | (or_sel & or1469);
  assign y1470 = (add_sel & s1470) | (sub_sel & sub1470) | (and_sel & and1470) | (or_sel & or1470);
  assign y1471 = (add_sel & s1471) | (sub_sel & sub1471) | (and_sel & and1471) | (or_sel & or1471);
  assign y1472 = (add_sel & s1472) | (sub_sel & sub1472) | (and_sel & and1472) | (or_sel & or1472);
  assign y1473 = (add_sel & s1473) | (sub_sel & sub1473) | (and_sel & and1473) | (or_sel & or1473);
  assign y1474 = (add_sel & s1474) | (sub_sel & sub1474) | (and_sel & and1474) | (or_sel & or1474);
  assign y1475 = (add_sel & s1475) | (sub_sel & sub1475) | (and_sel & and1475) | (or_sel & or1475);
  assign y1476 = (add_sel & s1476) | (sub_sel & sub1476) | (and_sel & and1476) | (or_sel & or1476);
  assign y1477 = (add_sel & s1477) | (sub_sel & sub1477) | (and_sel & and1477) | (or_sel & or1477);
  assign y1478 = (add_sel & s1478) | (sub_sel & sub1478) | (and_sel & and1478) | (or_sel & or1478);
  assign y1479 = (add_sel & s1479) | (sub_sel & sub1479) | (and_sel & and1479) | (or_sel & or1479);
  assign y1480 = (add_sel & s1480) | (sub_sel & sub1480) | (and_sel & and1480) | (or_sel & or1480);
  assign y1481 = (add_sel & s1481) | (sub_sel & sub1481) | (and_sel & and1481) | (or_sel & or1481);
  assign y1482 = (add_sel & s1482) | (sub_sel & sub1482) | (and_sel & and1482) | (or_sel & or1482);
  assign y1483 = (add_sel & s1483) | (sub_sel & sub1483) | (and_sel & and1483) | (or_sel & or1483);
  assign y1484 = (add_sel & s1484) | (sub_sel & sub1484) | (and_sel & and1484) | (or_sel & or1484);
  assign y1485 = (add_sel & s1485) | (sub_sel & sub1485) | (and_sel & and1485) | (or_sel & or1485);
  assign y1486 = (add_sel & s1486) | (sub_sel & sub1486) | (and_sel & and1486) | (or_sel & or1486);
  assign y1487 = (add_sel & s1487) | (sub_sel & sub1487) | (and_sel & and1487) | (or_sel & or1487);
  assign y1488 = (add_sel & s1488) | (sub_sel & sub1488) | (and_sel & and1488) | (or_sel & or1488);
  assign y1489 = (add_sel & s1489) | (sub_sel & sub1489) | (and_sel & and1489) | (or_sel & or1489);
  assign y1490 = (add_sel & s1490) | (sub_sel & sub1490) | (and_sel & and1490) | (or_sel & or1490);
  assign y1491 = (add_sel & s1491) | (sub_sel & sub1491) | (and_sel & and1491) | (or_sel & or1491);
  assign y1492 = (add_sel & s1492) | (sub_sel & sub1492) | (and_sel & and1492) | (or_sel & or1492);
  assign y1493 = (add_sel & s1493) | (sub_sel & sub1493) | (and_sel & and1493) | (or_sel & or1493);
  assign y1494 = (add_sel & s1494) | (sub_sel & sub1494) | (and_sel & and1494) | (or_sel & or1494);
  assign y1495 = (add_sel & s1495) | (sub_sel & sub1495) | (and_sel & and1495) | (or_sel & or1495);
  assign y1496 = (add_sel & s1496) | (sub_sel & sub1496) | (and_sel & and1496) | (or_sel & or1496);
  assign y1497 = (add_sel & s1497) | (sub_sel & sub1497) | (and_sel & and1497) | (or_sel & or1497);
  assign y1498 = (add_sel & s1498) | (sub_sel & sub1498) | (and_sel & and1498) | (or_sel & or1498);
  assign y1499 = (add_sel & s1499) | (sub_sel & sub1499) | (and_sel & and1499) | (or_sel & or1499);
  assign y1500 = (add_sel & s1500) | (sub_sel & sub1500) | (and_sel & and1500) | (or_sel & or1500);
  assign y1501 = (add_sel & s1501) | (sub_sel & sub1501) | (and_sel & and1501) | (or_sel & or1501);
  assign y1502 = (add_sel & s1502) | (sub_sel & sub1502) | (and_sel & and1502) | (or_sel & or1502);
  assign y1503 = (add_sel & s1503) | (sub_sel & sub1503) | (and_sel & and1503) | (or_sel & or1503);
  assign y1504 = (add_sel & s1504) | (sub_sel & sub1504) | (and_sel & and1504) | (or_sel & or1504);
  assign y1505 = (add_sel & s1505) | (sub_sel & sub1505) | (and_sel & and1505) | (or_sel & or1505);
  assign y1506 = (add_sel & s1506) | (sub_sel & sub1506) | (and_sel & and1506) | (or_sel & or1506);
  assign y1507 = (add_sel & s1507) | (sub_sel & sub1507) | (and_sel & and1507) | (or_sel & or1507);
  assign y1508 = (add_sel & s1508) | (sub_sel & sub1508) | (and_sel & and1508) | (or_sel & or1508);
  assign y1509 = (add_sel & s1509) | (sub_sel & sub1509) | (and_sel & and1509) | (or_sel & or1509);
  assign y1510 = (add_sel & s1510) | (sub_sel & sub1510) | (and_sel & and1510) | (or_sel & or1510);
  assign y1511 = (add_sel & s1511) | (sub_sel & sub1511) | (and_sel & and1511) | (or_sel & or1511);
  assign y1512 = (add_sel & s1512) | (sub_sel & sub1512) | (and_sel & and1512) | (or_sel & or1512);
  assign y1513 = (add_sel & s1513) | (sub_sel & sub1513) | (and_sel & and1513) | (or_sel & or1513);
  assign y1514 = (add_sel & s1514) | (sub_sel & sub1514) | (and_sel & and1514) | (or_sel & or1514);
  assign y1515 = (add_sel & s1515) | (sub_sel & sub1515) | (and_sel & and1515) | (or_sel & or1515);
  assign y1516 = (add_sel & s1516) | (sub_sel & sub1516) | (and_sel & and1516) | (or_sel & or1516);
  assign y1517 = (add_sel & s1517) | (sub_sel & sub1517) | (and_sel & and1517) | (or_sel & or1517);
  assign y1518 = (add_sel & s1518) | (sub_sel & sub1518) | (and_sel & and1518) | (or_sel & or1518);
  assign y1519 = (add_sel & s1519) | (sub_sel & sub1519) | (and_sel & and1519) | (or_sel & or1519);
  assign y1520 = (add_sel & s1520) | (sub_sel & sub1520) | (and_sel & and1520) | (or_sel & or1520);
  assign y1521 = (add_sel & s1521) | (sub_sel & sub1521) | (and_sel & and1521) | (or_sel & or1521);
  assign y1522 = (add_sel & s1522) | (sub_sel & sub1522) | (and_sel & and1522) | (or_sel & or1522);
  assign y1523 = (add_sel & s1523) | (sub_sel & sub1523) | (and_sel & and1523) | (or_sel & or1523);
  assign y1524 = (add_sel & s1524) | (sub_sel & sub1524) | (and_sel & and1524) | (or_sel & or1524);
  assign y1525 = (add_sel & s1525) | (sub_sel & sub1525) | (and_sel & and1525) | (or_sel & or1525);
  assign y1526 = (add_sel & s1526) | (sub_sel & sub1526) | (and_sel & and1526) | (or_sel & or1526);
  assign y1527 = (add_sel & s1527) | (sub_sel & sub1527) | (and_sel & and1527) | (or_sel & or1527);
  assign y1528 = (add_sel & s1528) | (sub_sel & sub1528) | (and_sel & and1528) | (or_sel & or1528);
  assign y1529 = (add_sel & s1529) | (sub_sel & sub1529) | (and_sel & and1529) | (or_sel & or1529);
  assign y1530 = (add_sel & s1530) | (sub_sel & sub1530) | (and_sel & and1530) | (or_sel & or1530);
  assign y1531 = (add_sel & s1531) | (sub_sel & sub1531) | (and_sel & and1531) | (or_sel & or1531);
  assign y1532 = (add_sel & s1532) | (sub_sel & sub1532) | (and_sel & and1532) | (or_sel & or1532);
  assign y1533 = (add_sel & s1533) | (sub_sel & sub1533) | (and_sel & and1533) | (or_sel & or1533);
  assign y1534 = (add_sel & s1534) | (sub_sel & sub1534) | (and_sel & and1534) | (or_sel & or1534);
  assign y1535 = (add_sel & s1535) | (sub_sel & sub1535) | (and_sel & and1535) | (or_sel & or1535);
  assign y1536 = (add_sel & s1536) | (sub_sel & sub1536) | (and_sel & and1536) | (or_sel & or1536);
  assign y1537 = (add_sel & s1537) | (sub_sel & sub1537) | (and_sel & and1537) | (or_sel & or1537);
  assign y1538 = (add_sel & s1538) | (sub_sel & sub1538) | (and_sel & and1538) | (or_sel & or1538);
  assign y1539 = (add_sel & s1539) | (sub_sel & sub1539) | (and_sel & and1539) | (or_sel & or1539);
  assign y1540 = (add_sel & s1540) | (sub_sel & sub1540) | (and_sel & and1540) | (or_sel & or1540);
  assign y1541 = (add_sel & s1541) | (sub_sel & sub1541) | (and_sel & and1541) | (or_sel & or1541);
  assign y1542 = (add_sel & s1542) | (sub_sel & sub1542) | (and_sel & and1542) | (or_sel & or1542);
  assign y1543 = (add_sel & s1543) | (sub_sel & sub1543) | (and_sel & and1543) | (or_sel & or1543);
  assign y1544 = (add_sel & s1544) | (sub_sel & sub1544) | (and_sel & and1544) | (or_sel & or1544);
  assign y1545 = (add_sel & s1545) | (sub_sel & sub1545) | (and_sel & and1545) | (or_sel & or1545);
  assign y1546 = (add_sel & s1546) | (sub_sel & sub1546) | (and_sel & and1546) | (or_sel & or1546);
  assign y1547 = (add_sel & s1547) | (sub_sel & sub1547) | (and_sel & and1547) | (or_sel & or1547);
  assign y1548 = (add_sel & s1548) | (sub_sel & sub1548) | (and_sel & and1548) | (or_sel & or1548);
  assign y1549 = (add_sel & s1549) | (sub_sel & sub1549) | (and_sel & and1549) | (or_sel & or1549);
  assign y1550 = (add_sel & s1550) | (sub_sel & sub1550) | (and_sel & and1550) | (or_sel & or1550);
  assign y1551 = (add_sel & s1551) | (sub_sel & sub1551) | (and_sel & and1551) | (or_sel & or1551);
  assign y1552 = (add_sel & s1552) | (sub_sel & sub1552) | (and_sel & and1552) | (or_sel & or1552);
  assign y1553 = (add_sel & s1553) | (sub_sel & sub1553) | (and_sel & and1553) | (or_sel & or1553);
  assign y1554 = (add_sel & s1554) | (sub_sel & sub1554) | (and_sel & and1554) | (or_sel & or1554);
  assign y1555 = (add_sel & s1555) | (sub_sel & sub1555) | (and_sel & and1555) | (or_sel & or1555);
  assign y1556 = (add_sel & s1556) | (sub_sel & sub1556) | (and_sel & and1556) | (or_sel & or1556);
  assign y1557 = (add_sel & s1557) | (sub_sel & sub1557) | (and_sel & and1557) | (or_sel & or1557);
  assign y1558 = (add_sel & s1558) | (sub_sel & sub1558) | (and_sel & and1558) | (or_sel & or1558);
  assign y1559 = (add_sel & s1559) | (sub_sel & sub1559) | (and_sel & and1559) | (or_sel & or1559);
  assign y1560 = (add_sel & s1560) | (sub_sel & sub1560) | (and_sel & and1560) | (or_sel & or1560);
  assign y1561 = (add_sel & s1561) | (sub_sel & sub1561) | (and_sel & and1561) | (or_sel & or1561);
  assign y1562 = (add_sel & s1562) | (sub_sel & sub1562) | (and_sel & and1562) | (or_sel & or1562);
  assign y1563 = (add_sel & s1563) | (sub_sel & sub1563) | (and_sel & and1563) | (or_sel & or1563);
  assign y1564 = (add_sel & s1564) | (sub_sel & sub1564) | (and_sel & and1564) | (or_sel & or1564);
  assign y1565 = (add_sel & s1565) | (sub_sel & sub1565) | (and_sel & and1565) | (or_sel & or1565);
  assign y1566 = (add_sel & s1566) | (sub_sel & sub1566) | (and_sel & and1566) | (or_sel & or1566);
  assign y1567 = (add_sel & s1567) | (sub_sel & sub1567) | (and_sel & and1567) | (or_sel & or1567);
  assign y1568 = (add_sel & s1568) | (sub_sel & sub1568) | (and_sel & and1568) | (or_sel & or1568);
  assign y1569 = (add_sel & s1569) | (sub_sel & sub1569) | (and_sel & and1569) | (or_sel & or1569);
  assign y1570 = (add_sel & s1570) | (sub_sel & sub1570) | (and_sel & and1570) | (or_sel & or1570);
  assign y1571 = (add_sel & s1571) | (sub_sel & sub1571) | (and_sel & and1571) | (or_sel & or1571);
  assign y1572 = (add_sel & s1572) | (sub_sel & sub1572) | (and_sel & and1572) | (or_sel & or1572);
  assign y1573 = (add_sel & s1573) | (sub_sel & sub1573) | (and_sel & and1573) | (or_sel & or1573);
  assign y1574 = (add_sel & s1574) | (sub_sel & sub1574) | (and_sel & and1574) | (or_sel & or1574);
  assign y1575 = (add_sel & s1575) | (sub_sel & sub1575) | (and_sel & and1575) | (or_sel & or1575);
  assign y1576 = (add_sel & s1576) | (sub_sel & sub1576) | (and_sel & and1576) | (or_sel & or1576);
  assign y1577 = (add_sel & s1577) | (sub_sel & sub1577) | (and_sel & and1577) | (or_sel & or1577);
  assign y1578 = (add_sel & s1578) | (sub_sel & sub1578) | (and_sel & and1578) | (or_sel & or1578);
  assign y1579 = (add_sel & s1579) | (sub_sel & sub1579) | (and_sel & and1579) | (or_sel & or1579);
  assign y1580 = (add_sel & s1580) | (sub_sel & sub1580) | (and_sel & and1580) | (or_sel & or1580);
  assign y1581 = (add_sel & s1581) | (sub_sel & sub1581) | (and_sel & and1581) | (or_sel & or1581);
  assign y1582 = (add_sel & s1582) | (sub_sel & sub1582) | (and_sel & and1582) | (or_sel & or1582);
  assign y1583 = (add_sel & s1583) | (sub_sel & sub1583) | (and_sel & and1583) | (or_sel & or1583);
  assign y1584 = (add_sel & s1584) | (sub_sel & sub1584) | (and_sel & and1584) | (or_sel & or1584);
  assign y1585 = (add_sel & s1585) | (sub_sel & sub1585) | (and_sel & and1585) | (or_sel & or1585);
  assign y1586 = (add_sel & s1586) | (sub_sel & sub1586) | (and_sel & and1586) | (or_sel & or1586);
  assign y1587 = (add_sel & s1587) | (sub_sel & sub1587) | (and_sel & and1587) | (or_sel & or1587);
  assign y1588 = (add_sel & s1588) | (sub_sel & sub1588) | (and_sel & and1588) | (or_sel & or1588);
  assign y1589 = (add_sel & s1589) | (sub_sel & sub1589) | (and_sel & and1589) | (or_sel & or1589);
  assign y1590 = (add_sel & s1590) | (sub_sel & sub1590) | (and_sel & and1590) | (or_sel & or1590);
  assign y1591 = (add_sel & s1591) | (sub_sel & sub1591) | (and_sel & and1591) | (or_sel & or1591);
  assign y1592 = (add_sel & s1592) | (sub_sel & sub1592) | (and_sel & and1592) | (or_sel & or1592);
  assign y1593 = (add_sel & s1593) | (sub_sel & sub1593) | (and_sel & and1593) | (or_sel & or1593);
  assign y1594 = (add_sel & s1594) | (sub_sel & sub1594) | (and_sel & and1594) | (or_sel & or1594);
  assign y1595 = (add_sel & s1595) | (sub_sel & sub1595) | (and_sel & and1595) | (or_sel & or1595);
  assign y1596 = (add_sel & s1596) | (sub_sel & sub1596) | (and_sel & and1596) | (or_sel & or1596);
  assign y1597 = (add_sel & s1597) | (sub_sel & sub1597) | (and_sel & and1597) | (or_sel & or1597);
  assign y1598 = (add_sel & s1598) | (sub_sel & sub1598) | (and_sel & and1598) | (or_sel & or1598);
  assign y1599 = (add_sel & s1599) | (sub_sel & sub1599) | (and_sel & and1599) | (or_sel & or1599);
  assign y1600 = (add_sel & s1600) | (sub_sel & sub1600) | (and_sel & and1600) | (or_sel & or1600);
  assign y1601 = (add_sel & s1601) | (sub_sel & sub1601) | (and_sel & and1601) | (or_sel & or1601);
  assign y1602 = (add_sel & s1602) | (sub_sel & sub1602) | (and_sel & and1602) | (or_sel & or1602);
  assign y1603 = (add_sel & s1603) | (sub_sel & sub1603) | (and_sel & and1603) | (or_sel & or1603);
  assign y1604 = (add_sel & s1604) | (sub_sel & sub1604) | (and_sel & and1604) | (or_sel & or1604);
  assign y1605 = (add_sel & s1605) | (sub_sel & sub1605) | (and_sel & and1605) | (or_sel & or1605);
  assign y1606 = (add_sel & s1606) | (sub_sel & sub1606) | (and_sel & and1606) | (or_sel & or1606);
  assign y1607 = (add_sel & s1607) | (sub_sel & sub1607) | (and_sel & and1607) | (or_sel & or1607);
  assign y1608 = (add_sel & s1608) | (sub_sel & sub1608) | (and_sel & and1608) | (or_sel & or1608);
  assign y1609 = (add_sel & s1609) | (sub_sel & sub1609) | (and_sel & and1609) | (or_sel & or1609);
  assign y1610 = (add_sel & s1610) | (sub_sel & sub1610) | (and_sel & and1610) | (or_sel & or1610);
  assign y1611 = (add_sel & s1611) | (sub_sel & sub1611) | (and_sel & and1611) | (or_sel & or1611);
  assign y1612 = (add_sel & s1612) | (sub_sel & sub1612) | (and_sel & and1612) | (or_sel & or1612);
  assign y1613 = (add_sel & s1613) | (sub_sel & sub1613) | (and_sel & and1613) | (or_sel & or1613);
  assign y1614 = (add_sel & s1614) | (sub_sel & sub1614) | (and_sel & and1614) | (or_sel & or1614);
  assign y1615 = (add_sel & s1615) | (sub_sel & sub1615) | (and_sel & and1615) | (or_sel & or1615);
  assign y1616 = (add_sel & s1616) | (sub_sel & sub1616) | (and_sel & and1616) | (or_sel & or1616);
  assign y1617 = (add_sel & s1617) | (sub_sel & sub1617) | (and_sel & and1617) | (or_sel & or1617);
  assign y1618 = (add_sel & s1618) | (sub_sel & sub1618) | (and_sel & and1618) | (or_sel & or1618);
  assign y1619 = (add_sel & s1619) | (sub_sel & sub1619) | (and_sel & and1619) | (or_sel & or1619);
  assign y1620 = (add_sel & s1620) | (sub_sel & sub1620) | (and_sel & and1620) | (or_sel & or1620);
  assign y1621 = (add_sel & s1621) | (sub_sel & sub1621) | (and_sel & and1621) | (or_sel & or1621);
  assign y1622 = (add_sel & s1622) | (sub_sel & sub1622) | (and_sel & and1622) | (or_sel & or1622);
  assign y1623 = (add_sel & s1623) | (sub_sel & sub1623) | (and_sel & and1623) | (or_sel & or1623);
  assign y1624 = (add_sel & s1624) | (sub_sel & sub1624) | (and_sel & and1624) | (or_sel & or1624);
  assign y1625 = (add_sel & s1625) | (sub_sel & sub1625) | (and_sel & and1625) | (or_sel & or1625);
  assign y1626 = (add_sel & s1626) | (sub_sel & sub1626) | (and_sel & and1626) | (or_sel & or1626);
  assign y1627 = (add_sel & s1627) | (sub_sel & sub1627) | (and_sel & and1627) | (or_sel & or1627);
  assign y1628 = (add_sel & s1628) | (sub_sel & sub1628) | (and_sel & and1628) | (or_sel & or1628);
  assign y1629 = (add_sel & s1629) | (sub_sel & sub1629) | (and_sel & and1629) | (or_sel & or1629);
  assign y1630 = (add_sel & s1630) | (sub_sel & sub1630) | (and_sel & and1630) | (or_sel & or1630);
  assign y1631 = (add_sel & s1631) | (sub_sel & sub1631) | (and_sel & and1631) | (or_sel & or1631);
  assign y1632 = (add_sel & s1632) | (sub_sel & sub1632) | (and_sel & and1632) | (or_sel & or1632);
  assign y1633 = (add_sel & s1633) | (sub_sel & sub1633) | (and_sel & and1633) | (or_sel & or1633);
  assign y1634 = (add_sel & s1634) | (sub_sel & sub1634) | (and_sel & and1634) | (or_sel & or1634);
  assign y1635 = (add_sel & s1635) | (sub_sel & sub1635) | (and_sel & and1635) | (or_sel & or1635);
  assign y1636 = (add_sel & s1636) | (sub_sel & sub1636) | (and_sel & and1636) | (or_sel & or1636);
  assign y1637 = (add_sel & s1637) | (sub_sel & sub1637) | (and_sel & and1637) | (or_sel & or1637);
  assign y1638 = (add_sel & s1638) | (sub_sel & sub1638) | (and_sel & and1638) | (or_sel & or1638);
  assign y1639 = (add_sel & s1639) | (sub_sel & sub1639) | (and_sel & and1639) | (or_sel & or1639);
  assign y1640 = (add_sel & s1640) | (sub_sel & sub1640) | (and_sel & and1640) | (or_sel & or1640);
  assign y1641 = (add_sel & s1641) | (sub_sel & sub1641) | (and_sel & and1641) | (or_sel & or1641);
  assign y1642 = (add_sel & s1642) | (sub_sel & sub1642) | (and_sel & and1642) | (or_sel & or1642);
  assign y1643 = (add_sel & s1643) | (sub_sel & sub1643) | (and_sel & and1643) | (or_sel & or1643);
  assign y1644 = (add_sel & s1644) | (sub_sel & sub1644) | (and_sel & and1644) | (or_sel & or1644);
  assign y1645 = (add_sel & s1645) | (sub_sel & sub1645) | (and_sel & and1645) | (or_sel & or1645);
  assign y1646 = (add_sel & s1646) | (sub_sel & sub1646) | (and_sel & and1646) | (or_sel & or1646);
  assign y1647 = (add_sel & s1647) | (sub_sel & sub1647) | (and_sel & and1647) | (or_sel & or1647);
  assign y1648 = (add_sel & s1648) | (sub_sel & sub1648) | (and_sel & and1648) | (or_sel & or1648);
  assign y1649 = (add_sel & s1649) | (sub_sel & sub1649) | (and_sel & and1649) | (or_sel & or1649);
  assign y1650 = (add_sel & s1650) | (sub_sel & sub1650) | (and_sel & and1650) | (or_sel & or1650);
  assign y1651 = (add_sel & s1651) | (sub_sel & sub1651) | (and_sel & and1651) | (or_sel & or1651);
  assign y1652 = (add_sel & s1652) | (sub_sel & sub1652) | (and_sel & and1652) | (or_sel & or1652);
  assign y1653 = (add_sel & s1653) | (sub_sel & sub1653) | (and_sel & and1653) | (or_sel & or1653);
  assign y1654 = (add_sel & s1654) | (sub_sel & sub1654) | (and_sel & and1654) | (or_sel & or1654);
  assign y1655 = (add_sel & s1655) | (sub_sel & sub1655) | (and_sel & and1655) | (or_sel & or1655);
  assign y1656 = (add_sel & s1656) | (sub_sel & sub1656) | (and_sel & and1656) | (or_sel & or1656);
  assign y1657 = (add_sel & s1657) | (sub_sel & sub1657) | (and_sel & and1657) | (or_sel & or1657);
  assign y1658 = (add_sel & s1658) | (sub_sel & sub1658) | (and_sel & and1658) | (or_sel & or1658);
  assign y1659 = (add_sel & s1659) | (sub_sel & sub1659) | (and_sel & and1659) | (or_sel & or1659);
  assign y1660 = (add_sel & s1660) | (sub_sel & sub1660) | (and_sel & and1660) | (or_sel & or1660);
  assign y1661 = (add_sel & s1661) | (sub_sel & sub1661) | (and_sel & and1661) | (or_sel & or1661);
  assign y1662 = (add_sel & s1662) | (sub_sel & sub1662) | (and_sel & and1662) | (or_sel & or1662);
  assign y1663 = (add_sel & s1663) | (sub_sel & sub1663) | (and_sel & and1663) | (or_sel & or1663);
  assign y1664 = (add_sel & s1664) | (sub_sel & sub1664) | (and_sel & and1664) | (or_sel & or1664);
  assign y1665 = (add_sel & s1665) | (sub_sel & sub1665) | (and_sel & and1665) | (or_sel & or1665);
  assign y1666 = (add_sel & s1666) | (sub_sel & sub1666) | (and_sel & and1666) | (or_sel & or1666);
  assign y1667 = (add_sel & s1667) | (sub_sel & sub1667) | (and_sel & and1667) | (or_sel & or1667);
  assign y1668 = (add_sel & s1668) | (sub_sel & sub1668) | (and_sel & and1668) | (or_sel & or1668);
  assign y1669 = (add_sel & s1669) | (sub_sel & sub1669) | (and_sel & and1669) | (or_sel & or1669);
  assign y1670 = (add_sel & s1670) | (sub_sel & sub1670) | (and_sel & and1670) | (or_sel & or1670);
  assign y1671 = (add_sel & s1671) | (sub_sel & sub1671) | (and_sel & and1671) | (or_sel & or1671);
  assign y1672 = (add_sel & s1672) | (sub_sel & sub1672) | (and_sel & and1672) | (or_sel & or1672);
  assign y1673 = (add_sel & s1673) | (sub_sel & sub1673) | (and_sel & and1673) | (or_sel & or1673);
  assign y1674 = (add_sel & s1674) | (sub_sel & sub1674) | (and_sel & and1674) | (or_sel & or1674);
  assign y1675 = (add_sel & s1675) | (sub_sel & sub1675) | (and_sel & and1675) | (or_sel & or1675);
  assign y1676 = (add_sel & s1676) | (sub_sel & sub1676) | (and_sel & and1676) | (or_sel & or1676);
  assign y1677 = (add_sel & s1677) | (sub_sel & sub1677) | (and_sel & and1677) | (or_sel & or1677);
  assign y1678 = (add_sel & s1678) | (sub_sel & sub1678) | (and_sel & and1678) | (or_sel & or1678);
  assign y1679 = (add_sel & s1679) | (sub_sel & sub1679) | (and_sel & and1679) | (or_sel & or1679);
  assign y1680 = (add_sel & s1680) | (sub_sel & sub1680) | (and_sel & and1680) | (or_sel & or1680);
  assign y1681 = (add_sel & s1681) | (sub_sel & sub1681) | (and_sel & and1681) | (or_sel & or1681);
  assign y1682 = (add_sel & s1682) | (sub_sel & sub1682) | (and_sel & and1682) | (or_sel & or1682);
  assign y1683 = (add_sel & s1683) | (sub_sel & sub1683) | (and_sel & and1683) | (or_sel & or1683);
  assign y1684 = (add_sel & s1684) | (sub_sel & sub1684) | (and_sel & and1684) | (or_sel & or1684);
  assign y1685 = (add_sel & s1685) | (sub_sel & sub1685) | (and_sel & and1685) | (or_sel & or1685);
  assign y1686 = (add_sel & s1686) | (sub_sel & sub1686) | (and_sel & and1686) | (or_sel & or1686);
  assign y1687 = (add_sel & s1687) | (sub_sel & sub1687) | (and_sel & and1687) | (or_sel & or1687);
  assign y1688 = (add_sel & s1688) | (sub_sel & sub1688) | (and_sel & and1688) | (or_sel & or1688);
  assign y1689 = (add_sel & s1689) | (sub_sel & sub1689) | (and_sel & and1689) | (or_sel & or1689);
  assign y1690 = (add_sel & s1690) | (sub_sel & sub1690) | (and_sel & and1690) | (or_sel & or1690);
  assign y1691 = (add_sel & s1691) | (sub_sel & sub1691) | (and_sel & and1691) | (or_sel & or1691);
  assign y1692 = (add_sel & s1692) | (sub_sel & sub1692) | (and_sel & and1692) | (or_sel & or1692);
  assign y1693 = (add_sel & s1693) | (sub_sel & sub1693) | (and_sel & and1693) | (or_sel & or1693);
  assign y1694 = (add_sel & s1694) | (sub_sel & sub1694) | (and_sel & and1694) | (or_sel & or1694);
  assign y1695 = (add_sel & s1695) | (sub_sel & sub1695) | (and_sel & and1695) | (or_sel & or1695);
  assign y1696 = (add_sel & s1696) | (sub_sel & sub1696) | (and_sel & and1696) | (or_sel & or1696);
  assign y1697 = (add_sel & s1697) | (sub_sel & sub1697) | (and_sel & and1697) | (or_sel & or1697);
  assign y1698 = (add_sel & s1698) | (sub_sel & sub1698) | (and_sel & and1698) | (or_sel & or1698);
  assign y1699 = (add_sel & s1699) | (sub_sel & sub1699) | (and_sel & and1699) | (or_sel & or1699);
  assign y1700 = (add_sel & s1700) | (sub_sel & sub1700) | (and_sel & and1700) | (or_sel & or1700);
  assign y1701 = (add_sel & s1701) | (sub_sel & sub1701) | (and_sel & and1701) | (or_sel & or1701);
  assign y1702 = (add_sel & s1702) | (sub_sel & sub1702) | (and_sel & and1702) | (or_sel & or1702);
  assign y1703 = (add_sel & s1703) | (sub_sel & sub1703) | (and_sel & and1703) | (or_sel & or1703);
  assign y1704 = (add_sel & s1704) | (sub_sel & sub1704) | (and_sel & and1704) | (or_sel & or1704);
  assign y1705 = (add_sel & s1705) | (sub_sel & sub1705) | (and_sel & and1705) | (or_sel & or1705);
  assign y1706 = (add_sel & s1706) | (sub_sel & sub1706) | (and_sel & and1706) | (or_sel & or1706);
  assign y1707 = (add_sel & s1707) | (sub_sel & sub1707) | (and_sel & and1707) | (or_sel & or1707);
  assign y1708 = (add_sel & s1708) | (sub_sel & sub1708) | (and_sel & and1708) | (or_sel & or1708);
  assign y1709 = (add_sel & s1709) | (sub_sel & sub1709) | (and_sel & and1709) | (or_sel & or1709);
  assign y1710 = (add_sel & s1710) | (sub_sel & sub1710) | (and_sel & and1710) | (or_sel & or1710);
  assign y1711 = (add_sel & s1711) | (sub_sel & sub1711) | (and_sel & and1711) | (or_sel & or1711);
  assign y1712 = (add_sel & s1712) | (sub_sel & sub1712) | (and_sel & and1712) | (or_sel & or1712);
  assign y1713 = (add_sel & s1713) | (sub_sel & sub1713) | (and_sel & and1713) | (or_sel & or1713);
  assign y1714 = (add_sel & s1714) | (sub_sel & sub1714) | (and_sel & and1714) | (or_sel & or1714);
  assign y1715 = (add_sel & s1715) | (sub_sel & sub1715) | (and_sel & and1715) | (or_sel & or1715);
  assign y1716 = (add_sel & s1716) | (sub_sel & sub1716) | (and_sel & and1716) | (or_sel & or1716);
  assign y1717 = (add_sel & s1717) | (sub_sel & sub1717) | (and_sel & and1717) | (or_sel & or1717);
  assign y1718 = (add_sel & s1718) | (sub_sel & sub1718) | (and_sel & and1718) | (or_sel & or1718);
  assign y1719 = (add_sel & s1719) | (sub_sel & sub1719) | (and_sel & and1719) | (or_sel & or1719);
  assign y1720 = (add_sel & s1720) | (sub_sel & sub1720) | (and_sel & and1720) | (or_sel & or1720);
  assign y1721 = (add_sel & s1721) | (sub_sel & sub1721) | (and_sel & and1721) | (or_sel & or1721);
  assign y1722 = (add_sel & s1722) | (sub_sel & sub1722) | (and_sel & and1722) | (or_sel & or1722);
  assign y1723 = (add_sel & s1723) | (sub_sel & sub1723) | (and_sel & and1723) | (or_sel & or1723);
  assign y1724 = (add_sel & s1724) | (sub_sel & sub1724) | (and_sel & and1724) | (or_sel & or1724);
  assign y1725 = (add_sel & s1725) | (sub_sel & sub1725) | (and_sel & and1725) | (or_sel & or1725);
  assign y1726 = (add_sel & s1726) | (sub_sel & sub1726) | (and_sel & and1726) | (or_sel & or1726);
  assign y1727 = (add_sel & s1727) | (sub_sel & sub1727) | (and_sel & and1727) | (or_sel & or1727);
  assign y1728 = (add_sel & s1728) | (sub_sel & sub1728) | (and_sel & and1728) | (or_sel & or1728);
  assign y1729 = (add_sel & s1729) | (sub_sel & sub1729) | (and_sel & and1729) | (or_sel & or1729);
  assign y1730 = (add_sel & s1730) | (sub_sel & sub1730) | (and_sel & and1730) | (or_sel & or1730);
  assign y1731 = (add_sel & s1731) | (sub_sel & sub1731) | (and_sel & and1731) | (or_sel & or1731);
  assign y1732 = (add_sel & s1732) | (sub_sel & sub1732) | (and_sel & and1732) | (or_sel & or1732);
  assign y1733 = (add_sel & s1733) | (sub_sel & sub1733) | (and_sel & and1733) | (or_sel & or1733);
  assign y1734 = (add_sel & s1734) | (sub_sel & sub1734) | (and_sel & and1734) | (or_sel & or1734);
  assign y1735 = (add_sel & s1735) | (sub_sel & sub1735) | (and_sel & and1735) | (or_sel & or1735);
  assign y1736 = (add_sel & s1736) | (sub_sel & sub1736) | (and_sel & and1736) | (or_sel & or1736);
  assign y1737 = (add_sel & s1737) | (sub_sel & sub1737) | (and_sel & and1737) | (or_sel & or1737);
  assign y1738 = (add_sel & s1738) | (sub_sel & sub1738) | (and_sel & and1738) | (or_sel & or1738);
  assign y1739 = (add_sel & s1739) | (sub_sel & sub1739) | (and_sel & and1739) | (or_sel & or1739);
  assign y1740 = (add_sel & s1740) | (sub_sel & sub1740) | (and_sel & and1740) | (or_sel & or1740);
  assign y1741 = (add_sel & s1741) | (sub_sel & sub1741) | (and_sel & and1741) | (or_sel & or1741);
  assign y1742 = (add_sel & s1742) | (sub_sel & sub1742) | (and_sel & and1742) | (or_sel & or1742);
  assign y1743 = (add_sel & s1743) | (sub_sel & sub1743) | (and_sel & and1743) | (or_sel & or1743);
  assign y1744 = (add_sel & s1744) | (sub_sel & sub1744) | (and_sel & and1744) | (or_sel & or1744);
  assign y1745 = (add_sel & s1745) | (sub_sel & sub1745) | (and_sel & and1745) | (or_sel & or1745);
  assign y1746 = (add_sel & s1746) | (sub_sel & sub1746) | (and_sel & and1746) | (or_sel & or1746);
  assign y1747 = (add_sel & s1747) | (sub_sel & sub1747) | (and_sel & and1747) | (or_sel & or1747);
  assign y1748 = (add_sel & s1748) | (sub_sel & sub1748) | (and_sel & and1748) | (or_sel & or1748);
  assign y1749 = (add_sel & s1749) | (sub_sel & sub1749) | (and_sel & and1749) | (or_sel & or1749);
  assign y1750 = (add_sel & s1750) | (sub_sel & sub1750) | (and_sel & and1750) | (or_sel & or1750);
  assign y1751 = (add_sel & s1751) | (sub_sel & sub1751) | (and_sel & and1751) | (or_sel & or1751);
  assign y1752 = (add_sel & s1752) | (sub_sel & sub1752) | (and_sel & and1752) | (or_sel & or1752);
  assign y1753 = (add_sel & s1753) | (sub_sel & sub1753) | (and_sel & and1753) | (or_sel & or1753);
  assign y1754 = (add_sel & s1754) | (sub_sel & sub1754) | (and_sel & and1754) | (or_sel & or1754);
  assign y1755 = (add_sel & s1755) | (sub_sel & sub1755) | (and_sel & and1755) | (or_sel & or1755);
  assign y1756 = (add_sel & s1756) | (sub_sel & sub1756) | (and_sel & and1756) | (or_sel & or1756);
  assign y1757 = (add_sel & s1757) | (sub_sel & sub1757) | (and_sel & and1757) | (or_sel & or1757);
  assign y1758 = (add_sel & s1758) | (sub_sel & sub1758) | (and_sel & and1758) | (or_sel & or1758);
  assign y1759 = (add_sel & s1759) | (sub_sel & sub1759) | (and_sel & and1759) | (or_sel & or1759);
  assign y1760 = (add_sel & s1760) | (sub_sel & sub1760) | (and_sel & and1760) | (or_sel & or1760);
  assign y1761 = (add_sel & s1761) | (sub_sel & sub1761) | (and_sel & and1761) | (or_sel & or1761);
  assign y1762 = (add_sel & s1762) | (sub_sel & sub1762) | (and_sel & and1762) | (or_sel & or1762);
  assign y1763 = (add_sel & s1763) | (sub_sel & sub1763) | (and_sel & and1763) | (or_sel & or1763);
  assign y1764 = (add_sel & s1764) | (sub_sel & sub1764) | (and_sel & and1764) | (or_sel & or1764);
  assign y1765 = (add_sel & s1765) | (sub_sel & sub1765) | (and_sel & and1765) | (or_sel & or1765);
  assign y1766 = (add_sel & s1766) | (sub_sel & sub1766) | (and_sel & and1766) | (or_sel & or1766);
  assign y1767 = (add_sel & s1767) | (sub_sel & sub1767) | (and_sel & and1767) | (or_sel & or1767);
  assign y1768 = (add_sel & s1768) | (sub_sel & sub1768) | (and_sel & and1768) | (or_sel & or1768);
  assign y1769 = (add_sel & s1769) | (sub_sel & sub1769) | (and_sel & and1769) | (or_sel & or1769);
  assign y1770 = (add_sel & s1770) | (sub_sel & sub1770) | (and_sel & and1770) | (or_sel & or1770);
  assign y1771 = (add_sel & s1771) | (sub_sel & sub1771) | (and_sel & and1771) | (or_sel & or1771);
  assign y1772 = (add_sel & s1772) | (sub_sel & sub1772) | (and_sel & and1772) | (or_sel & or1772);
  assign y1773 = (add_sel & s1773) | (sub_sel & sub1773) | (and_sel & and1773) | (or_sel & or1773);
  assign y1774 = (add_sel & s1774) | (sub_sel & sub1774) | (and_sel & and1774) | (or_sel & or1774);
  assign y1775 = (add_sel & s1775) | (sub_sel & sub1775) | (and_sel & and1775) | (or_sel & or1775);
  assign y1776 = (add_sel & s1776) | (sub_sel & sub1776) | (and_sel & and1776) | (or_sel & or1776);
  assign y1777 = (add_sel & s1777) | (sub_sel & sub1777) | (and_sel & and1777) | (or_sel & or1777);
  assign y1778 = (add_sel & s1778) | (sub_sel & sub1778) | (and_sel & and1778) | (or_sel & or1778);
  assign y1779 = (add_sel & s1779) | (sub_sel & sub1779) | (and_sel & and1779) | (or_sel & or1779);
  assign y1780 = (add_sel & s1780) | (sub_sel & sub1780) | (and_sel & and1780) | (or_sel & or1780);
  assign y1781 = (add_sel & s1781) | (sub_sel & sub1781) | (and_sel & and1781) | (or_sel & or1781);
  assign y1782 = (add_sel & s1782) | (sub_sel & sub1782) | (and_sel & and1782) | (or_sel & or1782);
  assign y1783 = (add_sel & s1783) | (sub_sel & sub1783) | (and_sel & and1783) | (or_sel & or1783);
  assign y1784 = (add_sel & s1784) | (sub_sel & sub1784) | (and_sel & and1784) | (or_sel & or1784);
  assign y1785 = (add_sel & s1785) | (sub_sel & sub1785) | (and_sel & and1785) | (or_sel & or1785);
  assign y1786 = (add_sel & s1786) | (sub_sel & sub1786) | (and_sel & and1786) | (or_sel & or1786);
  assign y1787 = (add_sel & s1787) | (sub_sel & sub1787) | (and_sel & and1787) | (or_sel & or1787);
  assign y1788 = (add_sel & s1788) | (sub_sel & sub1788) | (and_sel & and1788) | (or_sel & or1788);
  assign y1789 = (add_sel & s1789) | (sub_sel & sub1789) | (and_sel & and1789) | (or_sel & or1789);
  assign y1790 = (add_sel & s1790) | (sub_sel & sub1790) | (and_sel & and1790) | (or_sel & or1790);
  assign y1791 = (add_sel & s1791) | (sub_sel & sub1791) | (and_sel & and1791) | (or_sel & or1791);
  assign y1792 = (add_sel & s1792) | (sub_sel & sub1792) | (and_sel & and1792) | (or_sel & or1792);
  assign y1793 = (add_sel & s1793) | (sub_sel & sub1793) | (and_sel & and1793) | (or_sel & or1793);
  assign y1794 = (add_sel & s1794) | (sub_sel & sub1794) | (and_sel & and1794) | (or_sel & or1794);
  assign y1795 = (add_sel & s1795) | (sub_sel & sub1795) | (and_sel & and1795) | (or_sel & or1795);
  assign y1796 = (add_sel & s1796) | (sub_sel & sub1796) | (and_sel & and1796) | (or_sel & or1796);
  assign y1797 = (add_sel & s1797) | (sub_sel & sub1797) | (and_sel & and1797) | (or_sel & or1797);
  assign y1798 = (add_sel & s1798) | (sub_sel & sub1798) | (and_sel & and1798) | (or_sel & or1798);
  assign y1799 = (add_sel & s1799) | (sub_sel & sub1799) | (and_sel & and1799) | (or_sel & or1799);
  assign y1800 = (add_sel & s1800) | (sub_sel & sub1800) | (and_sel & and1800) | (or_sel & or1800);
  assign y1801 = (add_sel & s1801) | (sub_sel & sub1801) | (and_sel & and1801) | (or_sel & or1801);
  assign y1802 = (add_sel & s1802) | (sub_sel & sub1802) | (and_sel & and1802) | (or_sel & or1802);
  assign y1803 = (add_sel & s1803) | (sub_sel & sub1803) | (and_sel & and1803) | (or_sel & or1803);
  assign y1804 = (add_sel & s1804) | (sub_sel & sub1804) | (and_sel & and1804) | (or_sel & or1804);
  assign y1805 = (add_sel & s1805) | (sub_sel & sub1805) | (and_sel & and1805) | (or_sel & or1805);
  assign y1806 = (add_sel & s1806) | (sub_sel & sub1806) | (and_sel & and1806) | (or_sel & or1806);
  assign y1807 = (add_sel & s1807) | (sub_sel & sub1807) | (and_sel & and1807) | (or_sel & or1807);
  assign y1808 = (add_sel & s1808) | (sub_sel & sub1808) | (and_sel & and1808) | (or_sel & or1808);
  assign y1809 = (add_sel & s1809) | (sub_sel & sub1809) | (and_sel & and1809) | (or_sel & or1809);
  assign y1810 = (add_sel & s1810) | (sub_sel & sub1810) | (and_sel & and1810) | (or_sel & or1810);
  assign y1811 = (add_sel & s1811) | (sub_sel & sub1811) | (and_sel & and1811) | (or_sel & or1811);
  assign y1812 = (add_sel & s1812) | (sub_sel & sub1812) | (and_sel & and1812) | (or_sel & or1812);
  assign y1813 = (add_sel & s1813) | (sub_sel & sub1813) | (and_sel & and1813) | (or_sel & or1813);
  assign y1814 = (add_sel & s1814) | (sub_sel & sub1814) | (and_sel & and1814) | (or_sel & or1814);
  assign y1815 = (add_sel & s1815) | (sub_sel & sub1815) | (and_sel & and1815) | (or_sel & or1815);
  assign y1816 = (add_sel & s1816) | (sub_sel & sub1816) | (and_sel & and1816) | (or_sel & or1816);
  assign y1817 = (add_sel & s1817) | (sub_sel & sub1817) | (and_sel & and1817) | (or_sel & or1817);
  assign y1818 = (add_sel & s1818) | (sub_sel & sub1818) | (and_sel & and1818) | (or_sel & or1818);
  assign y1819 = (add_sel & s1819) | (sub_sel & sub1819) | (and_sel & and1819) | (or_sel & or1819);
  assign y1820 = (add_sel & s1820) | (sub_sel & sub1820) | (and_sel & and1820) | (or_sel & or1820);
  assign y1821 = (add_sel & s1821) | (sub_sel & sub1821) | (and_sel & and1821) | (or_sel & or1821);
  assign y1822 = (add_sel & s1822) | (sub_sel & sub1822) | (and_sel & and1822) | (or_sel & or1822);
  assign y1823 = (add_sel & s1823) | (sub_sel & sub1823) | (and_sel & and1823) | (or_sel & or1823);
  assign y1824 = (add_sel & s1824) | (sub_sel & sub1824) | (and_sel & and1824) | (or_sel & or1824);
  assign y1825 = (add_sel & s1825) | (sub_sel & sub1825) | (and_sel & and1825) | (or_sel & or1825);
  assign y1826 = (add_sel & s1826) | (sub_sel & sub1826) | (and_sel & and1826) | (or_sel & or1826);
  assign y1827 = (add_sel & s1827) | (sub_sel & sub1827) | (and_sel & and1827) | (or_sel & or1827);
  assign y1828 = (add_sel & s1828) | (sub_sel & sub1828) | (and_sel & and1828) | (or_sel & or1828);
  assign y1829 = (add_sel & s1829) | (sub_sel & sub1829) | (and_sel & and1829) | (or_sel & or1829);
  assign y1830 = (add_sel & s1830) | (sub_sel & sub1830) | (and_sel & and1830) | (or_sel & or1830);
  assign y1831 = (add_sel & s1831) | (sub_sel & sub1831) | (and_sel & and1831) | (or_sel & or1831);
  assign y1832 = (add_sel & s1832) | (sub_sel & sub1832) | (and_sel & and1832) | (or_sel & or1832);
  assign y1833 = (add_sel & s1833) | (sub_sel & sub1833) | (and_sel & and1833) | (or_sel & or1833);
  assign y1834 = (add_sel & s1834) | (sub_sel & sub1834) | (and_sel & and1834) | (or_sel & or1834);
  assign y1835 = (add_sel & s1835) | (sub_sel & sub1835) | (and_sel & and1835) | (or_sel & or1835);
  assign y1836 = (add_sel & s1836) | (sub_sel & sub1836) | (and_sel & and1836) | (or_sel & or1836);
  assign y1837 = (add_sel & s1837) | (sub_sel & sub1837) | (and_sel & and1837) | (or_sel & or1837);
  assign y1838 = (add_sel & s1838) | (sub_sel & sub1838) | (and_sel & and1838) | (or_sel & or1838);
  assign y1839 = (add_sel & s1839) | (sub_sel & sub1839) | (and_sel & and1839) | (or_sel & or1839);
  assign y1840 = (add_sel & s1840) | (sub_sel & sub1840) | (and_sel & and1840) | (or_sel & or1840);
  assign y1841 = (add_sel & s1841) | (sub_sel & sub1841) | (and_sel & and1841) | (or_sel & or1841);
  assign y1842 = (add_sel & s1842) | (sub_sel & sub1842) | (and_sel & and1842) | (or_sel & or1842);
  assign y1843 = (add_sel & s1843) | (sub_sel & sub1843) | (and_sel & and1843) | (or_sel & or1843);
  assign y1844 = (add_sel & s1844) | (sub_sel & sub1844) | (and_sel & and1844) | (or_sel & or1844);
  assign y1845 = (add_sel & s1845) | (sub_sel & sub1845) | (and_sel & and1845) | (or_sel & or1845);
  assign y1846 = (add_sel & s1846) | (sub_sel & sub1846) | (and_sel & and1846) | (or_sel & or1846);
  assign y1847 = (add_sel & s1847) | (sub_sel & sub1847) | (and_sel & and1847) | (or_sel & or1847);
  assign y1848 = (add_sel & s1848) | (sub_sel & sub1848) | (and_sel & and1848) | (or_sel & or1848);
  assign y1849 = (add_sel & s1849) | (sub_sel & sub1849) | (and_sel & and1849) | (or_sel & or1849);
  assign y1850 = (add_sel & s1850) | (sub_sel & sub1850) | (and_sel & and1850) | (or_sel & or1850);
  assign y1851 = (add_sel & s1851) | (sub_sel & sub1851) | (and_sel & and1851) | (or_sel & or1851);
  assign y1852 = (add_sel & s1852) | (sub_sel & sub1852) | (and_sel & and1852) | (or_sel & or1852);
  assign y1853 = (add_sel & s1853) | (sub_sel & sub1853) | (and_sel & and1853) | (or_sel & or1853);
  assign y1854 = (add_sel & s1854) | (sub_sel & sub1854) | (and_sel & and1854) | (or_sel & or1854);
  assign y1855 = (add_sel & s1855) | (sub_sel & sub1855) | (and_sel & and1855) | (or_sel & or1855);
  assign y1856 = (add_sel & s1856) | (sub_sel & sub1856) | (and_sel & and1856) | (or_sel & or1856);
  assign y1857 = (add_sel & s1857) | (sub_sel & sub1857) | (and_sel & and1857) | (or_sel & or1857);
  assign y1858 = (add_sel & s1858) | (sub_sel & sub1858) | (and_sel & and1858) | (or_sel & or1858);
  assign y1859 = (add_sel & s1859) | (sub_sel & sub1859) | (and_sel & and1859) | (or_sel & or1859);
  assign y1860 = (add_sel & s1860) | (sub_sel & sub1860) | (and_sel & and1860) | (or_sel & or1860);
  assign y1861 = (add_sel & s1861) | (sub_sel & sub1861) | (and_sel & and1861) | (or_sel & or1861);
  assign y1862 = (add_sel & s1862) | (sub_sel & sub1862) | (and_sel & and1862) | (or_sel & or1862);
  assign y1863 = (add_sel & s1863) | (sub_sel & sub1863) | (and_sel & and1863) | (or_sel & or1863);
  assign y1864 = (add_sel & s1864) | (sub_sel & sub1864) | (and_sel & and1864) | (or_sel & or1864);
  assign y1865 = (add_sel & s1865) | (sub_sel & sub1865) | (and_sel & and1865) | (or_sel & or1865);
  assign y1866 = (add_sel & s1866) | (sub_sel & sub1866) | (and_sel & and1866) | (or_sel & or1866);
  assign y1867 = (add_sel & s1867) | (sub_sel & sub1867) | (and_sel & and1867) | (or_sel & or1867);
  assign y1868 = (add_sel & s1868) | (sub_sel & sub1868) | (and_sel & and1868) | (or_sel & or1868);
  assign y1869 = (add_sel & s1869) | (sub_sel & sub1869) | (and_sel & and1869) | (or_sel & or1869);
  assign y1870 = (add_sel & s1870) | (sub_sel & sub1870) | (and_sel & and1870) | (or_sel & or1870);
  assign y1871 = (add_sel & s1871) | (sub_sel & sub1871) | (and_sel & and1871) | (or_sel & or1871);
  assign y1872 = (add_sel & s1872) | (sub_sel & sub1872) | (and_sel & and1872) | (or_sel & or1872);
  assign y1873 = (add_sel & s1873) | (sub_sel & sub1873) | (and_sel & and1873) | (or_sel & or1873);
  assign y1874 = (add_sel & s1874) | (sub_sel & sub1874) | (and_sel & and1874) | (or_sel & or1874);
  assign y1875 = (add_sel & s1875) | (sub_sel & sub1875) | (and_sel & and1875) | (or_sel & or1875);
  assign y1876 = (add_sel & s1876) | (sub_sel & sub1876) | (and_sel & and1876) | (or_sel & or1876);
  assign y1877 = (add_sel & s1877) | (sub_sel & sub1877) | (and_sel & and1877) | (or_sel & or1877);
  assign y1878 = (add_sel & s1878) | (sub_sel & sub1878) | (and_sel & and1878) | (or_sel & or1878);
  assign y1879 = (add_sel & s1879) | (sub_sel & sub1879) | (and_sel & and1879) | (or_sel & or1879);
  assign y1880 = (add_sel & s1880) | (sub_sel & sub1880) | (and_sel & and1880) | (or_sel & or1880);
  assign y1881 = (add_sel & s1881) | (sub_sel & sub1881) | (and_sel & and1881) | (or_sel & or1881);
  assign y1882 = (add_sel & s1882) | (sub_sel & sub1882) | (and_sel & and1882) | (or_sel & or1882);
  assign y1883 = (add_sel & s1883) | (sub_sel & sub1883) | (and_sel & and1883) | (or_sel & or1883);
  assign y1884 = (add_sel & s1884) | (sub_sel & sub1884) | (and_sel & and1884) | (or_sel & or1884);
  assign y1885 = (add_sel & s1885) | (sub_sel & sub1885) | (and_sel & and1885) | (or_sel & or1885);
  assign y1886 = (add_sel & s1886) | (sub_sel & sub1886) | (and_sel & and1886) | (or_sel & or1886);
  assign y1887 = (add_sel & s1887) | (sub_sel & sub1887) | (and_sel & and1887) | (or_sel & or1887);
  assign y1888 = (add_sel & s1888) | (sub_sel & sub1888) | (and_sel & and1888) | (or_sel & or1888);
  assign y1889 = (add_sel & s1889) | (sub_sel & sub1889) | (and_sel & and1889) | (or_sel & or1889);
  assign y1890 = (add_sel & s1890) | (sub_sel & sub1890) | (and_sel & and1890) | (or_sel & or1890);
  assign y1891 = (add_sel & s1891) | (sub_sel & sub1891) | (and_sel & and1891) | (or_sel & or1891);
  assign y1892 = (add_sel & s1892) | (sub_sel & sub1892) | (and_sel & and1892) | (or_sel & or1892);
  assign y1893 = (add_sel & s1893) | (sub_sel & sub1893) | (and_sel & and1893) | (or_sel & or1893);
  assign y1894 = (add_sel & s1894) | (sub_sel & sub1894) | (and_sel & and1894) | (or_sel & or1894);
  assign y1895 = (add_sel & s1895) | (sub_sel & sub1895) | (and_sel & and1895) | (or_sel & or1895);
  assign y1896 = (add_sel & s1896) | (sub_sel & sub1896) | (and_sel & and1896) | (or_sel & or1896);
  assign y1897 = (add_sel & s1897) | (sub_sel & sub1897) | (and_sel & and1897) | (or_sel & or1897);
  assign y1898 = (add_sel & s1898) | (sub_sel & sub1898) | (and_sel & and1898) | (or_sel & or1898);
  assign y1899 = (add_sel & s1899) | (sub_sel & sub1899) | (and_sel & and1899) | (or_sel & or1899);
  assign y1900 = (add_sel & s1900) | (sub_sel & sub1900) | (and_sel & and1900) | (or_sel & or1900);
  assign y1901 = (add_sel & s1901) | (sub_sel & sub1901) | (and_sel & and1901) | (or_sel & or1901);
  assign y1902 = (add_sel & s1902) | (sub_sel & sub1902) | (and_sel & and1902) | (or_sel & or1902);
  assign y1903 = (add_sel & s1903) | (sub_sel & sub1903) | (and_sel & and1903) | (or_sel & or1903);
  assign y1904 = (add_sel & s1904) | (sub_sel & sub1904) | (and_sel & and1904) | (or_sel & or1904);
  assign y1905 = (add_sel & s1905) | (sub_sel & sub1905) | (and_sel & and1905) | (or_sel & or1905);
  assign y1906 = (add_sel & s1906) | (sub_sel & sub1906) | (and_sel & and1906) | (or_sel & or1906);
  assign y1907 = (add_sel & s1907) | (sub_sel & sub1907) | (and_sel & and1907) | (or_sel & or1907);
  assign y1908 = (add_sel & s1908) | (sub_sel & sub1908) | (and_sel & and1908) | (or_sel & or1908);
  assign y1909 = (add_sel & s1909) | (sub_sel & sub1909) | (and_sel & and1909) | (or_sel & or1909);
  assign y1910 = (add_sel & s1910) | (sub_sel & sub1910) | (and_sel & and1910) | (or_sel & or1910);
  assign y1911 = (add_sel & s1911) | (sub_sel & sub1911) | (and_sel & and1911) | (or_sel & or1911);
  assign y1912 = (add_sel & s1912) | (sub_sel & sub1912) | (and_sel & and1912) | (or_sel & or1912);
  assign y1913 = (add_sel & s1913) | (sub_sel & sub1913) | (and_sel & and1913) | (or_sel & or1913);
  assign y1914 = (add_sel & s1914) | (sub_sel & sub1914) | (and_sel & and1914) | (or_sel & or1914);
  assign y1915 = (add_sel & s1915) | (sub_sel & sub1915) | (and_sel & and1915) | (or_sel & or1915);
  assign y1916 = (add_sel & s1916) | (sub_sel & sub1916) | (and_sel & and1916) | (or_sel & or1916);
  assign y1917 = (add_sel & s1917) | (sub_sel & sub1917) | (and_sel & and1917) | (or_sel & or1917);
  assign y1918 = (add_sel & s1918) | (sub_sel & sub1918) | (and_sel & and1918) | (or_sel & or1918);
  assign y1919 = (add_sel & s1919) | (sub_sel & sub1919) | (and_sel & and1919) | (or_sel & or1919);
  assign y1920 = (add_sel & s1920) | (sub_sel & sub1920) | (and_sel & and1920) | (or_sel & or1920);
  assign y1921 = (add_sel & s1921) | (sub_sel & sub1921) | (and_sel & and1921) | (or_sel & or1921);
  assign y1922 = (add_sel & s1922) | (sub_sel & sub1922) | (and_sel & and1922) | (or_sel & or1922);
  assign y1923 = (add_sel & s1923) | (sub_sel & sub1923) | (and_sel & and1923) | (or_sel & or1923);
  assign y1924 = (add_sel & s1924) | (sub_sel & sub1924) | (and_sel & and1924) | (or_sel & or1924);
  assign y1925 = (add_sel & s1925) | (sub_sel & sub1925) | (and_sel & and1925) | (or_sel & or1925);
  assign y1926 = (add_sel & s1926) | (sub_sel & sub1926) | (and_sel & and1926) | (or_sel & or1926);
  assign y1927 = (add_sel & s1927) | (sub_sel & sub1927) | (and_sel & and1927) | (or_sel & or1927);
  assign y1928 = (add_sel & s1928) | (sub_sel & sub1928) | (and_sel & and1928) | (or_sel & or1928);
  assign y1929 = (add_sel & s1929) | (sub_sel & sub1929) | (and_sel & and1929) | (or_sel & or1929);
  assign y1930 = (add_sel & s1930) | (sub_sel & sub1930) | (and_sel & and1930) | (or_sel & or1930);
  assign y1931 = (add_sel & s1931) | (sub_sel & sub1931) | (and_sel & and1931) | (or_sel & or1931);
  assign y1932 = (add_sel & s1932) | (sub_sel & sub1932) | (and_sel & and1932) | (or_sel & or1932);
  assign y1933 = (add_sel & s1933) | (sub_sel & sub1933) | (and_sel & and1933) | (or_sel & or1933);
  assign y1934 = (add_sel & s1934) | (sub_sel & sub1934) | (and_sel & and1934) | (or_sel & or1934);
  assign y1935 = (add_sel & s1935) | (sub_sel & sub1935) | (and_sel & and1935) | (or_sel & or1935);
  assign y1936 = (add_sel & s1936) | (sub_sel & sub1936) | (and_sel & and1936) | (or_sel & or1936);
  assign y1937 = (add_sel & s1937) | (sub_sel & sub1937) | (and_sel & and1937) | (or_sel & or1937);
  assign y1938 = (add_sel & s1938) | (sub_sel & sub1938) | (and_sel & and1938) | (or_sel & or1938);
  assign y1939 = (add_sel & s1939) | (sub_sel & sub1939) | (and_sel & and1939) | (or_sel & or1939);
  assign y1940 = (add_sel & s1940) | (sub_sel & sub1940) | (and_sel & and1940) | (or_sel & or1940);
  assign y1941 = (add_sel & s1941) | (sub_sel & sub1941) | (and_sel & and1941) | (or_sel & or1941);
  assign y1942 = (add_sel & s1942) | (sub_sel & sub1942) | (and_sel & and1942) | (or_sel & or1942);
  assign y1943 = (add_sel & s1943) | (sub_sel & sub1943) | (and_sel & and1943) | (or_sel & or1943);
  assign y1944 = (add_sel & s1944) | (sub_sel & sub1944) | (and_sel & and1944) | (or_sel & or1944);
  assign y1945 = (add_sel & s1945) | (sub_sel & sub1945) | (and_sel & and1945) | (or_sel & or1945);
  assign y1946 = (add_sel & s1946) | (sub_sel & sub1946) | (and_sel & and1946) | (or_sel & or1946);
  assign y1947 = (add_sel & s1947) | (sub_sel & sub1947) | (and_sel & and1947) | (or_sel & or1947);
  assign y1948 = (add_sel & s1948) | (sub_sel & sub1948) | (and_sel & and1948) | (or_sel & or1948);
  assign y1949 = (add_sel & s1949) | (sub_sel & sub1949) | (and_sel & and1949) | (or_sel & or1949);
  assign y1950 = (add_sel & s1950) | (sub_sel & sub1950) | (and_sel & and1950) | (or_sel & or1950);
  assign y1951 = (add_sel & s1951) | (sub_sel & sub1951) | (and_sel & and1951) | (or_sel & or1951);
  assign y1952 = (add_sel & s1952) | (sub_sel & sub1952) | (and_sel & and1952) | (or_sel & or1952);
  assign y1953 = (add_sel & s1953) | (sub_sel & sub1953) | (and_sel & and1953) | (or_sel & or1953);
  assign y1954 = (add_sel & s1954) | (sub_sel & sub1954) | (and_sel & and1954) | (or_sel & or1954);
  assign y1955 = (add_sel & s1955) | (sub_sel & sub1955) | (and_sel & and1955) | (or_sel & or1955);
  assign y1956 = (add_sel & s1956) | (sub_sel & sub1956) | (and_sel & and1956) | (or_sel & or1956);
  assign y1957 = (add_sel & s1957) | (sub_sel & sub1957) | (and_sel & and1957) | (or_sel & or1957);
  assign y1958 = (add_sel & s1958) | (sub_sel & sub1958) | (and_sel & and1958) | (or_sel & or1958);
  assign y1959 = (add_sel & s1959) | (sub_sel & sub1959) | (and_sel & and1959) | (or_sel & or1959);
  assign y1960 = (add_sel & s1960) | (sub_sel & sub1960) | (and_sel & and1960) | (or_sel & or1960);
  assign y1961 = (add_sel & s1961) | (sub_sel & sub1961) | (and_sel & and1961) | (or_sel & or1961);
  assign y1962 = (add_sel & s1962) | (sub_sel & sub1962) | (and_sel & and1962) | (or_sel & or1962);
  assign y1963 = (add_sel & s1963) | (sub_sel & sub1963) | (and_sel & and1963) | (or_sel & or1963);
  assign y1964 = (add_sel & s1964) | (sub_sel & sub1964) | (and_sel & and1964) | (or_sel & or1964);
  assign y1965 = (add_sel & s1965) | (sub_sel & sub1965) | (and_sel & and1965) | (or_sel & or1965);
  assign y1966 = (add_sel & s1966) | (sub_sel & sub1966) | (and_sel & and1966) | (or_sel & or1966);
  assign y1967 = (add_sel & s1967) | (sub_sel & sub1967) | (and_sel & and1967) | (or_sel & or1967);
  assign y1968 = (add_sel & s1968) | (sub_sel & sub1968) | (and_sel & and1968) | (or_sel & or1968);
  assign y1969 = (add_sel & s1969) | (sub_sel & sub1969) | (and_sel & and1969) | (or_sel & or1969);
  assign y1970 = (add_sel & s1970) | (sub_sel & sub1970) | (and_sel & and1970) | (or_sel & or1970);
  assign y1971 = (add_sel & s1971) | (sub_sel & sub1971) | (and_sel & and1971) | (or_sel & or1971);
  assign y1972 = (add_sel & s1972) | (sub_sel & sub1972) | (and_sel & and1972) | (or_sel & or1972);
  assign y1973 = (add_sel & s1973) | (sub_sel & sub1973) | (and_sel & and1973) | (or_sel & or1973);
  assign y1974 = (add_sel & s1974) | (sub_sel & sub1974) | (and_sel & and1974) | (or_sel & or1974);
  assign y1975 = (add_sel & s1975) | (sub_sel & sub1975) | (and_sel & and1975) | (or_sel & or1975);
  assign y1976 = (add_sel & s1976) | (sub_sel & sub1976) | (and_sel & and1976) | (or_sel & or1976);
  assign y1977 = (add_sel & s1977) | (sub_sel & sub1977) | (and_sel & and1977) | (or_sel & or1977);
  assign y1978 = (add_sel & s1978) | (sub_sel & sub1978) | (and_sel & and1978) | (or_sel & or1978);
  assign y1979 = (add_sel & s1979) | (sub_sel & sub1979) | (and_sel & and1979) | (or_sel & or1979);
  assign y1980 = (add_sel & s1980) | (sub_sel & sub1980) | (and_sel & and1980) | (or_sel & or1980);
  assign y1981 = (add_sel & s1981) | (sub_sel & sub1981) | (and_sel & and1981) | (or_sel & or1981);
  assign y1982 = (add_sel & s1982) | (sub_sel & sub1982) | (and_sel & and1982) | (or_sel & or1982);
  assign y1983 = (add_sel & s1983) | (sub_sel & sub1983) | (and_sel & and1983) | (or_sel & or1983);
  assign y1984 = (add_sel & s1984) | (sub_sel & sub1984) | (and_sel & and1984) | (or_sel & or1984);
  assign y1985 = (add_sel & s1985) | (sub_sel & sub1985) | (and_sel & and1985) | (or_sel & or1985);
  assign y1986 = (add_sel & s1986) | (sub_sel & sub1986) | (and_sel & and1986) | (or_sel & or1986);
  assign y1987 = (add_sel & s1987) | (sub_sel & sub1987) | (and_sel & and1987) | (or_sel & or1987);
  assign y1988 = (add_sel & s1988) | (sub_sel & sub1988) | (and_sel & and1988) | (or_sel & or1988);
  assign y1989 = (add_sel & s1989) | (sub_sel & sub1989) | (and_sel & and1989) | (or_sel & or1989);
  assign y1990 = (add_sel & s1990) | (sub_sel & sub1990) | (and_sel & and1990) | (or_sel & or1990);
  assign y1991 = (add_sel & s1991) | (sub_sel & sub1991) | (and_sel & and1991) | (or_sel & or1991);
  assign y1992 = (add_sel & s1992) | (sub_sel & sub1992) | (and_sel & and1992) | (or_sel & or1992);
  assign y1993 = (add_sel & s1993) | (sub_sel & sub1993) | (and_sel & and1993) | (or_sel & or1993);
  assign y1994 = (add_sel & s1994) | (sub_sel & sub1994) | (and_sel & and1994) | (or_sel & or1994);
  assign y1995 = (add_sel & s1995) | (sub_sel & sub1995) | (and_sel & and1995) | (or_sel & or1995);
  assign y1996 = (add_sel & s1996) | (sub_sel & sub1996) | (and_sel & and1996) | (or_sel & or1996);
  assign y1997 = (add_sel & s1997) | (sub_sel & sub1997) | (and_sel & and1997) | (or_sel & or1997);
  assign y1998 = (add_sel & s1998) | (sub_sel & sub1998) | (and_sel & and1998) | (or_sel & or1998);
  assign y1999 = (add_sel & s1999) | (sub_sel & sub1999) | (and_sel & and1999) | (or_sel & or1999);
  assign y2000 = (add_sel & s2000) | (sub_sel & sub2000) | (and_sel & and2000) | (or_sel & or2000);
  assign y2001 = (add_sel & s2001) | (sub_sel & sub2001) | (and_sel & and2001) | (or_sel & or2001);
  assign y2002 = (add_sel & s2002) | (sub_sel & sub2002) | (and_sel & and2002) | (or_sel & or2002);
  assign y2003 = (add_sel & s2003) | (sub_sel & sub2003) | (and_sel & and2003) | (or_sel & or2003);
  assign y2004 = (add_sel & s2004) | (sub_sel & sub2004) | (and_sel & and2004) | (or_sel & or2004);
  assign y2005 = (add_sel & s2005) | (sub_sel & sub2005) | (and_sel & and2005) | (or_sel & or2005);
  assign y2006 = (add_sel & s2006) | (sub_sel & sub2006) | (and_sel & and2006) | (or_sel & or2006);
  assign y2007 = (add_sel & s2007) | (sub_sel & sub2007) | (and_sel & and2007) | (or_sel & or2007);
  assign y2008 = (add_sel & s2008) | (sub_sel & sub2008) | (and_sel & and2008) | (or_sel & or2008);
  assign y2009 = (add_sel & s2009) | (sub_sel & sub2009) | (and_sel & and2009) | (or_sel & or2009);
  assign y2010 = (add_sel & s2010) | (sub_sel & sub2010) | (and_sel & and2010) | (or_sel & or2010);
  assign y2011 = (add_sel & s2011) | (sub_sel & sub2011) | (and_sel & and2011) | (or_sel & or2011);
  assign y2012 = (add_sel & s2012) | (sub_sel & sub2012) | (and_sel & and2012) | (or_sel & or2012);
  assign y2013 = (add_sel & s2013) | (sub_sel & sub2013) | (and_sel & and2013) | (or_sel & or2013);
  assign y2014 = (add_sel & s2014) | (sub_sel & sub2014) | (and_sel & and2014) | (or_sel & or2014);
  assign y2015 = (add_sel & s2015) | (sub_sel & sub2015) | (and_sel & and2015) | (or_sel & or2015);
  assign y2016 = (add_sel & s2016) | (sub_sel & sub2016) | (and_sel & and2016) | (or_sel & or2016);
  assign y2017 = (add_sel & s2017) | (sub_sel & sub2017) | (and_sel & and2017) | (or_sel & or2017);
  assign y2018 = (add_sel & s2018) | (sub_sel & sub2018) | (and_sel & and2018) | (or_sel & or2018);
  assign y2019 = (add_sel & s2019) | (sub_sel & sub2019) | (and_sel & and2019) | (or_sel & or2019);
  assign y2020 = (add_sel & s2020) | (sub_sel & sub2020) | (and_sel & and2020) | (or_sel & or2020);
  assign y2021 = (add_sel & s2021) | (sub_sel & sub2021) | (and_sel & and2021) | (or_sel & or2021);
  assign y2022 = (add_sel & s2022) | (sub_sel & sub2022) | (and_sel & and2022) | (or_sel & or2022);
  assign y2023 = (add_sel & s2023) | (sub_sel & sub2023) | (and_sel & and2023) | (or_sel & or2023);
  assign y2024 = (add_sel & s2024) | (sub_sel & sub2024) | (and_sel & and2024) | (or_sel & or2024);
  assign y2025 = (add_sel & s2025) | (sub_sel & sub2025) | (and_sel & and2025) | (or_sel & or2025);
  assign y2026 = (add_sel & s2026) | (sub_sel & sub2026) | (and_sel & and2026) | (or_sel & or2026);
  assign y2027 = (add_sel & s2027) | (sub_sel & sub2027) | (and_sel & and2027) | (or_sel & or2027);
  assign y2028 = (add_sel & s2028) | (sub_sel & sub2028) | (and_sel & and2028) | (or_sel & or2028);
  assign y2029 = (add_sel & s2029) | (sub_sel & sub2029) | (and_sel & and2029) | (or_sel & or2029);
  assign y2030 = (add_sel & s2030) | (sub_sel & sub2030) | (and_sel & and2030) | (or_sel & or2030);
  assign y2031 = (add_sel & s2031) | (sub_sel & sub2031) | (and_sel & and2031) | (or_sel & or2031);
  assign y2032 = (add_sel & s2032) | (sub_sel & sub2032) | (and_sel & and2032) | (or_sel & or2032);
  assign y2033 = (add_sel & s2033) | (sub_sel & sub2033) | (and_sel & and2033) | (or_sel & or2033);
  assign y2034 = (add_sel & s2034) | (sub_sel & sub2034) | (and_sel & and2034) | (or_sel & or2034);
  assign y2035 = (add_sel & s2035) | (sub_sel & sub2035) | (and_sel & and2035) | (or_sel & or2035);
  assign y2036 = (add_sel & s2036) | (sub_sel & sub2036) | (and_sel & and2036) | (or_sel & or2036);
  assign y2037 = (add_sel & s2037) | (sub_sel & sub2037) | (and_sel & and2037) | (or_sel & or2037);
  assign y2038 = (add_sel & s2038) | (sub_sel & sub2038) | (and_sel & and2038) | (or_sel & or2038);
  assign y2039 = (add_sel & s2039) | (sub_sel & sub2039) | (and_sel & and2039) | (or_sel & or2039);
  assign y2040 = (add_sel & s2040) | (sub_sel & sub2040) | (and_sel & and2040) | (or_sel & or2040);
  assign y2041 = (add_sel & s2041) | (sub_sel & sub2041) | (and_sel & and2041) | (or_sel & or2041);
  assign y2042 = (add_sel & s2042) | (sub_sel & sub2042) | (and_sel & and2042) | (or_sel & or2042);
  assign y2043 = (add_sel & s2043) | (sub_sel & sub2043) | (and_sel & and2043) | (or_sel & or2043);
  assign y2044 = (add_sel & s2044) | (sub_sel & sub2044) | (and_sel & and2044) | (or_sel & or2044);
  assign y2045 = (add_sel & s2045) | (sub_sel & sub2045) | (and_sel & and2045) | (or_sel & or2045);
  assign y2046 = (add_sel & s2046) | (sub_sel & sub2046) | (and_sel & and2046) | (or_sel & or2046);
  assign y2047 = (add_sel & s2047) | (sub_sel & sub2047) | (and_sel & and2047) | (or_sel & or2047);
endmodule