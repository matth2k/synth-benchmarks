// IWLS benchmark module "C1355.iscas" printed on Wed May 29 16:27:40 2002
module C1355 (\1GAT(0) , \8GAT(1) , \15GAT(2) , \22GAT(3) , \29GAT(4) , \36GAT(5) , \43GAT(6) , \50GAT(7) , \57GAT(8) , \64GAT(9) , \71GAT(10) , \78GAT(11) , \85GAT(12) , \92GAT(13) , \99GAT(14) , \106GAT(15) , \113GAT(16) , \120GAT(17) , \127GAT(18) , \134GAT(19) , \141GAT(20) , \148GAT(21) , \155GAT(22) , \162GAT(23) , \169GAT(24) , \176GAT(25) , \183GAT(26) , \190GAT(27) , \197GAT(28) , \204GAT(29) , \211GAT(30) , \218GAT(31) , \225GAT(32) , \226GAT(33) , \227GAT(34) , \228GAT(35) , \229GAT(36) , \230GAT(37) , \231GAT(38) , \232GAT(39) , \233GAT(40) , \1324GAT(583) , \1325GAT(579) , \1326GAT(575) , \1327GAT(571) , \1328GAT(584) , \1329GAT(580) , \1330GAT(576) , \1331GAT(572) , \1332GAT(585) , \1333GAT(581) , \1334GAT(577) , \1335GAT(573) , \1336GAT(586) , \1337GAT(582) , \1338GAT(578) , \1339GAT(574) , \1340GAT(567) , \1341GAT(563) , \1342GAT(559) , \1343GAT(555) , \1344GAT(568) , \1345GAT(564) , \1346GAT(560) , \1347GAT(556) , \1348GAT(569) , \1349GAT(565) , \1350GAT(561) , \1351GAT(557) , \1352GAT(570) , \1353GAT(566) , \1354GAT(562) , \1355GAT(558) );
input
  \106GAT(15) ,
  \197GAT(28) ,
  \190GAT(27) ,
  \43GAT(6) ,
  \29GAT(4) ,
  \8GAT(1) ,
  \162GAT(23) ,
  \64GAT(9) ,
  \169GAT(24) ,
  \155GAT(22) ,
  \92GAT(13) ,
  \183GAT(26) ,
  \15GAT(2) ,
  \99GAT(14) ,
  \232GAT(39) ,
  \230GAT(37) ,
  \231GAT(38) ,
  \176GAT(25) ,
  \233GAT(40) ,
  \113GAT(16) ,
  \127GAT(18) ,
  \50GAT(7) ,
  \211GAT(30) ,
  \120GAT(17) ,
  \134GAT(19) ,
  \218GAT(31) ,
  \141GAT(20) ,
  \36GAT(5) ,
  \229GAT(36) ,
  \148GAT(21) ,
  \228GAT(35) ,
  \227GAT(34) ,
  \225GAT(32) ,
  \226GAT(33) ,
  \57GAT(8) ,
  \71GAT(10) ,
  \204GAT(29) ,
  \78GAT(11) ,
  \22GAT(3) ,
  \85GAT(12) ,
  \1GAT(0) ;
output
  \1333GAT(581) ,
  \1341GAT(563) ,
  \1332GAT(585) ,
  \1340GAT(567) ,
  \1330GAT(576) ,
  \1342GAT(559) ,
  \1326GAT(575) ,
  \1331GAT(572) ,
  \1327GAT(571) ,
  \1337GAT(582) ,
  \1343GAT(555) ,
  \1336GAT(586) ,
  \1345GAT(564) ,
  \1344GAT(568) ,
  \1334GAT(577) ,
  \1325GAT(579) ,
  \1352GAT(570) ,
  \1324GAT(583) ,
  \1351GAT(557) ,
  \1350GAT(561) ,
  \1335GAT(573) ,
  \1347GAT(556) ,
  \1346GAT(560) ,
  \1353GAT(566) ,
  \1349GAT(565) ,
  \1348GAT(569) ,
  \1329GAT(580) ,
  \1338GAT(578) ,
  \1355GAT(558) ,
  \1328GAT(584) ,
  \1354GAT(562) ,
  \1339GAT(574) ;
wire
  \601GAT(193) ,
  \483GAT(164) ,
  \812GAT(306) ,
  \1126GAT(402) ,
  \1308GAT(535) ,
  \480GAT(172) ,
  \423GAT(97) ,
  \1239GAT(484) ,
  \1229GAT(487) ,
  \1045GAT(411) ,
  \1283GAT(461) ,
  \588GAT(220) ,
  \415GAT(101) ,
  \456GAT(157) ,
  \1171GAT(445) ,
  \465GAT(151) ,
  \1260GAT(506) ,
  \589GAT(212) ,
  \1244GAT(514) ,
  \1309GAT(531) ,
  \972GAT(371) ,
  \971GAT(360) ,
  \803GAT(309) ,
  \969GAT(341) ,
  \949GAT(359) ,
  \486GAT(171) ,
  \414GAT(109) ,
  \1180GAT(442) ,
  \982GAT(377) ,
  \612GAT(238) ,
  \383GAT(102) ,
  \1236GAT(518) ,
  \1273GAT(464) ,
  \1263GAT(467) ,
  \622GAT(232) ,
  \754GAT(288) ,
  \504GAT(156) ,
  \637GAT(226) ,
  \764GAT(283) ,
  \534GAT(184) ,
  \968GAT(346) ,
  \991GAT(385) ,
  \1270GAT(501) ,
  \948GAT(364) ,
  \1156GAT(450) ,
  \645GAT(236) ,
  \1256GAT(508) ,
  \1090GAT(399) ,
  \477GAT(166) ,
  \471GAT(146) ,
  \642GAT(237) ,
  \1278GAT(497) ,
  \721GAT(265) ,
  \983GAT(378) ,
  \1316GAT(537) ,
  \1288GAT(492) ,
  \382GAT(104) ,
  \938GAT(372) ,
  \1300GAT(553) ,
  \1307GAT(542) ,
  \1114GAT(401) ,
  \1011GAT(388) ,
  \607GAT(239) ,
  \1141GAT(455) ,
  \1275GAT(460) ,
  \1306GAT(546) ,
  \712GAT(271) ,
  \381GAT(106) ,
  \474GAT(174) ,
  \583GAT(199) ,
  \773GAT(303) ,
  \525GAT(191) ,
  \957GAT(343) ,
  \552GAT(187) ,
  \590GAT(219) ,
  \1287GAT(470) ,
  \1261GAT(471) ,
  \1315GAT(524) ,
  \305GAT(53) ,
  \1246GAT(513) ,
  \970GAT(370) ,
  \742GAT(276) ,
  \1219GAT(429) ,
  \398GAT(141) ,
  \302GAT(56) ,
  \308GAT(50) ,
  \973GAT(365) ,
  \1314GAT(528) ,
  \1251GAT(477) ,
  \632GAT(230) ,
  \332GAT(75) ,
  \996GAT(389) ,
  \598GAT(203) ,
  \399GAT(133) ,
  \819GAT(320) ,
  \1266GAT(503) ,
  \380GAT(108) ,
  \1132GAT(458) ,
  \1036GAT(423) ,
  \1265GAT(463) ,
  \1240GAT(516) ,
  \329GAT(68) ,
  \765GAT(293) ,
  \1096GAT(408) ,
  \873GAT(333) ,
  \599GAT(195) ,
  \574GAT(216) ,
  \1277GAT(473) ,
  \976GAT(376) ,
  \1254GAT(509) ,
  \981GAT(384) ,
  \818GAT(328) ,
  \1317GAT(533) ,
  \782GAT(300) ,
  \966GAT(340) ,
  \691GAT(261) ,
  \1078GAT(418) ,
  \785GAT(299) ,
  \1230GAT(521) ,
  \975GAT(361) ,
  \1087GAT(403) ,
  \961GAT(355) ,
  \459GAT(154) ,
  \591GAT(211) ,
  \441GAT(167) ,
  \1257GAT(482) ,
  \432GAT(173) ,
  \755GAT(292) ,
  \669GAT(245) ,
  \408GAT(121) ,
  \733GAT(279) ,
  \421GAT(83) ,
  \1001GAT(387) ,
  \549GAT(188) ,
  \378GAT(112) ,
  \424GAT(89) ,
  \791GAT(297) ,
  \561GAT(180) ,
  \409GAT(113) ,
  \955GAT(338) ,
  \592GAT(217) ,
  \1144GAT(454) ,
  \980GAT(383) ,
  \1042GAT(415) ,
  \962GAT(350) ,
  \1285GAT(474) ,
  \425GAT(81) ,
  \418GAT(107) ,
  \1303GAT(541) ,
  \965GAT(345) ,
  \768GAT(281) ,
  \379GAT(110) ,
  \829GAT(315) ,
  \314GAT(79) ,
  \575GAT(215) ,
  \1264GAT(504) ,
  \489GAT(163) ,
  \690GAT(263) ,
  \1289GAT(466) ,
  \828GAT(323) ,
  \1304GAT(554) ,
  \767GAT(295) ,
  \1255GAT(486) ,
  \692GAT(259) ,
  \1312GAT(536) ,
  \986GAT(386) ,
  \770GAT(304) ,
  \815GAT(305) ,
  \758GAT(286) ,
  \1267GAT(459) ,
  \317GAT(71) ,
  \1093GAT(395) ,
  \579GAT(207) ,
  \724GAT(267) ,
  \410GAT(111) ,
  \260GAT(42) ,
  \977GAT(366) ,
  \1135GAT(457) ,
  \344GAT(62) ,
  \368GAT(132) ,
  \1274GAT(499) ,
  \1279GAT(469) ,
  \964GAT(356) ,
  \953GAT(342) ,
  \954GAT(352) ,
  \1120GAT(410) ,
  \806GAT(308) ,
  \1243GAT(476) ,
  \700GAT(251) ,
  \1284GAT(494) ,
  \1242GAT(515) ,
  \263GAT(41) ,
  \952GAT(348) ,
  \335GAT(67) ,
  \426GAT(176) ,
  \417GAT(85) ,
  \1232GAT(520) ,
  \1299GAT(540) ,
  \1305GAT(550) ,
  \1311GAT(523) ,
  \341GAT(55) ,
  \326GAT(76) ,
  \602GAT(240) ,
  \413GAT(87) ,
  \984GAT(379) ,
  \1225GAT(427) ,
  \1302GAT(545) ,
  \974GAT(375) ,
  \1084GAT(407) ,
  \323GAT(70) ,
  \1310GAT(527) ,
  \576GAT(213) ,
  \397GAT(119) ,
  \356GAT(59) ,
  \1108GAT(409) ,
  \369GAT(130) ,
  \1233GAT(479) ,
  \1069GAT(413) ,
  \396GAT(127) ,
  \1322GAT(530) ,
  \1198GAT(436) ,
  \353GAT(52) ,
  \567GAT(177) ,
  \693GAT(257) ,
  \1301GAT(549) ,
  \578GAT(208) ,
  \666GAT(248) ,
  \338GAT(63) ,
  \593GAT(209) ,
  \587GAT(214) ,
  \963GAT(339) ,
  \860GAT(334) ,
  \736GAT(278) ,
  \727GAT(266) ,
  \586GAT(222) ,
  \985GAT(380) ,
  \347GAT(54) ,
  \251GAT(45) ,
  \730GAT(280) ,
  \320GAT(78) ,
  \406GAT(137) ,
  \595GAT(198) ,
  \245GAT(47) ,
  \272GAT(74) ,
  \366GAT(136) ,
  \519GAT(145) ,
  \577GAT(210) ,
  \1129GAT(398) ,
  \395GAT(135) ,
  \1313GAT(532) ,
  \761GAT(290) ,
  \359GAT(51) ,
  \654GAT(229) ,
  \394GAT(143) ,
  \695GAT(260) ,
  \248GAT(46) ,
  \1241GAT(480) ,
  \1298GAT(544) ,
  \1216GAT(430) ,
  \564GAT(179) ,
  \678GAT(244) ,
  \555GAT(185) ,
  \278GAT(72) ,
  \834GAT(336) ,
  \776GAT(302) ,
  \1297GAT(548) ,
  \254GAT(44) ,
  \257GAT(43) ,
  \702GAT(256) ,
  \571GAT(223) ,
  \350GAT(60) ,
  \275GAT(73) ,
  \242GAT(48) ,
  \847GAT(335) ,
  \1147GAT(453) ,
  \956GAT(353) ,
  \384GAT(100) ,
  \687GAT(242) ,
  \1258GAT(507) ,
  \1276GAT(498) ,
  \522GAT(192) ,
  \1320GAT(538) ,
  \1286GAT(493) ,
  \1189GAT(439) ,
  \951GAT(337) ,
  \950GAT(347) ,
  \1323GAT(526) ,
  \657GAT(228) ,
  \1231GAT(483) ,
  \899GAT(329) ,
  \694GAT(264) ,
  \405GAT(115) ,
  \1250GAT(511) ,
  \825GAT(317) ,
  \570GAT(224) ,
  \375GAT(118) ,
  \404GAT(123) ,
  \367GAT(134) ,
  \407GAT(129) ,
  \1247GAT(485) ,
  \715GAT(270) ,
  \1237GAT(488) ,
  \1138GAT(456) ,
  \763GAT(296) ,
  \1075GAT(422) ,
  \1290GAT(491) ,
  \284GAT(66) ,
  \444GAT(165) ,
  \510GAT(155) ,
  \597GAT(196) ,
  \1159GAT(449) ,
  \374GAT(120) ,
  \967GAT(351) ,
  \794GAT(312) ,
  \824GAT(325) ,
  \1280GAT(496) ,
  \1099GAT(404) ,
  \703GAT(252) ,
  \1268GAT(502) ,
  \1207GAT(433) ,
  \960GAT(344) ,
  \1054GAT(416) ,
  \1123GAT(406) ,
  \266GAT(80) ,
  \704GAT(254) ,
  \1168GAT(446) ,
  \706GAT(272) ,
  \745GAT(275) ,
  \1321GAT(534) ,
  \376GAT(116) ,
  \958GAT(354) ,
  \697GAT(258) ,
  \287GAT(65) ,
  \940GAT(362) ,
  \675GAT(246) ,
  \573GAT(218) ,
  \281GAT(69) ,
  \365GAT(138) ,
  \660GAT(227) ,
  \468GAT(149) ,
  \1292GAT(551) ,
  \1245GAT(489) ,
  \402GAT(139) ,
  \435GAT(170) ,
  \311GAT(49) ,
  \447GAT(162) ,
  \269GAT(77) ,
  \1259GAT(478) ,
  \705GAT(250) ,
  \718GAT(268) ,
  \572GAT(221) ,
  \1204GAT(434) ,
  \1016GAT(393) ,
  \364GAT(140) ,
  \831GAT(314) ,
  \1269GAT(472) ,
  \979GAT(382) ,
  \492GAT(169) ,
  \1295GAT(539) ,
  \1186GAT(440) ,
  \830GAT(322) ,
  \1177GAT(443) ,
  \1252GAT(510) ,
  \827GAT(316) ,
  \1238GAT(517) ,
  \696GAT(262) ,
  \1066GAT(417) ,
  \701GAT(249) ,
  \684GAT(243) ,
  \942GAT(368) ,
  \584GAT(197) ,
  \1293GAT(547) ,
  \809GAT(307) ,
  \943GAT(357) ,
  \1026GAT(394) ,
  \296GAT(58) ,
  \978GAT(381) ,
  \371GAT(126) ,
  \363GAT(142) ,
  \401GAT(117) ,
  \826GAT(324) ,
  \299GAT(57) ,
  \495GAT(161) ,
  \377GAT(114) ,
  \1294GAT(543) ,
  \762GAT(284) ,
  \1195GAT(437) ,
  \698GAT(255) ,
  \543GAT(178) ,
  \663GAT(225) ,
  \403GAT(131) ,
  \1213GAT(431) ,
  \422GAT(105) ,
  \438GAT(168) ,
  \582GAT(200) ,
  \1192GAT(438) ,
  \797GAT(311) ,
  \941GAT(373) ,
  \513GAT(147) ,
  \821GAT(319) ,
  \1228GAT(522) ,
  \1039GAT(419) ,
  \400GAT(125) ,
  \450GAT(160) ,
  \820GAT(327) ,
  \1282GAT(495) ,
  \531GAT(186) ,
  \1048GAT(424) ,
  \370GAT(128) ,
  \362GAT(144) ,
  \945GAT(363) ,
  \672GAT(247) ,
  \1150GAT(452) ,
  \1031GAT(392) ,
  \411GAT(103) ,
  \600GAT(201) ,
  \779GAT(301) ,
  \832GAT(321) ,
  \290GAT(64) ,
  \1248GAT(512) ,
  \1006GAT(390) ,
  \558GAT(181) ,
  \293GAT(61) ,
  \1102GAT(400) ,
  \1081GAT(414) ,
  \596GAT(204) ,
  \912GAT(330) ,
  \1117GAT(397) ,
  \1235GAT(475) ,
  \1222GAT(428) ,
  \833GAT(313) ,
  \1165GAT(447) ,
  \648GAT(235) ,
  \699GAT(253) ,
  \1105GAT(396) ,
  \585GAT(194) ,
  \800GAT(310) ,
  \681GAT(241) ,
  \709GAT(269) ,
  \748GAT(274) ,
  \1111GAT(405) ,
  \1183GAT(441) ,
  \528GAT(190) ,
  \581GAT(202) ,
  \1210GAT(432) ,
  \947GAT(369) ,
  \1051GAT(420) ,
  \925GAT(332) ,
  \946GAT(358) ,
  \1057GAT(412) ,
  \507GAT(148) ,
  \453GAT(159) ,
  \392GAT(84) ,
  \1291GAT(462) ,
  \760GAT(285) ,
  \651GAT(233) ,
  \386GAT(96) ,
  \393GAT(82) ,
  \385GAT(98) ,
  \1174GAT(444) ,
  \757GAT(289) ,
  \429GAT(175) ,
  \1060GAT(425) ,
  \412GAT(95) ,
  \1021GAT(391) ,
  \739GAT(277) ,
  \1296GAT(552) ,
  \594GAT(206) ,
  \373GAT(122) ,
  \823GAT(318) ,
  \388GAT(92) ,
  \580GAT(205) ,
  \1281GAT(465) ,
  \537GAT(183) ,
  \1271GAT(468) ,
  \462GAT(152) ,
  \627GAT(231) ,
  \822GAT(326) ,
  \944GAT(374) ,
  \1319GAT(525) ,
  \419GAT(99) ,
  \391GAT(86) ,
  \387GAT(94) ,
  \751GAT(273) ,
  \390GAT(88) ,
  \1318GAT(529) ,
  \389GAT(90) ,
  \540GAT(182) ,
  \788GAT(298) ,
  \1072GAT(426) ,
  \1063GAT(421) ,
  \516GAT(153) ,
  \1262GAT(505) ,
  \1234GAT(519) ,
  \1249GAT(481) ,
  \416GAT(93) ,
  \939GAT(367) ,
  \1201GAT(435) ,
  \1153GAT(451) ,
  \372GAT(124) ,
  \546GAT(189) ,
  \769GAT(294) ,
  \756GAT(287) ,
  \501GAT(150) ,
  \1162GAT(448) ,
  \1253GAT(490) ,
  \498GAT(158) ,
  \766GAT(282) ,
  \617GAT(234) ,
  \886GAT(331) ,
  \959GAT(349) ,
  \1272GAT(500) ,
  \420GAT(91) ,
  \759GAT(291) ;
assign
  \601GAT(193)  = ~\567GAT(177)  | ~\519GAT(145) ,
  \483GAT(164)  = ~\401GAT(117)  | ~\400GAT(125) ,
  \812GAT(306)  = ~\788GAT(298)  | ~\660GAT(227) ,
  \1126GAT(402)  = \1031GAT(392)  & \912GAT(330) ,
  \1308GAT(535)  = ~\1261GAT(471)  | ~\1260GAT(506) ,
  \480GAT(172)  = ~\399GAT(133)  | ~\398GAT(141) ,
  \423GAT(97)  = ~\356GAT(59)  | ~\162GAT(23) ,
  \1239GAT(484)  = ~\1147GAT(453)  | ~\1051GAT(420) ,
  \1229GAT(487)  = ~\1132GAT(458)  | ~\1036GAT(423) ,
  \1045GAT(411)  = \996GAT(389)  & \873GAT(333) ,
  \1283GAT(461)  = ~\1213GAT(431)  | ~\1117GAT(397) ,
  \588GAT(220)  = ~\549GAT(188)  | ~\480GAT(172) ,
  \415GAT(101)  = ~\344GAT(62)  | ~\148GAT(21) ,
  \456GAT(157)  = ~\383GAT(102)  | ~\382GAT(104) ,
  \1171GAT(445)  = ~\1075GAT(422)  | ~\92GAT(13) ,
  \465GAT(151)  = ~\389GAT(90)  | ~\388GAT(92) ,
  \1260GAT(506)  = ~\1180GAT(442)  | ~\113GAT(16) ,
  \589GAT(212)  = ~\549GAT(188)  | ~\483GAT(164) ,
  \1244GAT(514)  = ~\1156GAT(450)  | ~\57GAT(8) ,
  \1309GAT(531)  = ~\1263GAT(467)  | ~\1262GAT(505) ,
  \972GAT(371)  = ~\847GAT(335) ,
  \971GAT(360)  = ~\873GAT(333) ,
  \803GAT(309)  = ~\779GAT(301)  | ~\651GAT(233) ,
  \969GAT(341)  = ~\899GAT(329) ,
  \949GAT(359)  = ~\873GAT(333) ,
  \486GAT(171)  = ~\403GAT(131)  | ~\402GAT(139) ,
  \414GAT(109)  = ~\344GAT(62)  | ~\120GAT(17) ,
  \1180GAT(442)  = ~\1084GAT(407)  | ~\113GAT(16) ,
  \982GAT(377)  = \899GAT(329)  & (\960GAT(344)  & (\959GAT(349)  & \958GAT(354) )),
  \612GAT(238)  = ~\575GAT(215)  | ~\574GAT(216) ,
  \383GAT(102)  = ~\296GAT(58)  | ~\148GAT(21) ,
  \1236GAT(518)  = ~\1144GAT(454)  | ~\29GAT(4) ,
  \1273GAT(464)  = ~\1198GAT(436)  | ~\1102GAT(400) ,
  \1263GAT(467)  = ~\1183GAT(441)  | ~\1087GAT(403) ,
  \622GAT(232)  = ~\579GAT(207)  | ~\578GAT(208) ,
  \754GAT(288)  = ~\730GAT(280)  | ~\242GAT(48) ,
  \504GAT(156)  = ~\415GAT(101)  | ~\414GAT(109) ,
  \637GAT(226)  = ~\585GAT(194)  | ~\584GAT(197) ,
  \764GAT(283)  = ~\745GAT(275)  | ~\257GAT(43) ,
  \534GAT(184)  = ~\453GAT(159)  | ~\450GAT(160) ,
  \968GAT(346)  = ~\912GAT(330) ,
  \991GAT(385)  = \985GAT(380)  | (\984GAT(379)  | (\983GAT(378)  | \982GAT(377) )),
  \1270GAT(501)  = ~\1195GAT(437)  | ~\148GAT(21) ,
  \948GAT(364)  = ~\860GAT(334) ,
  \1156GAT(450)  = ~\1060GAT(425)  | ~\57GAT(8) ,
  \645GAT(236)  = ~\589GAT(212)  | ~\588GAT(220) ,
  \1256GAT(508)  = ~\1174GAT(444)  | ~\99GAT(14) ,
  \1090GAT(399)  = \1016GAT(393)  & \912GAT(330) ,
  \477GAT(166)  = ~\397GAT(119)  | ~\396GAT(127) ,
  \471GAT(146)  = ~\393GAT(82)  | ~\392GAT(84) ,
  \642GAT(237)  = ~\587GAT(214)  | ~\586GAT(222) ,
  \1278GAT(497)  = ~\1207GAT(433)  | ~\176GAT(25) ,
  \721GAT(265)  = ~\701GAT(249)  | ~\700GAT(251) ,
  \983GAT(378)  = \963GAT(339)  & (\912GAT(330)  & (\962GAT(350)  & \961GAT(355) )),
  \1316GAT(537)  = ~\1277GAT(473)  | ~\1276GAT(498) ,
  \1288GAT(492)  = ~\1222GAT(428)  | ~\211GAT(30) ,
  \382GAT(104)  = ~\296GAT(58)  | ~\141GAT(20) ,
  \938GAT(372)  = ~\834GAT(336) ,
  \1300GAT(553)  = ~\1245GAT(489)  | ~\1244GAT(514) ,
  \1307GAT(542)  = ~\1259GAT(478)  | ~\1258GAT(507) ,
  \1114GAT(401)  = \1026GAT(394)  & \912GAT(330) ,
  \1011GAT(388)  = \986GAT(386)  & (\899GAT(329)  & (\957GAT(343)  & (\886GAT(331)  & \956GAT(353) ))),
  \607GAT(239)  = ~\573GAT(218)  | ~\572GAT(221) ,
  \1141GAT(455)  = ~\1045GAT(411)  | ~\22GAT(3) ,
  \1275GAT(460)  = ~\1201GAT(435)  | ~\1105GAT(396) ,
  \1306GAT(546)  = ~\1257GAT(482)  | ~\1256GAT(508) ,
  \712GAT(271)  = ~\695GAT(260)  | ~\694GAT(264) ,
  \381GAT(106)  = ~\293GAT(61)  | ~\134GAT(19) ,
  \474GAT(174)  = ~\395GAT(135)  | ~\394GAT(143) ,
  \583GAT(199)  = ~\540GAT(182)  | ~\465GAT(151) ,
  \773GAT(303)  = ~\757GAT(289)  | ~\756GAT(287) ,
  \525GAT(191)  = ~\435GAT(170)  | ~\432GAT(173) ,
  \957GAT(343)  = ~\912GAT(330) ,
  \552GAT(187)  = ~\489GAT(163)  | ~\486GAT(171) ,
  \590GAT(219)  = ~\552GAT(187)  | ~\486GAT(171) ,
  \1287GAT(470)  = ~\1219GAT(429)  | ~\1123GAT(406) ,
  \1261GAT(471)  = ~\1180GAT(442)  | ~\1084GAT(407) ,
  \1315GAT(524)  = ~\1275GAT(460)  | ~\1274GAT(499) ,
  \305GAT(53)  = ~\190GAT(27)  | ~\183GAT(26) ,
  \1246GAT(513)  = ~\1159GAT(449)  | ~\64GAT(9) ,
  \970GAT(370)  = ~\847GAT(335) ,
  \742GAT(276)  = ~\706GAT(272)  | ~\254GAT(44) ,
  \1219GAT(429)  = ~\1123GAT(406)  | ~\204GAT(29) ,
  \398GAT(141)  = ~\320GAT(78)  | ~\8GAT(1) ,
  \302GAT(56)  = ~\176GAT(25)  | ~\169GAT(24) ,
  \308GAT(50)  = ~\204GAT(29)  | ~\197GAT(28) ,
  \973GAT(365)  = ~\860GAT(334) ,
  \1314GAT(528)  = ~\1273GAT(464)  | ~\1272GAT(500) ,
  \1251GAT(477)  = ~\1165GAT(447)  | ~\1069GAT(413) ,
  \632GAT(230)  = ~\583GAT(199)  | ~\582GAT(200) ,
  \332GAT(75)  = ~\50GAT(7)  | ~\22GAT(3) ,
  \996GAT(389)  = \986GAT(386)  & (\951GAT(337)  & (\912GAT(330)  & (\950GAT(347)  & \925GAT(332) ))),
  \598GAT(203)  = ~\564GAT(179)  | ~\510GAT(155) ,
  \399GAT(133)  = ~\320GAT(78)  | ~\36GAT(5) ,
  \819GAT(320)  = ~\794GAT(312)  | ~\770GAT(304) ,
  \1266GAT(503)  = ~\1189GAT(439)  | ~\134GAT(19) ,
  \380GAT(108)  = ~\293GAT(61)  | ~\127GAT(18) ,
  \1132GAT(458)  = ~\1036GAT(423)  | ~\1GAT(0) ,
  \1036GAT(423)  = \996GAT(389)  & \834GAT(336) ,
  \1265GAT(463)  = ~\1186GAT(440)  | ~\1090GAT(399) ,
  \1240GAT(516)  = ~\1150GAT(452)  | ~\43GAT(6) ,
  \329GAT(68)  = ~\99GAT(14)  | ~\71GAT(10) ,
  \765GAT(293)  = ~\745GAT(275)  | ~\709GAT(269) ,
  \1096GAT(408)  = \1021GAT(391)  & \925GAT(332) ,
  \873GAT(333)  = ~\825GAT(317)  | ~\824GAT(325) ,
  \599GAT(195)  = ~\564GAT(179)  | ~\513GAT(147) ,
  \574GAT(216)  = ~\528GAT(190)  | ~\438GAT(168) ,
  \1277GAT(473)  = ~\1204GAT(434)  | ~\1108GAT(409) ,
  \976GAT(376)  = ~\834GAT(336) ,
  \1254GAT(509)  = ~\1171GAT(445)  | ~\92GAT(13) ,
  \981GAT(384)  = \949GAT(359)  & (\948GAT(364)  & (\947GAT(369)  & \834GAT(336) )),
  \818GAT(328)  = ~\794GAT(312)  | ~\642GAT(237) ,
  \1317GAT(533)  = ~\1279GAT(469)  | ~\1278GAT(497) ,
  \1333GAT(581)  = \1301GAT(549) ,
  \782GAT(300)  = ~\763GAT(296)  | ~\762GAT(284) ,
  \966GAT(340)  = ~\899GAT(329) ,
  \691GAT(261)  = ~\666GAT(248)  | ~\607GAT(239) ,
  \1078GAT(418)  = \1011GAT(388)  & \860GAT(334) ,
  \785GAT(299)  = ~\765GAT(293)  | ~\764GAT(283) ,
  \1230GAT(521)  = ~\1135GAT(457)  | ~\8GAT(1) ,
  \975GAT(361)  = ~\873GAT(333) ,
  \1087GAT(403)  = \1016GAT(393)  & \886GAT(331) ,
  \961GAT(355)  = ~\925GAT(332) ,
  \459GAT(154)  = ~\385GAT(98)  | ~\384GAT(100) ,
  \591GAT(211)  = ~\552GAT(187)  | ~\489GAT(163) ,
  \441GAT(167)  = ~\373GAT(122)  | ~\372GAT(124) ,
  \1257GAT(482)  = ~\1174GAT(444)  | ~\1078GAT(418) ,
  \432GAT(173)  = ~\367GAT(134)  | ~\366GAT(136) ,
  \755GAT(292)  = ~\730GAT(280)  | ~\718GAT(268) ,
  \669GAT(245)  = ~\617GAT(234)  | ~\612GAT(238) ,
  \408GAT(121)  = ~\335GAT(67)  | ~\78GAT(11) ,
  \733GAT(279)  = ~\721GAT(265)  | ~\245GAT(47) ,
  \421GAT(83)  = ~\353GAT(52)  | ~\211GAT(30) ,
  \1001GAT(387)  = \986GAT(386)  & (\899GAT(329)  & (\953GAT(342)  & (\952GAT(348)  & \925GAT(332) ))),
  \549GAT(188)  = ~\483GAT(164)  | ~\480GAT(172) ,
  \378GAT(112)  = ~\290GAT(64)  | ~\113GAT(16) ,
  \424GAT(89)  = ~\359GAT(51)  | ~\190GAT(27) ,
  \791GAT(297)  = ~\769GAT(294)  | ~\768GAT(281) ,
  \561GAT(180)  = ~\507GAT(148)  | ~\504GAT(156) ,
  \409GAT(113)  = ~\335GAT(67)  | ~\106GAT(15) ,
  \955GAT(338)  = ~\899GAT(329) ,
  \592GAT(217)  = ~\555GAT(185)  | ~\492GAT(169) ,
  \1144GAT(454)  = ~\1048GAT(424)  | ~\29GAT(4) ,
  \980GAT(383)  = \946GAT(358)  & (\945GAT(363)  & (\847GAT(335)  & \944GAT(374) )),
  \1042GAT(415)  = \996GAT(389)  & \860GAT(334) ,
  \962GAT(350)  = ~\886GAT(331) ,
  \1341GAT(563)  = \1309GAT(531) ,
  \1285GAT(474)  = ~\1216GAT(430)  | ~\1120GAT(410) ,
  \425GAT(81)  = ~\359GAT(51)  | ~\218GAT(31) ,
  \418GAT(107)  = ~\350GAT(60)  | ~\127GAT(18) ,
  \1303GAT(541)  = ~\1251GAT(477)  | ~\1250GAT(511) ,
  \1332GAT(585)  = \1300GAT(553) ,
  \965GAT(345)  = ~\912GAT(330) ,
  \768GAT(281)  = ~\751GAT(273)  | ~\263GAT(41) ,
  \379GAT(110)  = ~\290GAT(64)  | ~\120GAT(17) ,
  \1340GAT(567)  = \1308GAT(535) ,
  \829GAT(315)  = ~\809GAT(307)  | ~\785GAT(299) ,
  \314GAT(79)  = ~\29GAT(4)  | ~\1GAT(0) ,
  \575GAT(215)  = ~\528GAT(190)  | ~\441GAT(167) ,
  \1264GAT(504)  = ~\1186GAT(440)  | ~\127GAT(18) ,
  \489GAT(163)  = ~\405GAT(115)  | ~\404GAT(123) ,
  \690GAT(263)  = ~\666GAT(248)  | ~\602GAT(240) ,
  \1289GAT(466)  = ~\1222GAT(428)  | ~\1126GAT(402) ,
  \828GAT(323)  = ~\809GAT(307)  | ~\657GAT(228) ,
  \1304GAT(554)  = ~\1253GAT(490)  | ~\1252GAT(510) ,
  \767GAT(295)  = ~\748GAT(274)  | ~\712GAT(271) ,
  \1255GAT(486)  = ~\1171GAT(445)  | ~\1075GAT(422) ,
  \692GAT(259)  = ~\669GAT(245)  | ~\612GAT(238) ,
  \1312GAT(536)  = ~\1269GAT(472)  | ~\1268GAT(502) ,
  \986GAT(386)  = \981GAT(384)  | (\980GAT(383)  | (\979GAT(382)  | \978GAT(381) )),
  \770GAT(304)  = ~\755GAT(292)  | ~\754GAT(288) ,
  \815GAT(305)  = ~\791GAT(297)  | ~\663GAT(225) ,
  \758GAT(286)  = ~\736GAT(278)  | ~\248GAT(46) ,
  \1330GAT(576)  = \1298GAT(544) ,
  \1267GAT(459)  = ~\1189GAT(439)  | ~\1093GAT(395) ,
  \317GAT(71)  = ~\85GAT(12)  | ~\57GAT(8) ,
  \1093GAT(395)  = \1016GAT(393)  & \899GAT(329) ,
  \579GAT(207)  = ~\534GAT(184)  | ~\453GAT(159) ,
  \724GAT(267)  = ~\703GAT(252)  | ~\702GAT(256) ,
  \410GAT(111)  = ~\338GAT(63)  | ~\113GAT(16) ,
  \260GAT(42)  = \233GAT(40)  & \231GAT(38) ,
  \977GAT(366)  = ~\860GAT(334) ,
  \1135GAT(457)  = ~\1039GAT(419)  | ~\8GAT(1) ,
  \344GAT(62)  = ~\148GAT(21)  | ~\120GAT(17) ,
  \368GAT(132)  = ~\275GAT(73)  | ~\43GAT(6) ,
  \1274GAT(499)  = ~\1201GAT(435)  | ~\162GAT(23) ,
  \1279GAT(469)  = ~\1207GAT(433)  | ~\1111GAT(405) ,
  \964GAT(356)  = ~\925GAT(332) ,
  \953GAT(342)  = ~\912GAT(330) ,
  \954GAT(352)  = ~\925GAT(332) ,
  \1120GAT(410)  = \1031GAT(392)  & \925GAT(332) ,
  \806GAT(308)  = ~\782GAT(300)  | ~\654GAT(229) ,
  \1243GAT(476)  = ~\1153GAT(451)  | ~\1057GAT(412) ,
  \700GAT(251)  = ~\681GAT(241)  | ~\632GAT(230) ,
  \1284GAT(494)  = ~\1216GAT(430)  | ~\197GAT(28) ,
  \1242GAT(515)  = ~\1153GAT(451)  | ~\50GAT(7) ,
  \263GAT(41)  = \233GAT(40)  & \232GAT(39) ,
  \952GAT(348)  = ~\886GAT(331) ,
  \335GAT(67)  = ~\106GAT(15)  | ~\78GAT(11) ,
  \1342GAT(559)  = \1310GAT(527) ,
  \426GAT(176)  = ~\363GAT(142)  | ~\362GAT(144) ,
  \417GAT(85)  = ~\347GAT(54)  | ~\204GAT(29) ,
  \1232GAT(520)  = ~\1138GAT(456)  | ~\15GAT(2) ,
  \1299GAT(540)  = ~\1243GAT(476)  | ~\1242GAT(515) ,
  \1305GAT(550)  = ~\1255GAT(486)  | ~\1254GAT(509) ,
  \1311GAT(523)  = ~\1267GAT(459)  | ~\1266GAT(503) ,
  \341GAT(55)  = ~\197GAT(28)  | ~\169GAT(24) ,
  \326GAT(76)  = ~\43GAT(6)  | ~\15GAT(2) ,
  \602GAT(240)  = ~\571GAT(223)  | ~\570GAT(224) ,
  \413GAT(87)  = ~\341GAT(55)  | ~\197GAT(28) ,
  \984GAT(379)  = \966GAT(340)  & (\965GAT(345)  & (\886GAT(331)  & \964GAT(356) )),
  \1225GAT(427)  = ~\1129GAT(398)  | ~\218GAT(31) ,
  \1302GAT(545)  = ~\1249GAT(481)  | ~\1248GAT(512) ,
  \974GAT(375)  = ~\834GAT(336) ,
  \1084GAT(407)  = \1016GAT(393)  & \925GAT(332) ,
  \323GAT(70)  = ~\92GAT(13)  | ~\64GAT(9) ,
  \1310GAT(527)  = ~\1265GAT(463)  | ~\1264GAT(504) ,
  \576GAT(213)  = ~\531GAT(186)  | ~\444GAT(165) ,
  \397GAT(119)  = ~\317GAT(71)  | ~\85GAT(12) ,
  \356GAT(59)  = ~\162GAT(23)  | ~\134GAT(19) ,
  \1108GAT(409)  = \1026GAT(394)  & \925GAT(332) ,
  \369GAT(130)  = ~\275GAT(73)  | ~\50GAT(7) ,
  \1233GAT(479)  = ~\1138GAT(456)  | ~\1042GAT(415) ,
  \1069GAT(413)  = \1006GAT(390)  & \873GAT(333) ,
  \396GAT(127)  = ~\317GAT(71)  | ~\57GAT(8) ,
  \1322GAT(530)  = ~\1289GAT(466)  | ~\1288GAT(492) ,
  \1198GAT(436)  = ~\1102GAT(400)  | ~\155GAT(22) ,
  \353GAT(52)  = ~\211GAT(30)  | ~\183GAT(26) ,
  \567GAT(177)  = ~\519GAT(145)  | ~\516GAT(153) ,
  \693GAT(257)  = ~\669GAT(245)  | ~\617GAT(234) ,
  \1301GAT(549)  = ~\1247GAT(485)  | ~\1246GAT(513) ,
  \578GAT(208)  = ~\534GAT(184)  | ~\450GAT(160) ,
  \666GAT(248)  = ~\607GAT(239)  | ~\602GAT(240) ,
  \338GAT(63)  = ~\141GAT(20)  | ~\113GAT(16) ,
  \593GAT(209)  = ~\555GAT(185)  | ~\495GAT(161) ,
  \587GAT(214)  = ~\546GAT(189)  | ~\477GAT(166) ,
  \963GAT(339)  = ~\899GAT(329) ,
  \860GAT(334)  = ~\823GAT(318)  | ~\822GAT(326) ,
  \1326GAT(575)  = \1294GAT(543) ,
  \736GAT(278)  = ~\724GAT(267)  | ~\248GAT(46) ,
  \727GAT(266)  = ~\705GAT(250)  | ~\704GAT(254) ,
  \586GAT(222)  = ~\546GAT(189)  | ~\474GAT(174) ,
  \985GAT(380)  = \969GAT(341)  & (\968GAT(346)  & (\967GAT(351)  & \925GAT(332) )),
  \347GAT(54)  = ~\204GAT(29)  | ~\176GAT(25) ,
  \251GAT(45)  = \233GAT(40)  & \228GAT(35) ,
  \730GAT(280)  = ~\718GAT(268)  | ~\242GAT(48) ,
  \320GAT(78)  = ~\36GAT(5)  | ~\8GAT(1) ,
  \406GAT(137)  = ~\332GAT(75)  | ~\22GAT(3) ,
  \595GAT(198)  = ~\558GAT(181)  | ~\501GAT(150) ,
  \245GAT(47)  = \233GAT(40)  & \226GAT(33) ,
  \272GAT(74)  = ~\36GAT(5)  | ~\29GAT(4) ,
  \366GAT(136)  = ~\272GAT(74)  | ~\29GAT(4) ,
  \519GAT(145)  = ~\425GAT(81)  | ~\424GAT(89) ,
  \577GAT(210)  = ~\531GAT(186)  | ~\447GAT(162) ,
  \1129GAT(398)  = \1031GAT(392)  & \899GAT(329) ,
  \395GAT(135)  = ~\314GAT(79)  | ~\29GAT(4) ,
  \1313GAT(532)  = ~\1271GAT(468)  | ~\1270GAT(501) ,
  \761GAT(290)  = ~\739GAT(277)  | ~\727GAT(266) ,
  \359GAT(51)  = ~\218GAT(31)  | ~\190GAT(27) ,
  \654GAT(229)  = ~\595GAT(198)  | ~\594GAT(206) ,
  \394GAT(143)  = ~\314GAT(79)  | ~\1GAT(0) ,
  \1331GAT(572)  = \1299GAT(540) ,
  \695GAT(260)  = ~\672GAT(247)  | ~\612GAT(238) ,
  \248GAT(46)  = \233GAT(40)  & \227GAT(34) ,
  \1241GAT(480)  = ~\1150GAT(452)  | ~\1054GAT(416) ,
  \1298GAT(544)  = ~\1241GAT(480)  | ~\1240GAT(516) ,
  \1216GAT(430)  = ~\1120GAT(410)  | ~\197GAT(28) ,
  \564GAT(179)  = ~\513GAT(147)  | ~\510GAT(155) ,
  \678GAT(244)  = ~\627GAT(231)  | ~\622GAT(232) ,
  \1327GAT(571)  = \1295GAT(539) ,
  \555GAT(185)  = ~\495GAT(161)  | ~\492GAT(169) ,
  \278GAT(72)  = ~\64GAT(9)  | ~\57GAT(8) ,
  \834GAT(336)  = ~\819GAT(320)  | ~\818GAT(328) ,
  \776GAT(302)  = ~\759GAT(291)  | ~\758GAT(286) ,
  \1337GAT(582)  = \1305GAT(550) ,
  \1297GAT(548)  = ~\1239GAT(484)  | ~\1238GAT(517) ,
  \254GAT(44)  = \233GAT(40)  & \229GAT(36) ,
  \257GAT(43)  = \233GAT(40)  & \230GAT(37) ,
  \702GAT(256)  = ~\684GAT(243)  | ~\622GAT(232) ,
  \571GAT(223)  = ~\522GAT(192)  | ~\429GAT(175) ,
  \350GAT(60)  = ~\155GAT(22)  | ~\127GAT(18) ,
  \275GAT(73)  = ~\50GAT(7)  | ~\43GAT(6) ,
  \242GAT(48)  = \233GAT(40)  & \225GAT(32) ,
  \1343GAT(555)  = \1311GAT(523) ,
  \847GAT(335)  = ~\821GAT(319)  | ~\820GAT(327) ,
  \1147GAT(453)  = ~\1051GAT(420)  | ~\36GAT(5) ,
  \956GAT(353)  = ~\925GAT(332) ,
  \1336GAT(586)  = \1304GAT(554) ,
  \384GAT(100)  = ~\299GAT(57)  | ~\155GAT(22) ,
  \687GAT(242)  = ~\637GAT(226)  | ~\627GAT(231) ,
  \1258GAT(507)  = ~\1177GAT(443)  | ~\106GAT(15) ,
  \1276GAT(498)  = ~\1204GAT(434)  | ~\169GAT(24) ,
  \522GAT(192)  = ~\429GAT(175)  | ~\426GAT(176) ,
  \1320GAT(538)  = ~\1285GAT(474)  | ~\1284GAT(494) ,
  \1286GAT(493)  = ~\1219GAT(429)  | ~\204GAT(29) ,
  \1189GAT(439)  = ~\1093GAT(395)  | ~\134GAT(19) ,
  \951GAT(337)  = ~\899GAT(329) ,
  \950GAT(347)  = ~\886GAT(331) ,
  \1323GAT(526)  = ~\1291GAT(462)  | ~\1290GAT(491) ,
  \1345GAT(564)  = \1313GAT(532) ,
  \657GAT(228)  = ~\597GAT(196)  | ~\596GAT(204) ,
  \1231GAT(483)  = ~\1135GAT(457)  | ~\1039GAT(419) ,
  \899GAT(329)  = ~\833GAT(313)  | ~\832GAT(321) ,
  \1344GAT(568)  = \1312GAT(536) ,
  \694GAT(264)  = ~\672GAT(247)  | ~\602GAT(240) ,
  \405GAT(115)  = ~\329GAT(68)  | ~\99GAT(14) ,
  \1250GAT(511)  = ~\1165GAT(447)  | ~\78GAT(11) ,
  \825GAT(317)  = ~\803GAT(309)  | ~\779GAT(301) ,
  \570GAT(224)  = ~\522GAT(192)  | ~\426GAT(176) ,
  \375GAT(118)  = ~\284GAT(66)  | ~\92GAT(13) ,
  \404GAT(123)  = ~\329GAT(68)  | ~\71GAT(10) ,
  \367GAT(134)  = ~\272GAT(74)  | ~\36GAT(5) ,
  \1334GAT(577)  = \1302GAT(545) ,
  \407GAT(129)  = ~\332GAT(75)  | ~\50GAT(7) ,
  \1247GAT(485)  = ~\1159GAT(449)  | ~\1063GAT(421) ,
  \715GAT(270)  = ~\697GAT(258)  | ~\696GAT(262) ,
  \1237GAT(488)  = ~\1144GAT(454)  | ~\1048GAT(424) ,
  \1138GAT(456)  = ~\1042GAT(415)  | ~\15GAT(2) ,
  \763GAT(296)  = ~\742GAT(276)  | ~\706GAT(272) ,
  \1075GAT(422)  = \1011GAT(388)  & \847GAT(335) ,
  \1290GAT(491)  = ~\1225GAT(427)  | ~\218GAT(31) ,
  \1325GAT(579)  = \1293GAT(547) ,
  \284GAT(66)  = ~\92GAT(13)  | ~\85GAT(12) ,
  \444GAT(165)  = ~\375GAT(118)  | ~\374GAT(120) ,
  \510GAT(155)  = ~\419GAT(99)  | ~\418GAT(107) ,
  \597GAT(196)  = ~\561GAT(180)  | ~\507GAT(148) ,
  \1159GAT(449)  = ~\1063GAT(421)  | ~\64GAT(9) ,
  \374GAT(120)  = ~\284GAT(66)  | ~\85GAT(12) ,
  \967GAT(351)  = ~\886GAT(331) ,
  \794GAT(312)  = ~\770GAT(304)  | ~\642GAT(237) ,
  \824GAT(325)  = ~\803GAT(309)  | ~\651GAT(233) ,
  \1280GAT(496)  = ~\1210GAT(432)  | ~\183GAT(26) ,
  \1099GAT(404)  = \1021GAT(391)  & \886GAT(331) ,
  \703GAT(252)  = ~\684GAT(243)  | ~\632GAT(230) ,
  \1268GAT(502)  = ~\1192GAT(438)  | ~\141GAT(20) ,
  \1207GAT(433)  = ~\1111GAT(405)  | ~\176GAT(25) ,
  \1352GAT(570)  = \1320GAT(538) ,
  \960GAT(344)  = ~\912GAT(330) ,
  \1054GAT(416)  = \1001GAT(387)  & \860GAT(334) ,
  \1123GAT(406)  = \1031GAT(392)  & \886GAT(331) ,
  \266GAT(80)  = ~\8GAT(1)  | ~\1GAT(0) ,
  \704GAT(254)  = ~\687GAT(242)  | ~\627GAT(231) ,
  \1168GAT(446)  = ~\1072GAT(426)  | ~\85GAT(12) ,
  \706GAT(272)  = ~\691GAT(261)  | ~\690GAT(263) ,
  \745GAT(275)  = ~\709GAT(269)  | ~\257GAT(43) ,
  \1321GAT(534)  = ~\1287GAT(470)  | ~\1286GAT(493) ,
  \376GAT(116)  = ~\287GAT(65)  | ~\99GAT(14) ,
  \958GAT(354)  = ~\925GAT(332) ,
  \697GAT(258)  = ~\675GAT(246)  | ~\617GAT(234) ,
  \287GAT(65)  = ~\106GAT(15)  | ~\99GAT(14) ,
  \940GAT(362)  = ~\860GAT(334) ,
  \675GAT(246)  = ~\617GAT(234)  | ~\607GAT(239) ,
  \1324GAT(583)  = \1292GAT(551) ,
  \573GAT(218)  = ~\525GAT(191)  | ~\435GAT(170) ,
  \281GAT(69)  = ~\78GAT(11)  | ~\71GAT(10) ,
  \365GAT(138)  = ~\269GAT(77)  | ~\22GAT(3) ,
  \660GAT(227)  = ~\599GAT(195)  | ~\598GAT(203) ,
  \1351GAT(557)  = \1319GAT(525) ,
  \468GAT(149)  = ~\391GAT(86)  | ~\390GAT(88) ,
  \1292GAT(551)  = ~\1229GAT(487)  | ~\1228GAT(522) ,
  \1245GAT(489)  = ~\1156GAT(450)  | ~\1060GAT(425) ,
  \402GAT(139)  = ~\326GAT(76)  | ~\15GAT(2) ,
  \435GAT(170)  = ~\369GAT(130)  | ~\368GAT(132) ,
  \311GAT(49)  = ~\218GAT(31)  | ~\211GAT(30) ,
  \447GAT(162)  = ~\377GAT(114)  | ~\376GAT(116) ,
  \269GAT(77)  = ~\22GAT(3)  | ~\15GAT(2) ,
  \1259GAT(478)  = ~\1177GAT(443)  | ~\1081GAT(414) ,
  \705GAT(250)  = ~\687GAT(242)  | ~\637GAT(226) ,
  \718GAT(268)  = ~\699GAT(253)  | ~\698GAT(255) ,
  \572GAT(221)  = ~\525GAT(191)  | ~\432GAT(173) ,
  \1204GAT(434)  = ~\1108GAT(409)  | ~\169GAT(24) ,
  \1350GAT(561)  = \1318GAT(529) ,
  \1016GAT(393)  = \991GAT(385)  & (\971GAT(360)  & (\860GAT(334)  & (\970GAT(370)  & \834GAT(336) ))),
  \364GAT(140)  = ~\269GAT(77)  | ~\15GAT(2) ,
  \831GAT(314)  = ~\812GAT(306)  | ~\788GAT(298) ,
  \1269GAT(472)  = ~\1192GAT(438)  | ~\1096GAT(408) ,
  \979GAT(382)  = \943GAT(357)  & (\860GAT(334)  & (\942GAT(368)  & \941GAT(373) )),
  \492GAT(169)  = ~\407GAT(129)  | ~\406GAT(137) ,
  \1335GAT(573)  = \1303GAT(541) ,
  \1347GAT(556)  = \1315GAT(524) ,
  \1295GAT(539)  = ~\1235GAT(475)  | ~\1234GAT(519) ,
  \1186GAT(440)  = ~\1090GAT(399)  | ~\127GAT(18) ,
  \830GAT(322)  = ~\812GAT(306)  | ~\660GAT(227) ,
  \1177GAT(443)  = ~\1081GAT(414)  | ~\106GAT(15) ,
  \1252GAT(510)  = ~\1168GAT(446)  | ~\85GAT(12) ,
  \827GAT(316)  = ~\806GAT(308)  | ~\782GAT(300) ,
  \1238GAT(517)  = ~\1147GAT(453)  | ~\36GAT(5) ,
  \696GAT(262)  = ~\675GAT(246)  | ~\607GAT(239) ,
  \1066GAT(417)  = \1006GAT(390)  & \860GAT(334) ,
  \701GAT(249)  = ~\681GAT(241)  | ~\637GAT(226) ,
  \684GAT(243)  = ~\632GAT(230)  | ~\622GAT(232) ,
  \1346GAT(560)  = \1314GAT(528) ,
  \942GAT(368)  = ~\847GAT(335) ,
  \584GAT(197)  = ~\543GAT(178)  | ~\468GAT(149) ,
  \1293GAT(547)  = ~\1231GAT(483)  | ~\1230GAT(521) ,
  \809GAT(307)  = ~\785GAT(299)  | ~\657GAT(228) ,
  \943GAT(357)  = ~\873GAT(333) ,
  \1026GAT(394)  = \991GAT(385)  & (\975GAT(361)  & (\860GAT(334)  & (\847GAT(335)  & \974GAT(375) ))),
  \296GAT(58)  = ~\148GAT(21)  | ~\141GAT(20) ,
  \1353GAT(566)  = \1321GAT(534) ,
  \978GAT(381)  = \873GAT(333)  & (\940GAT(362)  & (\939GAT(367)  & \938GAT(372) )),
  \371GAT(126)  = ~\278GAT(72)  | ~\64GAT(9) ,
  \363GAT(142)  = ~\266GAT(80)  | ~\8GAT(1) ,
  \401GAT(117)  = ~\323GAT(70)  | ~\92GAT(13) ,
  \826GAT(324)  = ~\806GAT(308)  | ~\654GAT(229) ,
  \299GAT(57)  = ~\162GAT(23)  | ~\155GAT(22) ,
  \495GAT(161)  = ~\409GAT(113)  | ~\408GAT(121) ,
  \377GAT(114)  = ~\287GAT(65)  | ~\106GAT(15) ,
  \1294GAT(543)  = ~\1233GAT(479)  | ~\1232GAT(520) ,
  \762GAT(284)  = ~\742GAT(276)  | ~\254GAT(44) ,
  \1195GAT(437)  = ~\1099GAT(404)  | ~\148GAT(21) ,
  \698GAT(255)  = ~\678GAT(244)  | ~\622GAT(232) ,
  \543GAT(178)  = ~\471GAT(146)  | ~\468GAT(149) ,
  \663GAT(225)  = ~\601GAT(193)  | ~\600GAT(201) ,
  \403GAT(131)  = ~\326GAT(76)  | ~\43GAT(6) ,
  \1213GAT(431)  = ~\1117GAT(397)  | ~\190GAT(27) ,
  \422GAT(105)  = ~\356GAT(59)  | ~\134GAT(19) ,
  \438GAT(168)  = ~\371GAT(126)  | ~\370GAT(128) ,
  \582GAT(200)  = ~\540GAT(182)  | ~\462GAT(152) ,
  \1192GAT(438)  = ~\1096GAT(408)  | ~\141GAT(20) ,
  \797GAT(311)  = ~\773GAT(303)  | ~\645GAT(236) ,
  \941GAT(373)  = ~\834GAT(336) ,
  \513GAT(147)  = ~\421GAT(83)  | ~\420GAT(91) ,
  \821GAT(319)  = ~\797GAT(311)  | ~\773GAT(303) ,
  \1228GAT(522)  = ~\1132GAT(458)  | ~\1GAT(0) ,
  \1039GAT(419)  = \996GAT(389)  & \847GAT(335) ,
  \400GAT(125)  = ~\323GAT(70)  | ~\64GAT(9) ,
  \450GAT(160)  = ~\379GAT(110)  | ~\378GAT(112) ,
  \820GAT(327)  = ~\797GAT(311)  | ~\645GAT(236) ,
  \1282GAT(495)  = ~\1213GAT(431)  | ~\190GAT(27) ,
  \531GAT(186)  = ~\447GAT(162)  | ~\444GAT(165) ,
  \1048GAT(424)  = \1001GAT(387)  & \834GAT(336) ,
  \370GAT(128)  = ~\278GAT(72)  | ~\57GAT(8) ,
  \362GAT(144)  = ~\266GAT(80)  | ~\1GAT(0) ,
  \945GAT(363)  = ~\860GAT(334) ,
  \672GAT(247)  = ~\612GAT(238)  | ~\602GAT(240) ,
  \1150GAT(452)  = ~\1054GAT(416)  | ~\43GAT(6) ,
  \1031GAT(392)  = \991GAT(385)  & (\873GAT(333)  & (\977GAT(366)  & (\847GAT(335)  & \976GAT(376) ))),
  \411GAT(103)  = ~\338GAT(63)  | ~\141GAT(20) ,
  \1349GAT(565)  = \1317GAT(533) ,
  \600GAT(201)  = ~\567GAT(177)  | ~\516GAT(153) ,
  \779GAT(301)  = ~\761GAT(290)  | ~\760GAT(285) ,
  \832GAT(321)  = ~\815GAT(305)  | ~\663GAT(225) ,
  \290GAT(64)  = ~\120GAT(17)  | ~\113GAT(16) ,
  \1248GAT(512)  = ~\1162GAT(448)  | ~\71GAT(10) ,
  \1006GAT(390)  = \986GAT(386)  & (\955GAT(338)  & (\912GAT(330)  & (\886GAT(331)  & \954GAT(352) ))),
  \558GAT(181)  = ~\501GAT(150)  | ~\498GAT(158) ,
  \293GAT(61)  = ~\134GAT(19)  | ~\127GAT(18) ,
  \1102GAT(400)  = \1021GAT(391)  & \912GAT(330) ,
  \1081GAT(414)  = \1011GAT(388)  & \873GAT(333) ,
  \1348GAT(569)  = \1316GAT(537) ,
  \596GAT(204)  = ~\561GAT(180)  | ~\504GAT(156) ,
  \912GAT(330)  = ~\831GAT(314)  | ~\830GAT(322) ,
  \1117GAT(397)  = \1026GAT(394)  & \899GAT(329) ,
  \1235GAT(475)  = ~\1141GAT(455)  | ~\1045GAT(411) ,
  \1222GAT(428)  = ~\1126GAT(402)  | ~\211GAT(30) ,
  \1329GAT(580)  = \1297GAT(548) ,
  \833GAT(313)  = ~\815GAT(305)  | ~\791GAT(297) ,
  \1165GAT(447)  = ~\1069GAT(413)  | ~\78GAT(11) ,
  \648GAT(235)  = ~\591GAT(211)  | ~\590GAT(219) ,
  \699GAT(253)  = ~\678GAT(244)  | ~\627GAT(231) ,
  \1105GAT(396)  = \1021GAT(391)  & \899GAT(329) ,
  \585GAT(194)  = ~\543GAT(178)  | ~\471GAT(146) ,
  \1338GAT(578)  = \1306GAT(546) ,
  \800GAT(310)  = ~\776GAT(302)  | ~\648GAT(235) ,
  \681GAT(241)  = ~\637GAT(226)  | ~\632GAT(230) ,
  \709GAT(269)  = ~\693GAT(257)  | ~\692GAT(259) ,
  \748GAT(274)  = ~\712GAT(271)  | ~\260GAT(42) ,
  \1111GAT(405)  = \1026GAT(394)  & \886GAT(331) ,
  \1183GAT(441)  = ~\1087GAT(403)  | ~\120GAT(17) ,
  \528GAT(190)  = ~\441GAT(167)  | ~\438GAT(168) ,
  \581GAT(202)  = ~\537GAT(183)  | ~\459GAT(154) ,
  \1210GAT(432)  = ~\1114GAT(401)  | ~\183GAT(26) ,
  \947GAT(369)  = ~\847GAT(335) ,
  \1051GAT(420)  = \1001GAT(387)  & \847GAT(335) ,
  \925GAT(332)  = ~\827GAT(316)  | ~\826GAT(324) ,
  \1355GAT(558)  = \1323GAT(526) ,
  \946GAT(358)  = ~\873GAT(333) ,
  \1057GAT(412)  = \1001GAT(387)  & \873GAT(333) ,
  \507GAT(148)  = ~\417GAT(85)  | ~\416GAT(93) ,
  \453GAT(159)  = ~\381GAT(106)  | ~\380GAT(108) ,
  \392GAT(84)  = ~\311GAT(49)  | ~\211GAT(30) ,
  \1291GAT(462)  = ~\1225GAT(427)  | ~\1129GAT(398) ,
  \760GAT(285)  = ~\739GAT(277)  | ~\251GAT(45) ,
  \651GAT(233)  = ~\593GAT(209)  | ~\592GAT(217) ,
  \386GAT(96)  = ~\302GAT(56)  | ~\169GAT(24) ,
  \393GAT(82)  = ~\311GAT(49)  | ~\218GAT(31) ,
  \385GAT(98)  = ~\299GAT(57)  | ~\162GAT(23) ,
  \1174GAT(444)  = ~\1078GAT(418)  | ~\99GAT(14) ,
  \757GAT(289)  = ~\733GAT(279)  | ~\721GAT(265) ,
  \429GAT(175)  = ~\365GAT(138)  | ~\364GAT(140) ,
  \1060GAT(425)  = \1006GAT(390)  & \834GAT(336) ,
  \412GAT(95)  = ~\341GAT(55)  | ~\169GAT(24) ,
  \1021GAT(391)  = \991GAT(385)  & (\873GAT(333)  & (\973GAT(365)  & (\972GAT(371)  & \834GAT(336) ))),
  \1328GAT(584)  = \1296GAT(552) ,
  \739GAT(277)  = ~\727GAT(266)  | ~\251GAT(45) ,
  \1296GAT(552)  = ~\1237GAT(488)  | ~\1236GAT(518) ,
  \594GAT(206)  = ~\558GAT(181)  | ~\498GAT(158) ,
  \373GAT(122)  = ~\281GAT(69)  | ~\78GAT(11) ,
  \823GAT(318)  = ~\800GAT(310)  | ~\776GAT(302) ,
  \388GAT(92)  = ~\305GAT(53)  | ~\183GAT(26) ,
  \580GAT(205)  = ~\537GAT(183)  | ~\456GAT(157) ,
  \1281GAT(465)  = ~\1210GAT(432)  | ~\1114GAT(401) ,
  \537GAT(183)  = ~\459GAT(154)  | ~\456GAT(157) ,
  \1271GAT(468)  = ~\1195GAT(437)  | ~\1099GAT(404) ,
  \462GAT(152)  = ~\387GAT(94)  | ~\386GAT(96) ,
  \627GAT(231)  = ~\581GAT(202)  | ~\580GAT(205) ,
  \822GAT(326)  = ~\800GAT(310)  | ~\648GAT(235) ,
  \944GAT(374)  = ~\834GAT(336) ,
  \1319GAT(525)  = ~\1283GAT(461)  | ~\1282GAT(495) ,
  \419GAT(99)  = ~\350GAT(60)  | ~\155GAT(22) ,
  \1354GAT(562)  = \1322GAT(530) ,
  \391GAT(86)  = ~\308GAT(50)  | ~\204GAT(29) ,
  \387GAT(94)  = ~\302GAT(56)  | ~\176GAT(25) ,
  \751GAT(273)  = ~\715GAT(270)  | ~\263GAT(41) ,
  \390GAT(88)  = ~\308GAT(50)  | ~\197GAT(28) ,
  \1318GAT(529)  = ~\1281GAT(465)  | ~\1280GAT(496) ,
  \389GAT(90)  = ~\305GAT(53)  | ~\190GAT(27) ,
  \540GAT(182)  = ~\465GAT(151)  | ~\462GAT(152) ,
  \788GAT(298)  = ~\767GAT(295)  | ~\766GAT(282) ,
  \1072GAT(426)  = \1011GAT(388)  & \834GAT(336) ,
  \1063GAT(421)  = \1006GAT(390)  & \847GAT(335) ,
  \1339GAT(574)  = \1307GAT(542) ,
  \516GAT(153)  = ~\423GAT(97)  | ~\422GAT(105) ,
  \1262GAT(505)  = ~\1183GAT(441)  | ~\120GAT(17) ,
  \1234GAT(519)  = ~\1141GAT(455)  | ~\22GAT(3) ,
  \1249GAT(481)  = ~\1162GAT(448)  | ~\1066GAT(417) ,
  \416GAT(93)  = ~\347GAT(54)  | ~\176GAT(25) ,
  \939GAT(367)  = ~\847GAT(335) ,
  \1201GAT(435)  = ~\1105GAT(396)  | ~\162GAT(23) ,
  \1153GAT(451)  = ~\1057GAT(412)  | ~\50GAT(7) ,
  \372GAT(124)  = ~\281GAT(69)  | ~\71GAT(10) ,
  \546GAT(189)  = ~\477GAT(166)  | ~\474GAT(174) ,
  \769GAT(294)  = ~\751GAT(273)  | ~\715GAT(270) ,
  \756GAT(287)  = ~\733GAT(279)  | ~\245GAT(47) ,
  \501GAT(150)  = ~\413GAT(87)  | ~\412GAT(95) ,
  \1162GAT(448)  = ~\1066GAT(417)  | ~\71GAT(10) ,
  \1253GAT(490)  = ~\1168GAT(446)  | ~\1072GAT(426) ,
  \498GAT(158)  = ~\411GAT(103)  | ~\410GAT(111) ,
  \766GAT(282)  = ~\748GAT(274)  | ~\260GAT(42) ,
  \617GAT(234)  = ~\577GAT(210)  | ~\576GAT(213) ,
  \886GAT(331)  = ~\829GAT(315)  | ~\828GAT(323) ,
  \959GAT(349)  = ~\886GAT(331) ,
  \1272GAT(500)  = ~\1198GAT(436)  | ~\155GAT(22) ,
  \420GAT(91)  = ~\353GAT(52)  | ~\183GAT(26) ,
  \759GAT(291)  = ~\736GAT(278)  | ~\724GAT(267) ;
endmodule

