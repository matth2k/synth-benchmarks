module s38417 (
  CK,
  g1249,
  g1943,
  g2637,
  g3212,
  g3213,
  g3214,
  g3215,
  g3216,
  g3217,
  g3218,
  g3219,
  g3220,
  g3221,
  g3222,
  g3223,
  g3224,
  g3225,
  g3226,
  g3227,
  g3228,
  g3229,
  g3230,
  g3231,
  g3232,
  g3233,
  g3234,
  g51,
  g563,
  g4590,
  g25420,
  g25442,
  g25489,
  g8021,
  g7334,
  g24734,
  g8258,
  g8273,
  g5437,
  g5472,
  g5511,
  g5555,
  g6231,
  g6368,
  g6573,
  g6837,
  g7909,
  g7961,
  g8012,
  g8087,
  g8261,
  g8023,
  g26104,
  g5629,
  g5657,
  g5695,
  g5747,
  g6485,
  g6677,
  g6750,
  g6979,
  g7052,
  g7229,
  g7302,
  g7425,
  g8106,
  g8096,
  g3993,
  g8259,
  g4088,
  g16355,
  g8249,
  g16496,
  g16437,
  g8251,
  g4090,
  g6442,
  g8266,
  g8271,
  g4323,
  g8263,
  g4321,
  g4450,
  g16297,
  g8267,
  g8275,
  g4200,
  g8269,
  g7519,
  g16399,
  g25435,
  g5549,
  g5595,
  g5612,
  g5637,
  g8274,
  g6225,
  g8270,
  g8264,
  g8272,
  g5648,
  g5686,
  g5738,
  g5796,
  g6642,
  g6911,
  g6944,
  g7161,
  g7194,
  g7357,
  g7390,
  g7487,
  g8030,
  g8268,
  g26149,
  g5388,
  g8265,
  g27380,
  g6313,
  g6447,
  g6518,
  g6712,
  g6782,
  g7014,
  g7084,
  g7264,
  g7956,
  g8007,
  g8082,
  g8167,
  g26135,
  g8262,
  g8260,
  g6895,
  g8175
);
  input CK;
  wire CK;
  input g1249;
  wire g1249;
  input g1943;
  wire g1943;
  input g2637;
  wire g2637;
  input g3212;
  wire g3212;
  input g3213;
  wire g3213;
  input g3214;
  wire g3214;
  input g3215;
  wire g3215;
  input g3216;
  wire g3216;
  input g3217;
  wire g3217;
  input g3218;
  wire g3218;
  input g3219;
  wire g3219;
  input g3220;
  wire g3220;
  input g3221;
  wire g3221;
  input g3222;
  wire g3222;
  input g3223;
  wire g3223;
  input g3224;
  wire g3224;
  input g3225;
  wire g3225;
  input g3226;
  wire g3226;
  input g3227;
  wire g3227;
  input g3228;
  wire g3228;
  input g3229;
  wire g3229;
  input g3230;
  wire g3230;
  input g3231;
  wire g3231;
  input g3232;
  wire g3232;
  input g3233;
  wire g3233;
  input g3234;
  wire g3234;
  input g51;
  wire g51;
  input g563;
  wire g563;
  output g4590;
  wire g4590;
  output g25420;
  wire g25420;
  output g25442;
  wire g25442;
  output g25489;
  wire g25489;
  output g8021;
  wire g8021;
  output g7334;
  wire g7334;
  output g24734;
  wire g24734;
  output g8258;
  wire g8258;
  output g8273;
  wire g8273;
  output g5437;
  wire g5437;
  output g5472;
  wire g5472;
  output g5511;
  wire g5511;
  output g5555;
  wire g5555;
  output g6231;
  wire g6231;
  output g6368;
  wire g6368;
  output g6573;
  wire g6573;
  output g6837;
  wire g6837;
  output g7909;
  wire g7909;
  output g7961;
  wire g7961;
  output g8012;
  wire g8012;
  output g8087;
  wire g8087;
  output g8261;
  wire g8261;
  output g8023;
  wire g8023;
  output g26104;
  wire g26104;
  output g5629;
  wire g5629;
  output g5657;
  wire g5657;
  output g5695;
  wire g5695;
  output g5747;
  wire g5747;
  output g6485;
  wire g6485;
  output g6677;
  wire g6677;
  output g6750;
  wire g6750;
  output g6979;
  wire g6979;
  output g7052;
  wire g7052;
  output g7229;
  wire g7229;
  output g7302;
  wire g7302;
  output g7425;
  wire g7425;
  output g8106;
  wire g8106;
  output g8096;
  wire g8096;
  output g3993;
  wire g3993;
  output g8259;
  wire g8259;
  output g4088;
  wire g4088;
  output g16355;
  wire g16355;
  output g8249;
  wire g8249;
  output g16496;
  wire g16496;
  output g16437;
  wire g16437;
  output g8251;
  wire g8251;
  output g4090;
  wire g4090;
  output g6442;
  wire g6442;
  output g8266;
  wire g8266;
  output g8271;
  wire g8271;
  output g4323;
  wire g4323;
  output g8263;
  wire g8263;
  output g4321;
  wire g4321;
  output g4450;
  wire g4450;
  output g16297;
  wire g16297;
  output g8267;
  wire g8267;
  output g8275;
  wire g8275;
  output g4200;
  wire g4200;
  output g8269;
  wire g8269;
  output g7519;
  wire g7519;
  output g16399;
  wire g16399;
  output g25435;
  wire g25435;
  output g5549;
  wire g5549;
  output g5595;
  wire g5595;
  output g5612;
  wire g5612;
  output g5637;
  wire g5637;
  output g8274;
  wire g8274;
  output g6225;
  wire g6225;
  output g8270;
  wire g8270;
  output g8264;
  wire g8264;
  output g8272;
  wire g8272;
  output g5648;
  wire g5648;
  output g5686;
  wire g5686;
  output g5738;
  wire g5738;
  output g5796;
  wire g5796;
  output g6642;
  wire g6642;
  output g6911;
  wire g6911;
  output g6944;
  wire g6944;
  output g7161;
  wire g7161;
  output g7194;
  wire g7194;
  output g7357;
  wire g7357;
  output g7390;
  wire g7390;
  output g7487;
  wire g7487;
  output g8030;
  wire g8030;
  output g8268;
  wire g8268;
  output g26149;
  wire g26149;
  output g5388;
  wire g5388;
  output g8265;
  wire g8265;
  output g27380;
  wire g27380;
  output g6313;
  wire g6313;
  output g6447;
  wire g6447;
  output g6518;
  wire g6518;
  output g6712;
  wire g6712;
  output g6782;
  wire g6782;
  output g7014;
  wire g7014;
  output g7084;
  wire g7084;
  output g7264;
  wire g7264;
  output g7956;
  wire g7956;
  output g8007;
  wire g8007;
  output g8082;
  wire g8082;
  output g8167;
  wire g8167;
  output g26135;
  wire g26135;
  output g8262;
  wire g8262;
  output g8260;
  wire g8260;
  output g6895;
  wire g6895;
  output g8175;
  wire g8175;
  wire __0__;
  wire __1__;
  wire __2__;
  wire __3__;
  wire __4__;
  wire __5__;
  wire __6__;
  wire __7__;
  wire __8__;
  wire __9__;
  wire __10__;
  wire __11__;
  wire __12__;
  wire __13__;
  wire __14__;
  wire __15__;
  wire __16__;
  wire __17__;
  wire __18__;
  wire __19__;
  wire __20__;
  wire __21__;
  wire __22__;
  wire __23__;
  wire __24__;
  wire __25__;
  wire __26__;
  wire __27__;
  wire __28__;
  wire __29__;
  wire __30__;
  wire __31__;
  wire __32__;
  wire __33__;
  wire __34__;
  wire __35__;
  wire __36__;
  wire __37__;
  wire __38__;
  wire __39__;
  wire __40__;
  wire __41__;
  wire __42__;
  wire __43__;
  wire __44__;
  wire __45__;
  wire __46__;
  wire __47__;
  wire __48__;
  wire __49__;
  wire __50__;
  wire __51__;
  wire __52__;
  wire __53__;
  wire __54__;
  wire __55__;
  wire __56__;
  wire __57__;
  wire __58__;
  wire __59__;
  wire __60__;
  wire __61__;
  wire __62__;
  wire __63__;
  wire __64__;
  wire __65__;
  wire __66__;
  wire __67__;
  wire __68__;
  wire __69__;
  wire __70__;
  wire __71__;
  wire __72__;
  wire __73__;
  wire __74__;
  wire __75__;
  wire __76__;
  wire __77__;
  wire __78__;
  wire __79__;
  wire __80__;
  wire __81__;
  wire __82__;
  wire __83__;
  wire __84__;
  wire __85__;
  wire __86__;
  wire __87__;
  wire __88__;
  wire __89__;
  wire __90__;
  wire __91__;
  wire __92__;
  wire __93__;
  wire __94__;
  wire __95__;
  wire __96__;
  wire __97__;
  wire __98__;
  wire __99__;
  wire __100__;
  wire __101__;
  wire __102__;
  wire __103__;
  wire __104__;
  wire __105__;
  wire __106__;
  wire __107__;
  wire __108__;
  wire __109__;
  wire __110__;
  wire __111__;
  wire __112__;
  wire __113__;
  wire __114__;
  wire __115__;
  wire __116__;
  wire __117__;
  wire __118__;
  wire __119__;
  wire __120__;
  wire __121__;
  wire __122__;
  wire __123__;
  wire __124__;
  wire __125__;
  wire __126__;
  wire __127__;
  wire __128__;
  wire __129__;
  wire __130__;
  wire __131__;
  wire __132__;
  wire __133__;
  wire __134__;
  wire __135__;
  wire __136__;
  wire __137__;
  wire __138__;
  wire __139__;
  wire __140__;
  wire __141__;
  wire __142__;
  wire __143__;
  wire __144__;
  wire __145__;
  wire __146__;
  wire __147__;
  wire __148__;
  wire __149__;
  wire __150__;
  wire __151__;
  wire __152__;
  wire __153__;
  wire __154__;
  wire __155__;
  wire __156__;
  wire __157__;
  wire __158__;
  wire __159__;
  wire __160__;
  wire __161__;
  wire __162__;
  wire __163__;
  wire __164__;
  wire __165__;
  wire __166__;
  wire __167__;
  wire __168__;
  wire __169__;
  wire __170__;
  wire __171__;
  wire __172__;
  wire __173__;
  wire __174__;
  wire __175__;
  wire __176__;
  wire __177__;
  wire __178__;
  wire __179__;
  wire __180__;
  wire __181__;
  wire __182__;
  wire __183__;
  wire __184__;
  wire __185__;
  wire __186__;
  wire __187__;
  wire __188__;
  wire __189__;
  wire __190__;
  wire __191__;
  wire __192__;
  wire __193__;
  wire __194__;
  wire __195__;
  wire __196__;
  wire __197__;
  wire __198__;
  wire __199__;
  wire __200__;
  wire __201__;
  wire __202__;
  wire __203__;
  wire __204__;
  wire __205__;
  wire __206__;
  wire __207__;
  wire __208__;
  wire __209__;
  wire __210__;
  wire __211__;
  wire __212__;
  wire __213__;
  wire __214__;
  wire __215__;
  wire __216__;
  wire __217__;
  wire __218__;
  wire __219__;
  wire __220__;
  wire __221__;
  wire __222__;
  wire __223__;
  wire __224__;
  wire __225__;
  wire __226__;
  wire __227__;
  wire __228__;
  wire __229__;
  wire __230__;
  wire __231__;
  wire __232__;
  wire __233__;
  wire __234__;
  wire __235__;
  wire __236__;
  wire __237__;
  wire __238__;
  wire __239__;
  wire __240__;
  wire __241__;
  wire __242__;
  wire __243__;
  wire __244__;
  wire __245__;
  wire __246__;
  wire __247__;
  wire __248__;
  wire __249__;
  wire __250__;
  wire __251__;
  wire __252__;
  wire __253__;
  wire __254__;
  wire __255__;
  wire __256__;
  wire __257__;
  wire __258__;
  wire __259__;
  wire __260__;
  wire __261__;
  wire __262__;
  wire __263__;
  wire __264__;
  wire __265__;
  wire __266__;
  wire __267__;
  wire __268__;
  wire __269__;
  wire __270__;
  wire __271__;
  wire __272__;
  wire __273__;
  wire __274__;
  wire __275__;
  wire __276__;
  wire __277__;
  wire __278__;
  wire __279__;
  wire __280__;
  wire __281__;
  wire __282__;
  wire __283__;
  wire __284__;
  wire __285__;
  wire __286__;
  wire __287__;
  wire __288__;
  wire __289__;
  wire __290__;
  wire __291__;
  wire __292__;
  wire __293__;
  wire __294__;
  wire __295__;
  wire __296__;
  wire __297__;
  wire __298__;
  wire __299__;
  wire __300__;
  wire __301__;
  wire __302__;
  wire __303__;
  wire __304__;
  wire __305__;
  wire __306__;
  wire __307__;
  wire __308__;
  wire __309__;
  wire __310__;
  wire __311__;
  wire __312__;
  wire __313__;
  wire __314__;
  wire __315__;
  wire __316__;
  wire __317__;
  wire __318__;
  wire __319__;
  wire __320__;
  wire __321__;
  wire __322__;
  wire __323__;
  wire __324__;
  wire __325__;
  wire __326__;
  wire __327__;
  wire __328__;
  wire __329__;
  wire __330__;
  wire __331__;
  wire __332__;
  wire __333__;
  wire __334__;
  wire __335__;
  wire __336__;
  wire __337__;
  wire __338__;
  wire __339__;
  wire __340__;
  wire __341__;
  wire __342__;
  wire __343__;
  wire __344__;
  wire __345__;
  wire __346__;
  wire __347__;
  wire __348__;
  wire __349__;
  wire __350__;
  wire __351__;
  wire __352__;
  wire __353__;
  wire __354__;
  wire __355__;
  wire __356__;
  wire __357__;
  wire __358__;
  wire __359__;
  wire __360__;
  wire __361__;
  wire __362__;
  wire __363__;
  wire __364__;
  wire __365__;
  wire __366__;
  wire __367__;
  wire __368__;
  wire __369__;
  wire __370__;
  wire __371__;
  wire __372__;
  wire __373__;
  wire __374__;
  wire __375__;
  wire __376__;
  wire __377__;
  wire __378__;
  wire __379__;
  wire __380__;
  wire __381__;
  wire __382__;
  wire __383__;
  wire __384__;
  wire __385__;
  wire __386__;
  wire __387__;
  wire __388__;
  wire __389__;
  wire __390__;
  wire __391__;
  wire __392__;
  wire __393__;
  wire __394__;
  wire __395__;
  wire __396__;
  wire __397__;
  wire __398__;
  wire __399__;
  wire __400__;
  wire __401__;
  wire __402__;
  wire __403__;
  wire __404__;
  wire __405__;
  wire __406__;
  wire __407__;
  wire __408__;
  wire __409__;
  wire __410__;
  wire __411__;
  wire __412__;
  wire __413__;
  wire __414__;
  wire __415__;
  wire __416__;
  wire __417__;
  wire __418__;
  wire __419__;
  wire __420__;
  wire __421__;
  wire __422__;
  wire __423__;
  wire __424__;
  wire __425__;
  wire __426__;
  wire __427__;
  wire __428__;
  wire __429__;
  wire __430__;
  wire __431__;
  wire __432__;
  wire __433__;
  wire __434__;
  wire __435__;
  wire __436__;
  wire __437__;
  wire __438__;
  wire __439__;
  wire __440__;
  wire __441__;
  wire __442__;
  wire __443__;
  wire __444__;
  wire __445__;
  wire __446__;
  wire __447__;
  wire __448__;
  wire __449__;
  wire __450__;
  wire __451__;
  wire __452__;
  wire __453__;
  wire __454__;
  wire __455__;
  wire __456__;
  wire __457__;
  wire __458__;
  wire __459__;
  wire __460__;
  wire __461__;
  wire __462__;
  wire __463__;
  wire __464__;
  wire __465__;
  wire __466__;
  wire __467__;
  wire __468__;
  wire __469__;
  wire __470__;
  wire __471__;
  wire __472__;
  wire __473__;
  wire __474__;
  wire __475__;
  wire __476__;
  wire __477__;
  wire __478__;
  wire __479__;
  wire __480__;
  wire __481__;
  wire __482__;
  wire __483__;
  wire __484__;
  wire __485__;
  wire __486__;
  wire __487__;
  wire __488__;
  wire __489__;
  wire __490__;
  wire __491__;
  wire __492__;
  wire __493__;
  wire __494__;
  wire __495__;
  wire __496__;
  wire __497__;
  wire __498__;
  wire __499__;
  wire __500__;
  wire __501__;
  wire __502__;
  wire __503__;
  wire __504__;
  wire __505__;
  wire __506__;
  wire __507__;
  wire __508__;
  wire __509__;
  wire __510__;
  wire __511__;
  wire __512__;
  wire __513__;
  wire __514__;
  wire __515__;
  wire __516__;
  wire __517__;
  wire __518__;
  wire __519__;
  wire __520__;
  wire __521__;
  wire __522__;
  wire __523__;
  wire __524__;
  wire __525__;
  wire __526__;
  wire __527__;
  wire __528__;
  wire __529__;
  wire __530__;
  wire __531__;
  wire __532__;
  wire __533__;
  wire __534__;
  wire __535__;
  wire __536__;
  wire __537__;
  wire __538__;
  wire __539__;
  wire __540__;
  wire __541__;
  wire __542__;
  wire __543__;
  wire __544__;
  wire __545__;
  wire __546__;
  wire __547__;
  wire __548__;
  wire __549__;
  wire __550__;
  wire __551__;
  wire __552__;
  wire __553__;
  wire __554__;
  wire __555__;
  wire __556__;
  wire __557__;
  wire __558__;
  wire __559__;
  wire __560__;
  wire __561__;
  wire __562__;
  wire __563__;
  wire __564__;
  wire __565__;
  wire __566__;
  wire __567__;
  wire __568__;
  wire __569__;
  wire __570__;
  wire __571__;
  wire __572__;
  wire __573__;
  wire __574__;
  wire __575__;
  wire __576__;
  wire __577__;
  wire __578__;
  wire __579__;
  wire __580__;
  wire __581__;
  wire __582__;
  wire __583__;
  wire __584__;
  wire __585__;
  wire __586__;
  wire __587__;
  wire __588__;
  wire __589__;
  wire __590__;
  wire __591__;
  wire __592__;
  wire __593__;
  wire __594__;
  wire __595__;
  wire __596__;
  wire __597__;
  wire __598__;
  wire __599__;
  wire __600__;
  wire __601__;
  wire __602__;
  wire __603__;
  wire __604__;
  wire __605__;
  wire __606__;
  wire __607__;
  wire __608__;
  wire __609__;
  wire __610__;
  wire __611__;
  wire __612__;
  wire __613__;
  wire __614__;
  wire __615__;
  wire __616__;
  wire __617__;
  wire __618__;
  wire __619__;
  wire __620__;
  wire __621__;
  wire __622__;
  wire __623__;
  wire __624__;
  wire __625__;
  wire __626__;
  wire __627__;
  wire __628__;
  wire __629__;
  wire __630__;
  wire __631__;
  wire __632__;
  wire __633__;
  wire __634__;
  wire __635__;
  wire __636__;
  wire __637__;
  wire __638__;
  wire __639__;
  wire __640__;
  wire __641__;
  wire __642__;
  wire __643__;
  wire __644__;
  wire __645__;
  wire __646__;
  wire __647__;
  wire __648__;
  wire __649__;
  wire __650__;
  wire __651__;
  wire __652__;
  wire __653__;
  wire __654__;
  wire __655__;
  wire __656__;
  wire __657__;
  wire __658__;
  wire __659__;
  wire __660__;
  wire __661__;
  wire __662__;
  wire __663__;
  wire __664__;
  wire __665__;
  wire __666__;
  wire __667__;
  wire __668__;
  wire __669__;
  wire __670__;
  wire __671__;
  wire __672__;
  wire __673__;
  wire __674__;
  wire __675__;
  wire __676__;
  wire __677__;
  wire __678__;
  wire __679__;
  wire __680__;
  wire __681__;
  wire __682__;
  wire __683__;
  wire __684__;
  wire __685__;
  wire __686__;
  wire __687__;
  wire __688__;
  wire __689__;
  wire __690__;
  wire __691__;
  wire __692__;
  wire __693__;
  wire __694__;
  wire __695__;
  wire __696__;
  wire __697__;
  wire __698__;
  wire __699__;
  wire __700__;
  wire __701__;
  wire __702__;
  wire __703__;
  wire __704__;
  wire __705__;
  wire __706__;
  wire __707__;
  wire __708__;
  wire __709__;
  wire __710__;
  wire __711__;
  wire __712__;
  wire __713__;
  wire __714__;
  wire __715__;
  wire __716__;
  wire __717__;
  wire __718__;
  wire __719__;
  wire __720__;
  wire __721__;
  wire __722__;
  wire __723__;
  wire __724__;
  wire __725__;
  wire __726__;
  wire __727__;
  wire __728__;
  wire __729__;
  wire __730__;
  wire __731__;
  wire __732__;
  wire __733__;
  wire __734__;
  wire __735__;
  wire __736__;
  wire __737__;
  wire __738__;
  wire __739__;
  wire __740__;
  wire __741__;
  wire __742__;
  wire __743__;
  wire __744__;
  wire __745__;
  wire __746__;
  wire __747__;
  wire __748__;
  wire __749__;
  wire __750__;
  wire __751__;
  wire __752__;
  wire __753__;
  wire __754__;
  wire __755__;
  wire __756__;
  wire __757__;
  wire __758__;
  wire __759__;
  wire __760__;
  wire __761__;
  wire __762__;
  wire __763__;
  wire __764__;
  wire __765__;
  wire __766__;
  wire __767__;
  wire __768__;
  wire __769__;
  wire __770__;
  wire __771__;
  wire __772__;
  wire __773__;
  wire __774__;
  wire __775__;
  wire __776__;
  wire __777__;
  wire __778__;
  wire __779__;
  wire __780__;
  wire __781__;
  wire __782__;
  wire __783__;
  wire __784__;
  wire __785__;
  wire __786__;
  wire __787__;
  wire __788__;
  wire __789__;
  wire __790__;
  wire __791__;
  wire __792__;
  wire __793__;
  wire __794__;
  wire __795__;
  wire __796__;
  wire __797__;
  wire __798__;
  wire __799__;
  wire __800__;
  wire __801__;
  wire __802__;
  wire __803__;
  wire __804__;
  wire __805__;
  wire __806__;
  wire __807__;
  wire __808__;
  wire __809__;
  wire __810__;
  wire __811__;
  wire __812__;
  wire __813__;
  wire __814__;
  wire __815__;
  wire __816__;
  wire __817__;
  wire __818__;
  wire __819__;
  wire __820__;
  wire __821__;
  wire __822__;
  wire __823__;
  wire __824__;
  wire __825__;
  wire __826__;
  wire __827__;
  wire __828__;
  wire __829__;
  wire __830__;
  wire __831__;
  wire __832__;
  wire __833__;
  wire __834__;
  wire __835__;
  wire __836__;
  wire __837__;
  wire __838__;
  wire __839__;
  wire __840__;
  wire __841__;
  wire __842__;
  wire __843__;
  wire __844__;
  wire __845__;
  wire __846__;
  wire __847__;
  wire __848__;
  wire __849__;
  wire __850__;
  wire __851__;
  wire __852__;
  wire __853__;
  wire __854__;
  wire __855__;
  wire __856__;
  wire __857__;
  wire __858__;
  wire __859__;
  wire __860__;
  wire __861__;
  wire __862__;
  wire __863__;
  wire __864__;
  wire __865__;
  wire __866__;
  wire __867__;
  wire __868__;
  wire __869__;
  wire __870__;
  wire __871__;
  wire __872__;
  wire __873__;
  wire __874__;
  wire __875__;
  wire __876__;
  wire __877__;
  wire __878__;
  wire __879__;
  wire __880__;
  wire __881__;
  wire __882__;
  wire __883__;
  wire __884__;
  wire __885__;
  wire __886__;
  wire __887__;
  wire __888__;
  wire __889__;
  wire __890__;
  wire __891__;
  wire __892__;
  wire __893__;
  wire __894__;
  wire __895__;
  wire __896__;
  wire __897__;
  wire __898__;
  wire __899__;
  wire __900__;
  wire __901__;
  wire __902__;
  wire __903__;
  wire __904__;
  wire __905__;
  wire __906__;
  wire __907__;
  wire __908__;
  wire __909__;
  wire __910__;
  wire __911__;
  wire __912__;
  wire __913__;
  wire __914__;
  wire __915__;
  wire __916__;
  wire __917__;
  wire __918__;
  wire __919__;
  wire __920__;
  wire __921__;
  wire __922__;
  wire __923__;
  wire __924__;
  wire __925__;
  wire __926__;
  wire __927__;
  wire __928__;
  wire __929__;
  wire __930__;
  wire __931__;
  wire __932__;
  wire __933__;
  wire __934__;
  wire __935__;
  wire __936__;
  wire __937__;
  wire __938__;
  wire __939__;
  wire __940__;
  wire __941__;
  wire __942__;
  wire __943__;
  wire __944__;
  wire __945__;
  wire __946__;
  wire __947__;
  wire __948__;
  wire __949__;
  wire __950__;
  wire __951__;
  wire __952__;
  wire __953__;
  wire __954__;
  wire __955__;
  wire __956__;
  wire __957__;
  wire __958__;
  wire __959__;
  wire __960__;
  wire __961__;
  wire __962__;
  wire __963__;
  wire __964__;
  wire __965__;
  wire __966__;
  wire __967__;
  wire __968__;
  wire __969__;
  wire __970__;
  wire __971__;
  wire __972__;
  wire __973__;
  wire __974__;
  wire __975__;
  wire __976__;
  wire __977__;
  wire __978__;
  wire __979__;
  wire __980__;
  wire __981__;
  wire __982__;
  wire __983__;
  wire __984__;
  wire __985__;
  wire __986__;
  wire __987__;
  wire __988__;
  wire __989__;
  wire __990__;
  wire __991__;
  wire __992__;
  wire __993__;
  wire __994__;
  wire __995__;
  wire __996__;
  wire __997__;
  wire __998__;
  wire __999__;
  wire __1000__;
  wire __1001__;
  wire __1002__;
  wire __1003__;
  wire __1004__;
  wire __1005__;
  wire __1006__;
  wire __1007__;
  wire __1008__;
  wire __1009__;
  wire __1010__;
  wire __1011__;
  wire __1012__;
  wire __1013__;
  wire __1014__;
  wire __1015__;
  wire __1016__;
  wire __1017__;
  wire __1018__;
  wire __1019__;
  wire __1020__;
  wire __1021__;
  wire __1022__;
  wire __1023__;
  wire __1024__;
  wire __1025__;
  wire __1026__;
  wire __1027__;
  wire __1028__;
  wire __1029__;
  wire __1030__;
  wire __1031__;
  wire __1032__;
  wire __1033__;
  wire __1034__;
  wire __1035__;
  wire __1036__;
  wire __1037__;
  wire __1038__;
  wire __1039__;
  wire __1040__;
  wire __1041__;
  wire __1042__;
  wire __1043__;
  wire __1044__;
  wire __1045__;
  wire __1046__;
  wire __1047__;
  wire __1048__;
  wire __1049__;
  wire __1050__;
  wire __1051__;
  wire __1052__;
  wire __1053__;
  wire __1054__;
  wire __1055__;
  wire __1056__;
  wire __1057__;
  wire __1058__;
  wire __1059__;
  wire __1060__;
  wire __1061__;
  wire __1062__;
  wire __1063__;
  wire __1064__;
  wire __1065__;
  wire __1066__;
  wire __1067__;
  wire __1068__;
  wire __1069__;
  wire __1070__;
  wire __1071__;
  wire __1072__;
  wire __1073__;
  wire __1074__;
  wire __1075__;
  wire __1076__;
  wire __1077__;
  wire __1078__;
  wire __1079__;
  wire __1080__;
  wire __1081__;
  wire __1082__;
  wire __1083__;
  wire __1084__;
  wire __1085__;
  wire __1086__;
  wire __1087__;
  wire __1088__;
  wire __1089__;
  wire __1090__;
  wire __1091__;
  wire __1092__;
  wire __1093__;
  wire __1094__;
  wire __1095__;
  wire __1096__;
  wire __1097__;
  wire __1098__;
  wire __1099__;
  wire __1100__;
  wire __1101__;
  wire __1102__;
  wire __1103__;
  wire __1104__;
  wire __1105__;
  wire __1106__;
  wire __1107__;
  wire __1108__;
  wire __1109__;
  wire __1110__;
  wire __1111__;
  wire __1112__;
  wire __1113__;
  wire __1114__;
  wire __1115__;
  wire __1116__;
  wire __1117__;
  wire __1118__;
  wire __1119__;
  wire __1120__;
  wire __1121__;
  wire __1122__;
  wire __1123__;
  wire __1124__;
  wire __1125__;
  wire __1126__;
  wire __1127__;
  wire __1128__;
  wire __1129__;
  wire __1130__;
  wire __1131__;
  wire __1132__;
  wire __1133__;
  wire __1134__;
  wire __1135__;
  wire __1136__;
  wire __1137__;
  wire __1138__;
  wire __1139__;
  wire __1140__;
  wire __1141__;
  wire __1142__;
  wire __1143__;
  wire __1144__;
  wire __1145__;
  wire __1146__;
  wire __1147__;
  wire __1148__;
  wire __1149__;
  wire __1150__;
  wire __1151__;
  wire __1152__;
  wire __1153__;
  wire __1154__;
  wire __1155__;
  wire __1156__;
  wire __1157__;
  wire __1158__;
  wire __1159__;
  wire __1160__;
  wire __1161__;
  wire __1162__;
  wire __1163__;
  wire __1164__;
  wire __1165__;
  wire __1166__;
  wire __1167__;
  wire __1168__;
  wire __1169__;
  wire __1170__;
  wire __1171__;
  wire __1172__;
  wire __1173__;
  wire __1174__;
  wire __1175__;
  wire __1176__;
  wire __1177__;
  wire __1178__;
  wire __1179__;
  wire __1180__;
  wire __1181__;
  wire __1182__;
  wire __1183__;
  wire __1184__;
  wire __1185__;
  wire __1186__;
  wire __1187__;
  wire __1188__;
  wire __1189__;
  wire __1190__;
  wire __1191__;
  wire __1192__;
  wire __1193__;
  wire __1194__;
  wire __1195__;
  wire __1196__;
  wire __1197__;
  wire __1198__;
  wire __1199__;
  wire __1200__;
  wire __1201__;
  wire __1202__;
  wire __1203__;
  wire __1204__;
  wire __1205__;
  wire __1206__;
  wire __1207__;
  wire __1208__;
  wire __1209__;
  wire __1210__;
  wire __1211__;
  wire __1212__;
  wire __1213__;
  wire __1214__;
  wire __1215__;
  wire __1216__;
  wire __1217__;
  wire __1218__;
  wire __1219__;
  wire __1220__;
  wire __1221__;
  wire __1222__;
  wire __1223__;
  wire __1224__;
  wire __1225__;
  wire __1226__;
  wire __1227__;
  wire __1228__;
  wire __1229__;
  wire __1230__;
  wire __1231__;
  wire __1232__;
  wire __1233__;
  wire __1234__;
  wire __1235__;
  wire __1236__;
  wire __1237__;
  wire __1238__;
  wire __1239__;
  wire __1240__;
  wire __1241__;
  wire __1242__;
  wire __1243__;
  wire __1244__;
  wire __1245__;
  wire __1246__;
  wire __1247__;
  wire __1248__;
  wire __1249__;
  wire __1250__;
  wire __1251__;
  wire __1252__;
  wire __1253__;
  wire __1254__;
  wire __1255__;
  wire __1256__;
  wire __1257__;
  wire __1258__;
  wire __1259__;
  wire __1260__;
  wire __1261__;
  wire __1262__;
  wire __1263__;
  wire __1264__;
  wire __1265__;
  wire __1266__;
  wire __1267__;
  wire __1268__;
  wire __1269__;
  wire __1270__;
  wire __1271__;
  wire __1272__;
  wire __1273__;
  wire __1274__;
  wire __1275__;
  wire __1276__;
  wire __1277__;
  wire __1278__;
  wire __1279__;
  wire __1280__;
  wire __1281__;
  wire __1282__;
  wire __1283__;
  wire __1284__;
  wire __1285__;
  wire __1286__;
  wire __1287__;
  wire __1288__;
  wire __1289__;
  wire __1290__;
  wire __1291__;
  wire __1292__;
  wire __1293__;
  wire __1294__;
  wire __1295__;
  wire __1296__;
  wire __1297__;
  wire __1298__;
  wire __1299__;
  wire __1300__;
  wire __1301__;
  wire __1302__;
  wire __1303__;
  wire __1304__;
  wire __1305__;
  wire __1306__;
  wire __1307__;
  wire __1308__;
  wire __1309__;
  wire __1310__;
  wire __1311__;
  wire __1312__;
  wire __1313__;
  wire __1314__;
  wire __1315__;
  wire __1316__;
  wire __1317__;
  wire __1318__;
  wire __1319__;
  wire __1320__;
  wire __1321__;
  wire __1322__;
  wire __1323__;
  wire __1324__;
  wire __1325__;
  wire __1326__;
  wire __1327__;
  wire __1328__;
  wire __1329__;
  wire __1330__;
  wire __1331__;
  wire __1332__;
  wire __1333__;
  wire __1334__;
  wire __1335__;
  wire __1336__;
  wire __1337__;
  wire __1338__;
  wire __1339__;
  wire __1340__;
  wire __1341__;
  wire __1342__;
  wire __1343__;
  wire __1344__;
  wire __1345__;
  wire __1346__;
  wire __1347__;
  wire __1348__;
  wire __1349__;
  wire __1350__;
  wire __1351__;
  wire __1352__;
  wire __1353__;
  wire __1354__;
  wire __1355__;
  wire __1356__;
  wire __1357__;
  wire __1358__;
  wire __1359__;
  wire __1360__;
  wire __1361__;
  wire __1362__;
  wire __1363__;
  wire __1364__;
  wire __1365__;
  wire __1366__;
  wire __1367__;
  wire __1368__;
  wire __1369__;
  wire __1370__;
  wire __1371__;
  wire __1372__;
  wire __1373__;
  wire __1374__;
  wire __1375__;
  wire __1376__;
  wire __1377__;
  wire __1378__;
  wire __1379__;
  wire __1380__;
  wire __1381__;
  wire __1382__;
  wire __1383__;
  wire __1384__;
  wire __1385__;
  wire __1386__;
  wire __1387__;
  wire __1388__;
  wire __1389__;
  wire __1390__;
  wire __1391__;
  wire __1392__;
  wire __1393__;
  wire __1394__;
  wire __1395__;
  wire __1396__;
  wire __1397__;
  wire __1398__;
  wire __1399__;
  wire __1400__;
  wire __1401__;
  wire __1402__;
  wire __1403__;
  wire __1404__;
  wire __1405__;
  wire __1406__;
  wire __1407__;
  wire __1408__;
  wire __1409__;
  wire __1410__;
  wire __1411__;
  wire __1412__;
  wire __1413__;
  wire __1414__;
  wire __1415__;
  wire __1416__;
  wire __1417__;
  wire __1418__;
  wire __1419__;
  wire __1420__;
  wire __1421__;
  wire __1422__;
  wire __1423__;
  wire __1424__;
  wire __1425__;
  wire __1426__;
  wire __1427__;
  wire __1428__;
  wire __1429__;
  wire __1430__;
  wire __1431__;
  wire __1432__;
  wire __1433__;
  wire __1434__;
  wire __1435__;
  wire __1436__;
  wire __1437__;
  wire __1438__;
  wire __1439__;
  wire __1440__;
  wire __1441__;
  wire __1442__;
  wire __1443__;
  wire __1444__;
  wire __1445__;
  wire __1446__;
  wire __1447__;
  wire __1448__;
  wire __1449__;
  wire __1450__;
  wire __1451__;
  wire __1452__;
  wire __1453__;
  wire __1454__;
  wire __1455__;
  wire __1456__;
  wire __1457__;
  wire __1458__;
  wire __1459__;
  wire __1460__;
  wire __1461__;
  wire __1462__;
  wire __1463__;
  wire __1464__;
  wire __1465__;
  wire __1466__;
  wire __1467__;
  wire __1468__;
  wire __1469__;
  wire __1470__;
  wire __1471__;
  wire __1472__;
  wire __1473__;
  wire __1474__;
  wire __1475__;
  wire __1476__;
  wire __1477__;
  wire __1478__;
  wire __1479__;
  wire __1480__;
  wire __1481__;
  wire __1482__;
  wire __1483__;
  wire __1484__;
  wire __1485__;
  wire __1486__;
  wire __1487__;
  wire __1488__;
  wire __1489__;
  wire __1490__;
  wire __1491__;
  wire __1492__;
  wire __1493__;
  wire __1494__;
  wire __1495__;
  wire __1496__;
  wire __1497__;
  wire __1498__;
  wire __1499__;
  wire __1500__;
  wire __1501__;
  wire __1502__;
  wire __1503__;
  wire __1504__;
  wire __1505__;
  wire __1506__;
  wire __1507__;
  wire __1508__;
  wire __1509__;
  wire __1510__;
  wire __1511__;
  wire __1512__;
  wire __1513__;
  wire __1514__;
  wire __1515__;
  wire __1516__;
  wire __1517__;
  wire __1518__;
  wire __1519__;
  wire __1520__;
  wire __1521__;
  wire __1522__;
  wire __1523__;
  wire __1524__;
  wire __1525__;
  wire __1526__;
  wire __1527__;
  wire __1528__;
  wire __1529__;
  wire __1530__;
  wire __1531__;
  wire __1532__;
  wire __1533__;
  wire __1536__;
  wire __1537__;
  wire __1538__;
  wire __1539__;
  wire __1540__;
  wire __1541__;
  wire __1542__;
  wire __1543__;
  wire __1544__;
  wire __1545__;
  wire __1546__;
  wire __1547__;
  wire __1548__;
  wire __1549__;
  wire __1550__;
  wire __1551__;
  wire __1552__;
  wire __1553__;
  wire __1554__;
  wire __1555__;
  wire __1556__;
  wire __1557__;
  wire __1558__;
  wire __1559__;
  wire __1560__;
  wire __1561__;
  wire __1562__;
  wire __1563__;
  wire __1564__;
  wire __1565__;
  wire __1566__;
  wire __1567__;
  wire __1568__;
  wire __1569__;
  wire __1570__;
  wire __1571__;
  wire __1572__;
  wire __1573__;
  wire __1574__;
  wire __1575__;
  wire __1576__;
  wire __1577__;
  wire __1578__;
  wire __1579__;
  wire __1580__;
  wire __1581__;
  wire __1582__;
  wire __1583__;
  wire __1584__;
  wire __1585__;
  wire __1586__;
  wire __1587__;
  wire __1588__;
  wire __1589__;
  wire __1590__;
  wire __1591__;
  wire __1592__;
  wire __1593__;
  wire __1594__;
  wire __1595__;
  wire __1596__;
  wire __1597__;
  wire __1598__;
  wire __1599__;
  wire __1600__;
  wire __1601__;
  wire __1602__;
  wire __1603__;
  wire __1604__;
  wire __1605__;
  wire __1606__;
  wire __1607__;
  wire __1608__;
  wire __1609__;
  wire __1610__;
  wire __1611__;
  wire __1612__;
  wire __1613__;
  wire __1614__;
  wire __1615__;
  wire __1616__;
  wire __1617__;
  wire __1618__;
  wire __1619__;
  wire __1620__;
  wire __1621__;
  wire __1622__;
  wire __1623__;
  wire __1624__;
  wire __1625__;
  wire __1626__;
  wire __1627__;
  wire __1628__;
  wire __1629__;
  wire __1630__;
  wire __1631__;
  wire __1632__;
  wire __1633__;
  wire __1634__;
  wire __1635__;
  wire __1636__;
  wire __1637__;
  wire __1638__;
  wire __1639__;
  wire __1640__;
  wire __1641__;
  wire __1642__;
  wire __1643__;
  wire __1644__;
  wire __1645__;
  wire __1646__;
  wire __1647__;
  wire __1648__;
  wire __1649__;
  wire __1650__;
  wire __1651__;
  wire __1652__;
  wire __1653__;
  wire __1654__;
  wire __1655__;
  wire __1656__;
  wire __1657__;
  wire __1658__;
  wire __1659__;
  wire __1660__;
  wire __1661__;
  wire __1662__;
  wire __1663__;
  wire __1664__;
  wire __1665__;
  wire __1666__;
  wire __1667__;
  wire __1668__;
  wire __1669__;
  wire __1670__;
  wire __1671__;
  wire __1672__;
  wire __1673__;
  wire __1674__;
  wire __1675__;
  wire __1676__;
  wire __1677__;
  wire __1678__;
  wire __1679__;
  wire __1680__;
  wire __1681__;
  wire __1682__;
  wire __1683__;
  wire __1684__;
  wire __1685__;
  wire __1686__;
  wire __1687__;
  wire __1688__;
  wire __1689__;
  wire __1690__;
  wire __1691__;
  wire __1692__;
  wire __1693__;
  wire __1694__;
  wire __1695__;
  wire __1696__;
  wire __1697__;
  wire __1698__;
  wire __1699__;
  wire __1700__;
  wire __1701__;
  wire __1702__;
  wire __1703__;
  wire __1704__;
  wire __1705__;
  wire __1706__;
  wire __1707__;
  wire __1708__;
  wire __1709__;
  wire __1710__;
  wire __1711__;
  wire __1712__;
  wire __1713__;
  wire __1714__;
  wire __1715__;
  wire __1716__;
  wire __1717__;
  wire __1718__;
  wire __1719__;
  wire __1720__;
  wire __1721__;
  wire __1722__;
  wire __1723__;
  wire __1724__;
  wire __1725__;
  wire __1726__;
  wire __1727__;
  wire __1728__;
  wire __1729__;
  wire __1730__;
  wire __1731__;
  wire __1732__;
  wire __1733__;
  wire __1734__;
  wire __1735__;
  wire __1736__;
  wire __1737__;
  wire __1738__;
  wire __1739__;
  wire __1740__;
  wire __1741__;
  wire __1742__;
  wire __1743__;
  wire __1744__;
  wire __1745__;
  wire __1746__;
  wire __1747__;
  wire __1748__;
  wire __1749__;
  wire __1750__;
  wire __1751__;
  wire __1752__;
  wire __1753__;
  wire __1754__;
  wire __1755__;
  wire __1756__;
  wire __1757__;
  wire __1758__;
  wire __1759__;
  wire __1760__;
  wire __1761__;
  wire __1762__;
  wire __1763__;
  wire __1764__;
  wire __1765__;
  wire __1766__;
  wire __1767__;
  wire __1768__;
  wire __1769__;
  wire __1770__;
  wire __1771__;
  wire __1772__;
  wire __1773__;
  wire __1774__;
  wire __1775__;
  wire __1776__;
  wire __1777__;
  wire __1778__;
  wire __1779__;
  wire __1780__;
  wire __1781__;
  wire __1782__;
  wire __1783__;
  wire __1784__;
  wire __1785__;
  wire __1786__;
  wire __1787__;
  wire __1788__;
  wire __1789__;
  wire __1790__;
  wire __1791__;
  wire __1792__;
  wire __1793__;
  wire __1794__;
  wire __1795__;
  wire __1796__;
  wire __1797__;
  wire __1798__;
  wire __1799__;
  wire __1800__;
  wire __1801__;
  wire __1802__;
  wire __1803__;
  wire __1804__;
  wire __1805__;
  wire __1806__;
  wire __1807__;
  wire __1808__;
  wire __1809__;
  wire __1810__;
  wire __1811__;
  wire __1812__;
  wire __1813__;
  wire __1814__;
  wire __1815__;
  wire __1816__;
  wire __1817__;
  wire __1818__;
  wire __1819__;
  wire __1820__;
  wire __1821__;
  wire __1822__;
  wire __1823__;
  wire __1824__;
  wire __1825__;
  wire __1826__;
  wire __1827__;
  wire __1828__;
  wire __1829__;
  wire __1830__;
  wire __1831__;
  wire __1832__;
  wire __1833__;
  wire __1834__;
  wire __1835__;
  wire __1836__;
  wire __1837__;
  wire __1838__;
  wire __1839__;
  wire __1840__;
  wire __1841__;
  wire __1842__;
  wire __1843__;
  wire __1844__;
  wire __1845__;
  wire __1846__;
  wire __1847__;
  wire __1848__;
  wire __1849__;
  wire __1850__;
  wire __1851__;
  wire __1852__;
  wire __1853__;
  wire __1854__;
  wire __1855__;
  wire __1856__;
  wire __1857__;
  wire __1858__;
  wire __1859__;
  wire __1860__;
  wire __1861__;
  wire __1862__;
  wire __1863__;
  wire __1864__;
  wire __1865__;
  wire __1866__;
  wire __1867__;
  wire __1868__;
  wire __1869__;
  wire __1870__;
  wire __1871__;
  wire __1872__;
  wire __1873__;
  wire __1874__;
  wire __1875__;
  wire __1876__;
  wire __1877__;
  wire __1878__;
  wire __1879__;
  wire __1880__;
  wire __1881__;
  wire __1882__;
  wire __1883__;
  wire __1884__;
  wire __1885__;
  wire __1886__;
  wire __1887__;
  wire __1888__;
  wire __1889__;
  wire __1890__;
  wire __1891__;
  wire __1892__;
  wire __1893__;
  wire __1894__;
  wire __1895__;
  wire __1896__;
  wire __1897__;
  wire __1898__;
  wire __1899__;
  wire __1900__;
  wire __1901__;
  wire __1902__;
  wire __1903__;
  wire __1904__;
  wire __1905__;
  wire __1906__;
  wire __1907__;
  wire __1908__;
  wire __1909__;
  wire __1910__;
  wire __1911__;
  wire __1912__;
  wire __1913__;
  wire __1914__;
  wire __1915__;
  wire __1916__;
  wire __1917__;
  wire __1918__;
  wire __1919__;
  wire __1920__;
  wire __1921__;
  wire __1922__;
  wire __1923__;
  wire __1924__;
  wire __1925__;
  wire __1926__;
  wire __1927__;
  wire __1928__;
  wire __1929__;
  wire __1930__;
  wire __1931__;
  wire __1932__;
  wire __1933__;
  wire __1934__;
  wire __1935__;
  wire __1936__;
  wire __1937__;
  wire __1938__;
  wire __1939__;
  wire __1940__;
  wire __1941__;
  wire __1942__;
  wire __1943__;
  wire __1944__;
  wire __1945__;
  wire __1946__;
  wire __1947__;
  wire __1948__;
  wire __1949__;
  wire __1950__;
  wire __1951__;
  wire __1952__;
  wire __1953__;
  wire __1954__;
  wire __1955__;
  wire __1956__;
  wire __1957__;
  wire __1958__;
  wire __1959__;
  wire __1960__;
  wire __1961__;
  wire __1962__;
  wire __1963__;
  wire __1964__;
  wire __1965__;
  wire __1966__;
  wire __1967__;
  wire __1968__;
  wire __1969__;
  wire __1970__;
  wire __1971__;
  wire __1972__;
  wire __1973__;
  wire __1974__;
  wire __1975__;
  wire __1976__;
  wire __1977__;
  wire __1978__;
  wire __1979__;
  wire __1980__;
  wire __1981__;
  wire __1982__;
  wire __1983__;
  wire __1984__;
  wire __1985__;
  wire __1986__;
  wire __1987__;
  wire __1988__;
  wire __1989__;
  wire __1990__;
  wire __1991__;
  wire __1992__;
  wire __1993__;
  wire __1994__;
  wire __1995__;
  wire __1996__;
  wire __1997__;
  wire __1998__;
  wire __1999__;
  wire __2000__;
  wire __2001__;
  wire __2002__;
  wire __2003__;
  wire __2004__;
  wire __2005__;
  wire __2006__;
  wire __2007__;
  wire __2008__;
  wire __2009__;
  wire __2010__;
  wire __2011__;
  wire __2012__;
  wire __2013__;
  wire __2014__;
  wire __2015__;
  wire __2016__;
  wire __2017__;
  wire __2018__;
  wire __2019__;
  wire __2020__;
  wire __2021__;
  wire __2022__;
  wire __2023__;
  wire __2024__;
  wire __2025__;
  wire __2026__;
  wire __2027__;
  wire __2028__;
  wire __2029__;
  wire __2030__;
  wire __2031__;
  wire __2032__;
  wire __2033__;
  wire __2034__;
  wire __2035__;
  wire __2036__;
  wire __2037__;
  wire __2038__;
  wire __2039__;
  wire __2040__;
  wire __2041__;
  wire __2042__;
  wire __2043__;
  wire __2044__;
  wire __2045__;
  wire __2046__;
  wire __2047__;
  wire __2048__;
  wire __2049__;
  wire __2050__;
  wire __2051__;
  wire __2052__;
  wire __2053__;
  wire __2054__;
  wire __2055__;
  wire __2056__;
  wire __2057__;
  wire __2058__;
  wire __2059__;
  wire __2060__;
  wire __2061__;
  wire __2062__;
  wire __2063__;
  wire __2064__;
  wire __2065__;
  wire __2066__;
  wire __2067__;
  wire __2068__;
  wire __2069__;
  wire __2070__;
  wire __2071__;
  wire __2072__;
  wire __2073__;
  wire __2074__;
  wire __2075__;
  wire __2076__;
  wire __2077__;
  wire __2078__;
  wire __2079__;
  wire __2080__;
  wire __2081__;
  wire __2082__;
  wire __2083__;
  wire __2084__;
  wire __2085__;
  wire __2086__;
  wire __2087__;
  wire __2088__;
  wire __2089__;
  wire __2090__;
  wire __2091__;
  wire __2092__;
  wire __2093__;
  wire __2094__;
  wire __2095__;
  wire __2096__;
  wire __2097__;
  wire __2098__;
  wire __2099__;
  wire __2100__;
  wire __2101__;
  wire __2102__;
  wire __2103__;
  wire __2104__;
  wire __2105__;
  wire __2106__;
  wire __2107__;
  wire __2108__;
  wire __2109__;
  wire __2110__;
  wire __2111__;
  wire __2112__;
  wire __2113__;
  wire __2114__;
  wire __2115__;
  wire __2116__;
  wire __2117__;
  wire __2118__;
  wire __2119__;
  wire __2120__;
  wire __2121__;
  wire __2122__;
  wire __2123__;
  wire __2124__;
  wire __2125__;
  wire __2126__;
  wire __2127__;
  wire __2128__;
  wire __2129__;
  wire __2130__;
  wire __2131__;
  wire __2132__;
  wire __2133__;
  wire __2134__;
  wire __2135__;
  wire __2136__;
  wire __2137__;
  wire __2138__;
  wire __2139__;
  wire __2140__;
  wire __2141__;
  wire __2142__;
  wire __2143__;
  wire __2144__;
  wire __2145__;
  wire __2146__;
  wire __2147__;
  wire __2148__;
  wire __2149__;
  wire __2150__;
  wire __2151__;
  wire __2152__;
  wire __2153__;
  wire __2154__;
  wire __2155__;
  wire __2156__;
  wire __2157__;
  wire __2158__;
  wire __2159__;
  wire __2160__;
  wire __2161__;
  wire __2162__;
  wire __2163__;
  wire __2164__;
  wire __2165__;
  wire __2166__;
  wire __2167__;
  wire __2168__;
  wire __2169__;
  wire __2170__;
  wire __2171__;
  wire __2172__;
  wire __2173__;
  wire __2174__;
  wire __2175__;
  wire __2176__;
  wire __2177__;
  wire __2178__;
  wire __2179__;
  wire __2180__;
  wire __2181__;
  wire __2182__;
  wire __2183__;
  wire __2184__;
  wire __2185__;
  wire __2186__;
  wire __2187__;
  wire __2188__;
  wire __2189__;
  wire __2190__;
  wire __2191__;
  wire __2192__;
  wire __2193__;
  wire __2194__;
  wire __2195__;
  wire __2196__;
  wire __2197__;
  wire __2198__;
  wire __2199__;
  wire __2200__;
  wire __2201__;
  wire __2202__;
  wire __2203__;
  wire __2204__;
  wire __2205__;
  wire __2206__;
  wire __2207__;
  wire __2208__;
  wire __2209__;
  wire __2210__;
  wire __2211__;
  wire __2212__;
  wire __2213__;
  wire __2214__;
  wire __2215__;
  wire __2216__;
  wire __2217__;
  wire __2218__;
  wire __2219__;
  wire __2220__;
  wire __2221__;
  wire __2222__;
  wire __2223__;
  wire __2224__;
  wire __2225__;
  wire __2226__;
  wire __2227__;
  wire __2228__;
  wire __2229__;
  wire __2230__;
  wire __2231__;
  wire __2232__;
  wire __2233__;
  wire __2234__;
  wire __2235__;
  wire __2236__;
  wire __2237__;
  wire __2238__;
  wire __2239__;
  wire __2240__;
  wire __2241__;
  wire __2242__;
  wire __2243__;
  wire __2244__;
  wire __2245__;
  wire __2246__;
  wire __2247__;
  wire __2248__;
  wire __2249__;
  wire __2250__;
  wire __2251__;
  wire __2252__;
  wire __2253__;
  wire __2254__;
  wire __2255__;
  wire __2256__;
  wire __2257__;
  wire __2258__;
  wire __2259__;
  wire __2260__;
  wire __2261__;
  wire __2262__;
  wire __2263__;
  wire __2264__;
  wire __2265__;
  wire __2266__;
  wire __2267__;
  wire __2268__;
  wire __2269__;
  wire __2270__;
  wire __2271__;
  wire __2272__;
  wire __2273__;
  wire __2274__;
  wire __2275__;
  wire __2276__;
  wire __2277__;
  wire __2278__;
  wire __2279__;
  wire __2280__;
  wire __2281__;
  wire __2282__;
  wire __2283__;
  wire __2284__;
  wire __2285__;
  wire __2286__;
  wire __2287__;
  wire __2288__;
  wire __2289__;
  wire __2290__;
  wire __2291__;
  wire __2292__;
  wire __2293__;
  wire __2294__;
  wire __2295__;
  wire __2296__;
  wire __2297__;
  wire __2298__;
  wire __2299__;
  wire __2300__;
  wire __2301__;
  wire __2302__;
  wire __2303__;
  wire __2304__;
  wire __2305__;
  wire __2306__;
  wire __2307__;
  wire __2308__;
  wire __2309__;
  wire __2310__;
  wire __2311__;
  wire __2312__;
  wire __2313__;
  wire __2314__;
  wire __2315__;
  wire __2316__;
  wire __2317__;
  wire __2318__;
  wire __2319__;
  wire __2320__;
  wire __2321__;
  wire __2322__;
  wire __2323__;
  wire __2324__;
  wire __2325__;
  wire __2326__;
  wire __2327__;
  wire __2328__;
  wire __2329__;
  wire __2330__;
  wire __2331__;
  wire __2332__;
  wire __2333__;
  wire __2334__;
  wire __2335__;
  wire __2336__;
  wire __2337__;
  wire __2338__;
  wire __2339__;
  wire __2340__;
  wire __2341__;
  wire __2342__;
  wire __2343__;
  wire __2344__;
  wire __2345__;
  wire __2346__;
  wire __2347__;
  wire __2348__;
  wire __2349__;
  wire __2350__;
  wire __2351__;
  wire __2352__;
  wire __2353__;
  wire __2354__;
  wire __2355__;
  wire __2356__;
  wire __2357__;
  wire __2358__;
  wire __2359__;
  wire __2360__;
  wire __2361__;
  wire __2362__;
  wire __2363__;
  wire __2364__;
  wire __2365__;
  wire __2366__;
  wire __2367__;
  wire __2368__;
  wire __2369__;
  wire __2370__;
  wire __2371__;
  wire __2372__;
  wire __2373__;
  wire __2374__;
  wire __2375__;
  wire __2376__;
  wire __2377__;
  wire __2378__;
  wire __2379__;
  wire __2380__;
  wire __2381__;
  wire __2382__;
  wire __2383__;
  wire __2384__;
  wire __2385__;
  wire __2386__;
  wire __2387__;
  wire __2388__;
  wire __2389__;
  wire __2390__;
  wire __2391__;
  wire __2392__;
  wire __2393__;
  wire __2394__;
  wire __2395__;
  wire __2396__;
  wire __2397__;
  wire __2398__;
  wire __2399__;
  wire __2400__;
  wire __2401__;
  wire __2402__;
  wire __2403__;
  wire __2404__;
  wire __2405__;
  wire __2406__;
  wire __2407__;
  wire __2408__;
  wire __2409__;
  wire __2410__;
  wire __2411__;
  wire __2412__;
  wire __2413__;
  wire __2414__;
  wire __2415__;
  wire __2416__;
  wire __2417__;
  wire __2418__;
  wire __2419__;
  wire __2420__;
  wire __2421__;
  wire __2422__;
  wire __2423__;
  wire __2424__;
  wire __2425__;
  wire __2426__;
  wire __2427__;
  wire __2428__;
  wire __2429__;
  wire __2430__;
  wire __2431__;
  wire __2432__;
  wire __2433__;
  wire __2434__;
  wire __2435__;
  wire __2436__;
  wire __2437__;
  wire __2438__;
  wire __2439__;
  wire __2440__;
  wire __2441__;
  wire __2442__;
  wire __2443__;
  wire __2444__;
  wire __2445__;
  wire __2446__;
  wire __2447__;
  wire __2448__;
  wire __2449__;
  wire __2450__;
  wire __2451__;
  wire __2452__;
  wire __2453__;
  wire __2454__;
  wire __2455__;
  wire __2456__;
  wire __2457__;
  wire __2458__;
  wire __2459__;
  wire __2460__;
  wire __2461__;
  wire __2462__;
  wire __2463__;
  wire __2464__;
  wire __2465__;
  wire __2466__;
  wire __2467__;
  wire __2468__;
  wire __2469__;
  wire __2470__;
  wire __2471__;
  wire __2472__;
  wire __2473__;
  wire __2474__;
  wire __2475__;
  wire __2476__;
  wire __2477__;
  wire __2478__;
  wire __2479__;
  wire __2480__;
  wire __2481__;
  wire __2482__;
  wire __2483__;
  wire __2484__;
  wire __2485__;
  wire __2486__;
  wire __2487__;
  wire __2488__;
  wire __2489__;
  wire __2490__;
  wire __2491__;
  wire __2492__;
  wire __2493__;
  wire __2494__;
  wire __2495__;
  wire __2496__;
  wire __2497__;
  wire __2498__;
  wire __2499__;
  wire __2500__;
  wire __2501__;
  wire __2502__;
  wire __2503__;
  wire __2504__;
  wire __2505__;
  wire __2506__;
  wire __2507__;
  wire __2508__;
  wire __2509__;
  wire __2510__;
  wire __2511__;
  wire __2512__;
  wire __2513__;
  wire __2514__;
  wire __2515__;
  wire __2516__;
  wire __2517__;
  wire __2518__;
  wire __2519__;
  wire __2520__;
  wire __2521__;
  wire __2522__;
  wire __2523__;
  wire __2524__;
  wire __2525__;
  wire __2526__;
  wire __2527__;
  wire __2528__;
  wire __2529__;
  wire __2530__;
  wire __2531__;
  wire __2532__;
  wire __2533__;
  wire __2534__;
  wire __2535__;
  wire __2536__;
  wire __2537__;
  wire __2538__;
  wire __2539__;
  wire __2540__;
  wire __2541__;
  wire __2542__;
  wire __2543__;
  wire __2544__;
  wire __2545__;
  wire __2546__;
  wire __2547__;
  wire __2548__;
  wire __2549__;
  wire __2550__;
  wire __2551__;
  wire __2552__;
  wire __2553__;
  wire __2554__;
  wire __2555__;
  wire __2556__;
  wire __2557__;
  wire __2558__;
  wire __2559__;
  wire __2560__;
  wire __2561__;
  wire __2562__;
  wire __2563__;
  wire __2564__;
  wire __2565__;
  wire __2566__;
  wire __2567__;
  wire __2568__;
  wire __2569__;
  wire __2570__;
  wire __2571__;
  wire __2572__;
  wire __2573__;
  wire __2574__;
  wire __2575__;
  wire __2576__;
  wire __2577__;
  wire __2578__;
  wire __2579__;
  wire __2580__;
  wire __2581__;
  wire __2582__;
  wire __2583__;
  wire __2584__;
  wire __2585__;
  wire __2586__;
  wire __2587__;
  wire __2588__;
  wire __2589__;
  wire __2590__;
  wire __2591__;
  wire __2592__;
  wire __2593__;
  wire __2594__;
  wire __2595__;
  wire __2596__;
  wire __2597__;
  wire __2598__;
  wire __2599__;
  wire __2600__;
  wire __2601__;
  wire __2602__;
  wire __2603__;
  wire __2604__;
  wire __2605__;
  wire __2606__;
  wire __2607__;
  wire __2608__;
  wire __2609__;
  wire __2610__;
  wire __2611__;
  wire __2612__;
  wire __2613__;
  wire __2614__;
  wire __2615__;
  wire __2616__;
  wire __2617__;
  wire __2618__;
  wire __2619__;
  wire __2620__;
  wire __2621__;
  wire __2622__;
  wire __2623__;
  wire __2624__;
  wire __2625__;
  wire __2626__;
  wire __2627__;
  wire __2628__;
  wire __2629__;
  wire __2630__;
  wire __2631__;
  wire __2632__;
  wire __2633__;
  wire __2634__;
  wire __2635__;
  wire __2636__;
  wire __2637__;
  wire __2638__;
  wire __2639__;
  wire __2640__;
  wire __2641__;
  wire __2642__;
  wire __2643__;
  wire __2644__;
  wire __2645__;
  wire __2646__;
  wire __2647__;
  wire __2648__;
  wire __2649__;
  wire __2650__;
  wire __2651__;
  wire __2652__;
  wire __2653__;
  wire __2654__;
  wire __2655__;
  wire __2656__;
  wire __2657__;
  wire __2658__;
  wire __2659__;
  wire __2660__;
  wire __2661__;
  wire __2662__;
  wire __2663__;
  wire __2664__;
  wire __2665__;
  wire __2666__;
  wire __2667__;
  wire __2668__;
  wire __2669__;
  wire __2670__;
  wire __2671__;
  wire __2672__;
  wire __2673__;
  wire __2674__;
  wire __2675__;
  wire __2676__;
  wire __2677__;
  wire __2678__;
  wire __2679__;
  wire __2680__;
  wire __2681__;
  wire __2682__;
  wire __2683__;
  wire __2684__;
  wire __2685__;
  wire __2686__;
  wire __2687__;
  wire __2688__;
  wire __2689__;
  wire __2690__;
  wire __2691__;
  wire __2692__;
  wire __2693__;
  wire __2694__;
  wire __2695__;
  wire __2696__;
  wire __2697__;
  wire __2698__;
  wire __2699__;
  wire __2700__;
  wire __2701__;
  wire __2702__;
  wire __2703__;
  wire __2704__;
  wire __2705__;
  wire __2706__;
  wire __2707__;
  wire __2708__;
  wire __2709__;
  wire __2710__;
  wire __2711__;
  wire __2712__;
  wire __2713__;
  wire __2714__;
  wire __2715__;
  wire __2716__;
  wire __2717__;
  wire __2718__;
  wire __2719__;
  wire __2720__;
  wire __2721__;
  wire __2722__;
  wire __2723__;
  wire __2724__;
  wire __2725__;
  wire __2726__;
  wire __2727__;
  wire __2728__;
  wire __2729__;
  wire __2730__;
  wire __2731__;
  wire __2732__;
  wire __2733__;
  wire __2734__;
  wire __2735__;
  wire __2736__;
  wire __2737__;
  wire __2738__;
  wire __2739__;
  wire __2740__;
  wire __2741__;
  wire __2742__;
  wire __2743__;
  wire __2744__;
  wire __2745__;
  wire __2746__;
  wire __2747__;
  wire __2748__;
  wire __2749__;
  wire __2750__;
  wire __2751__;
  wire __2752__;
  wire __2753__;
  wire __2754__;
  wire __2755__;
  wire __2756__;
  wire __2757__;
  wire __2758__;
  wire __2759__;
  wire __2760__;
  wire __2761__;
  wire __2762__;
  wire __2763__;
  wire __2764__;
  wire __2765__;
  wire __2766__;
  wire __2767__;
  wire __2768__;
  wire __2769__;
  wire __2770__;
  wire __2771__;
  wire __2772__;
  wire __2773__;
  wire __2774__;
  wire __2775__;
  wire __2776__;
  wire __2777__;
  wire __2778__;
  wire __2779__;
  wire __2780__;
  wire __2781__;
  wire __2782__;
  wire __2783__;
  wire __2784__;
  wire __2785__;
  wire __2786__;
  wire __2787__;
  wire __2788__;
  wire __2789__;
  wire __2790__;
  wire __2791__;
  wire __2792__;
  wire __2793__;
  wire __2794__;
  wire __2795__;
  wire __2796__;
  wire __2797__;
  wire __2798__;
  wire __2799__;
  wire __2800__;
  wire __2801__;
  wire __2802__;
  wire __2803__;
  wire __2804__;
  wire __2805__;
  wire __2806__;
  wire __2807__;
  wire __2808__;
  wire __2809__;
  wire __2810__;
  wire __2811__;
  wire __2812__;
  wire __2813__;
  wire __2814__;
  wire __2815__;
  wire __2816__;
  wire __2817__;
  wire __2818__;
  wire __2819__;
  wire __2820__;
  wire __2821__;
  wire __2822__;
  wire __2823__;
  wire __2824__;
  wire __2825__;
  wire __2826__;
  wire __2827__;
  wire __2828__;
  wire __2829__;
  wire __2830__;
  wire __2831__;
  wire __2832__;
  wire __2833__;
  wire __2834__;
  wire __2835__;
  wire __2836__;
  wire __2837__;
  wire __2838__;
  wire __2839__;
  wire __2840__;
  wire __2841__;
  wire __2842__;
  wire __2843__;
  wire __2844__;
  wire __2845__;
  wire __2846__;
  wire __2847__;
  wire __2848__;
  wire __2849__;
  wire __2850__;
  wire __2851__;
  wire __2852__;
  wire __2853__;
  wire __2854__;
  wire __2855__;
  wire __2856__;
  wire __2857__;
  wire __2858__;
  wire __2859__;
  wire __2860__;
  wire __2861__;
  wire __2862__;
  wire __2863__;
  wire __2864__;
  wire __2865__;
  wire __2866__;
  wire __2867__;
  wire __2868__;
  wire __2869__;
  wire __2870__;
  wire __2871__;
  wire __2872__;
  wire __2873__;
  wire __2874__;
  wire __2875__;
  wire __2876__;
  wire __2877__;
  wire __2878__;
  wire __2879__;
  wire __2880__;
  wire __2881__;
  wire __2882__;
  wire __2883__;
  wire __2884__;
  wire __2885__;
  wire __2886__;
  wire __2887__;
  wire __2888__;
  wire __2889__;
  wire __2890__;
  wire __2891__;
  wire __2892__;
  wire __2893__;
  wire __2894__;
  wire __2895__;
  wire __2896__;
  wire __2897__;
  wire __2898__;
  wire __2899__;
  wire __2900__;
  wire __2901__;
  wire __2902__;
  wire __2903__;
  wire __2904__;
  wire __2905__;
  wire __2906__;
  wire __2907__;
  wire __2908__;
  wire __2909__;
  wire __2910__;
  wire __2911__;
  wire __2912__;
  wire __2913__;
  wire __2914__;
  wire __2915__;
  wire __2916__;
  wire __2917__;
  wire __2918__;
  wire __2919__;
  wire __2920__;
  wire __2921__;
  wire __2922__;
  wire __2923__;
  wire __2924__;
  wire __2925__;
  wire __2926__;
  wire __2927__;
  wire __2928__;
  wire __2929__;
  wire __2930__;
  wire __2931__;
  wire __2932__;
  wire __2933__;
  wire __2934__;
  wire __2935__;
  wire __2936__;
  wire __2937__;
  wire __2938__;
  wire __2939__;
  wire __2940__;
  wire __2941__;
  wire __2942__;
  wire __2943__;
  wire __2944__;
  wire __2945__;
  wire __2946__;
  wire __2947__;
  wire __2948__;
  wire __2949__;
  wire __2950__;
  wire __2951__;
  wire __2952__;
  wire __2953__;
  wire __2954__;
  wire __2955__;
  wire __2956__;
  wire __2957__;
  wire __2958__;
  wire __2959__;
  wire __2960__;
  wire __2961__;
  wire __2962__;
  wire __2963__;
  wire __2964__;
  wire __2965__;
  wire __2966__;
  wire __2967__;
  wire __2968__;
  wire __2969__;
  wire __2970__;
  wire __2971__;
  wire __2972__;
  wire __2973__;
  wire __2974__;
  wire __2975__;
  wire __2976__;
  wire __2977__;
  wire __2978__;
  wire __2979__;
  wire __2980__;
  wire __2981__;
  wire __2982__;
  wire __2983__;
  wire __2984__;
  wire __2985__;
  wire __2986__;
  wire __2987__;
  wire __2988__;
  wire __2989__;
  wire __2990__;
  wire __2991__;
  wire __2992__;
  wire __2993__;
  wire __2994__;
  wire __2995__;
  wire __2996__;
  wire __2997__;
  wire __2998__;
  wire __2999__;
  wire __3000__;
  wire __3001__;
  wire __3002__;
  wire __3003__;
  wire __3004__;
  wire __3005__;
  wire __3006__;
  wire __3007__;
  wire __3008__;
  wire __3009__;
  wire __3010__;
  wire __3011__;
  wire __3012__;
  wire __3013__;
  wire __3014__;
  wire __3015__;
  wire __3016__;
  wire __3017__;
  wire __3018__;
  wire __3019__;
  wire __3020__;
  wire __3021__;
  wire __3022__;
  wire __3023__;
  wire __3024__;
  wire __3025__;
  wire __3026__;
  wire __3027__;
  wire __3028__;
  wire __3029__;
  wire __3030__;
  wire __3031__;
  wire __3032__;
  wire __3033__;
  wire __3034__;
  wire __3035__;
  wire __3036__;
  wire __3037__;
  wire __3038__;
  wire __3039__;
  wire __3040__;
  wire __3041__;
  wire __3042__;
  wire __3043__;
  wire __3044__;
  wire __3045__;
  wire __3046__;
  wire __3047__;
  wire __3048__;
  wire __3049__;
  wire __3050__;
  wire __3051__;
  wire __3052__;
  wire __3053__;
  wire __3054__;
  wire __3055__;
  wire __3056__;
  wire __3057__;
  wire __3058__;
  wire __3059__;
  wire __3060__;
  wire __3061__;
  wire __3062__;
  wire __3063__;
  wire __3064__;
  wire __3065__;
  wire __3066__;
  wire __3067__;
  wire __3068__;
  wire __3069__;
  wire __3070__;
  wire __3071__;
  wire __3072__;
  wire __3073__;
  wire __3074__;
  wire __3075__;
  wire __3076__;
  wire __3077__;
  wire __3078__;
  wire __3079__;
  wire __3080__;
  wire __3081__;
  wire __3082__;
  wire __3083__;
  wire __3084__;
  wire __3085__;
  wire __3086__;
  wire __3087__;
  wire __3088__;
  wire __3089__;
  wire __3090__;
  wire __3091__;
  wire __3092__;
  wire __3093__;
  wire __3094__;
  wire __3095__;
  wire __3096__;
  wire __3097__;
  wire __3098__;
  wire __3099__;
  wire __3100__;
  wire __3101__;
  wire __3102__;
  wire __3103__;
  wire __3104__;
  wire __3105__;
  wire __3106__;
  wire __3107__;
  wire __3108__;
  wire __3109__;
  wire __3110__;
  wire __3111__;
  wire __3112__;
  wire __3113__;
  wire __3114__;
  wire __3115__;
  wire __3116__;
  wire __3117__;
  wire __3118__;
  wire __3119__;
  wire __3120__;
  wire __3121__;
  wire __3122__;
  wire __3123__;
  wire __3124__;
  wire __3125__;
  wire __3126__;
  wire __3127__;
  wire __3128__;
  wire __3129__;
  wire __3130__;
  wire __3131__;
  wire __3132__;
  wire __3133__;
  wire __3134__;
  wire __3135__;
  wire __3136__;
  wire __3137__;
  wire __3138__;
  wire __3139__;
  wire __3140__;
  wire __3141__;
  wire __3142__;
  wire __3143__;
  wire __3144__;
  wire __3145__;
  wire __3146__;
  wire __3147__;
  wire __3148__;
  wire __3149__;
  wire __3150__;
  wire __3151__;
  wire __3152__;
  wire __3153__;
  wire __3154__;
  wire __3155__;
  wire __3156__;
  wire __3157__;
  wire __3158__;
  wire __3159__;
  wire __3160__;
  wire __3161__;
  wire __3162__;
  wire __3163__;
  wire __3164__;
  wire __3165__;
  wire __3166__;
  wire __3167__;
  wire __3168__;
  wire __3169__;
  wire __3170__;
  wire __3171__;
  wire __3172__;
  wire __3173__;
  wire __3174__;
  wire __3175__;
  wire __3176__;
  wire __3177__;
  wire __3178__;
  wire __3179__;
  wire __3180__;
  wire __3181__;
  wire __3182__;
  wire __3183__;
  wire __3184__;
  wire __3185__;
  wire __3186__;
  wire __3187__;
  wire __3188__;
  wire __3189__;
  wire __3190__;
  wire __3191__;
  wire __3192__;
  wire __3193__;
  wire __3194__;
  wire __3195__;
  wire __3196__;
  wire __3197__;
  wire __3198__;
  wire __3199__;
  wire __3200__;
  wire __3201__;
  wire __3202__;
  wire __3203__;
  wire __3204__;
  wire __3205__;
  wire __3206__;
  wire __3207__;
  wire __3208__;
  wire __3209__;
  wire __3210__;
  wire __3211__;
  wire __3212__;
  wire __3213__;
  wire __3214__;
  wire __3215__;
  wire __3216__;
  wire __3217__;
  wire __3218__;
  wire __3219__;
  wire __3220__;
  wire __3221__;
  wire __3222__;
  wire __3223__;
  wire __3224__;
  wire __3225__;
  wire __3226__;
  wire __3227__;
  wire __3228__;
  wire __3229__;
  wire __3230__;
  wire __3231__;
  wire __3232__;
  wire __3233__;
  wire __3234__;
  wire __3235__;
  wire __3236__;
  wire __3237__;
  wire __3238__;
  wire __3239__;
  wire __3240__;
  wire __3241__;
  wire __3242__;
  wire __3243__;
  wire __3244__;
  wire __3245__;
  wire __3246__;
  wire __3247__;
  wire __3248__;
  wire __3249__;
  wire __3250__;
  wire __3251__;
  wire __3252__;
  wire __3253__;
  wire __3254__;
  wire __3255__;
  wire __3256__;
  wire __3257__;
  wire __3258__;
  wire __3259__;
  wire __3260__;
  wire __3261__;
  wire __3262__;
  wire __3263__;
  wire __3264__;
  wire __3265__;
  wire __3266__;
  wire __3267__;
  wire __3268__;
  wire __3269__;
  wire __3270__;
  wire __3271__;
  wire __3272__;
  wire __3273__;
  wire __3274__;
  wire __3275__;
  wire __3276__;
  wire __3277__;
  wire __3278__;
  wire __3279__;
  wire __3280__;
  wire __3281__;
  wire __3282__;
  wire __3283__;
  wire __3284__;
  wire __3285__;
  wire __3286__;
  wire __3287__;
  wire __3288__;
  wire __3289__;
  wire __3290__;
  wire __3291__;
  wire __3292__;
  wire __3293__;
  wire __3294__;
  wire __3295__;
  wire __3296__;
  wire __3297__;
  wire __3298__;
  wire __3299__;
  wire __3300__;
  wire __3301__;
  wire __3302__;
  wire __3303__;
  wire __3304__;
  wire __3305__;
  wire __3306__;
  wire __3307__;
  wire __3308__;
  wire __3309__;
  wire __3310__;
  wire __3311__;
  wire __3312__;
  wire __3313__;
  wire __3314__;
  wire __3315__;
  wire __3316__;
  wire __3317__;
  wire __3318__;
  wire __3319__;
  wire __3320__;
  wire __3321__;
  wire __3322__;
  wire __3323__;
  wire __3324__;
  wire __3325__;
  wire __3326__;
  wire __3327__;
  wire __3328__;
  wire __3329__;
  wire __3330__;
  wire __3331__;
  wire __3332__;
  wire __3333__;
  wire __3334__;
  wire __3335__;
  wire __3336__;
  wire __3337__;
  wire __3338__;
  wire __3339__;
  wire __3340__;
  wire __3341__;
  wire __3342__;
  wire __3343__;
  wire __3344__;
  wire __3345__;
  wire __3346__;
  wire __3347__;
  wire __3348__;
  wire __3349__;
  wire __3350__;
  wire __3351__;
  wire __3352__;
  wire __3353__;
  wire __3354__;
  wire __3355__;
  wire __3356__;
  wire __3357__;
  wire __3358__;
  wire __3359__;
  wire __3360__;
  wire __3361__;
  wire __3362__;
  wire __3363__;
  wire __3364__;
  wire __3365__;
  wire __3366__;
  wire __3367__;
  wire __3368__;
  wire __3369__;
  wire __3370__;
  wire __3371__;
  wire __3372__;
  wire __3373__;
  wire __3374__;
  wire __3375__;
  wire __3376__;
  wire __3377__;
  wire __3378__;
  wire __3379__;
  wire __3380__;
  wire __3381__;
  wire __3382__;
  wire __3383__;
  wire __3384__;
  wire __3385__;
  wire __3386__;
  wire __3387__;
  wire __3388__;
  wire __3389__;
  wire __3390__;
  wire __3391__;
  wire __3392__;
  wire __3393__;
  wire __3394__;
  wire __3395__;
  wire __3396__;
  wire __3397__;
  wire __3398__;
  wire __3399__;
  wire __3400__;
  wire __3401__;
  wire __3402__;
  wire __3403__;
  wire __3404__;
  wire __3405__;
  wire __3406__;
  wire __3407__;
  wire __3408__;
  wire __3409__;
  wire __3410__;
  wire __3411__;
  wire __3412__;
  wire __3413__;
  wire __3414__;
  wire __3415__;
  wire __3416__;
  wire __3417__;
  wire __3418__;
  wire __3419__;
  wire __3420__;
  wire __3421__;
  wire __3422__;
  wire __3423__;
  wire __3424__;
  wire __3425__;
  wire __3426__;
  wire __3427__;
  wire __3428__;
  wire __3429__;
  wire __3430__;
  wire __3431__;
  wire __3432__;
  wire __3433__;
  wire __3434__;
  wire __3435__;
  wire __3436__;
  wire __3437__;
  wire __3438__;
  wire __3439__;
  wire __3440__;
  wire __3441__;
  wire __3442__;
  wire __3443__;
  wire __3444__;
  wire __3445__;
  wire __3446__;
  wire __3447__;
  wire __3448__;
  wire __3449__;
  wire __3450__;
  wire __3451__;
  wire __3452__;
  wire __3453__;
  wire __3454__;
  wire __3455__;
  wire __3456__;
  wire __3457__;
  wire __3458__;
  wire __3459__;
  wire __3460__;
  wire __3461__;
  wire __3462__;
  wire __3463__;
  wire __3464__;
  wire __3465__;
  wire __3466__;
  wire __3467__;
  wire __3468__;
  wire __3469__;
  wire __3470__;
  wire __3471__;
  wire __3472__;
  wire __3473__;
  wire __3474__;
  wire __3475__;
  wire __3476__;
  wire __3477__;
  wire __3478__;
  wire __3479__;
  wire __3480__;
  wire __3481__;
  wire __3482__;
  wire __3483__;
  wire __3484__;
  wire __3485__;
  wire __3486__;
  wire __3487__;
  wire __3488__;
  wire __3489__;
  wire __3490__;
  wire __3491__;
  wire __3492__;
  wire __3493__;
  wire __3494__;
  wire __3495__;
  wire __3496__;
  wire __3497__;
  wire __3498__;
  wire __3499__;
  wire __3500__;
  wire __3501__;
  wire __3502__;
  wire __3503__;
  wire __3504__;
  wire __3505__;
  wire __3506__;
  wire __3507__;
  wire __3508__;
  wire __3509__;
  wire __3510__;
  wire __3511__;
  wire __3512__;
  wire __3513__;
  wire __3514__;
  wire __3515__;
  wire __3516__;
  wire __3517__;
  wire __3518__;
  wire __3519__;
  wire __3520__;
  wire __3521__;
  wire __3522__;
  wire __3523__;
  wire __3524__;
  wire __3525__;
  wire __3526__;
  wire __3527__;
  wire __3528__;
  wire __3529__;
  wire __3530__;
  wire __3531__;
  wire __3532__;
  wire __3533__;
  wire __3534__;
  wire __3535__;
  wire __3536__;
  wire __3537__;
  wire __3538__;
  wire __3539__;
  wire __3540__;
  wire __3541__;
  wire __3542__;
  wire __3543__;
  wire __3544__;
  wire __3545__;
  wire __3546__;
  wire __3547__;
  wire __3548__;
  wire __3549__;
  wire __3550__;
  wire __3551__;
  wire __3552__;
  wire __3553__;
  wire __3554__;
  wire __3555__;
  wire __3556__;
  wire __3557__;
  wire __3558__;
  wire __3559__;
  wire __3560__;
  wire __3561__;
  wire __3562__;
  wire __3563__;
  wire __3564__;
  wire __3565__;
  wire __3566__;
  wire __3567__;
  wire __3568__;
  wire __3569__;
  wire __3570__;
  wire __3571__;
  wire __3572__;
  wire __3573__;
  wire __3574__;
  wire __3575__;
  wire __3576__;
  wire __3577__;
  wire __3578__;
  wire __3579__;
  wire __3580__;
  wire __3581__;
  wire __3582__;
  wire __3583__;
  wire __3584__;
  wire __3585__;
  wire __3586__;
  wire __3587__;
  wire __3588__;
  wire __3589__;
  wire __3590__;
  wire __3591__;
  wire __3592__;
  wire __3593__;
  wire __3594__;
  wire __3595__;
  wire __3596__;
  wire __3597__;
  wire __3598__;
  wire __3599__;
  wire __3600__;
  wire __3601__;
  wire __3602__;
  wire __3603__;
  wire __3604__;
  wire __3605__;
  wire __3606__;
  wire __3607__;
  wire __3608__;
  wire __3609__;
  wire __3610__;
  wire __3611__;
  wire __3612__;
  wire __3613__;
  wire __3614__;
  wire __3615__;
  wire __3616__;
  wire __3617__;
  wire __3618__;
  wire __3619__;
  wire __3620__;
  wire __3621__;
  wire __3622__;
  wire __3623__;
  wire __3624__;
  wire __3625__;
  wire __3626__;
  wire __3627__;
  wire __3628__;
  wire __3629__;
  wire __3630__;
  wire __3631__;
  wire __3632__;
  wire __3633__;
  wire __3634__;
  wire __3635__;
  wire __3636__;
  wire __3637__;
  wire __3638__;
  wire __3639__;
  wire __3640__;
  wire __3641__;
  wire __3642__;
  wire __3643__;
  wire __3644__;
  wire __3645__;
  wire __3646__;
  wire __3647__;
  wire __3648__;
  wire __3649__;
  wire __3650__;
  wire __3651__;
  wire __3652__;
  wire __3653__;
  wire __3654__;
  wire __3655__;
  wire __3656__;
  wire __3657__;
  wire __3658__;
  wire __3659__;
  wire __3660__;
  wire __3661__;
  wire __3662__;
  wire __3663__;
  wire __3664__;
  wire __3665__;
  wire __3666__;
  wire __3667__;
  wire __3668__;
  wire __3669__;
  wire __3670__;
  wire __3671__;
  wire __3672__;
  wire __3673__;
  wire __3674__;
  wire __3675__;
  wire __3676__;
  wire __3677__;
  wire __3678__;
  wire __3679__;
  wire __3680__;
  wire __3681__;
  wire __3682__;
  INV __3683__ (
    .I(__1457__),
    .O(__0__)
  );
  INV __3684__ (
    .I(__1456__),
    .O(__1__)
  );
  INV __3685__ (
    .I(__1455__),
    .O(__2__)
  );
  INV __3686__ (
    .I(__1408__),
    .O(__3__)
  );
  INV __3687__ (
    .I(__1413__),
    .O(__4__)
  );
  INV __3688__ (
    .I(__1454__),
    .O(__5__)
  );
  INV __3689__ (
    .I(__1412__),
    .O(__6__)
  );
  INV __3690__ (
    .I(__1453__),
    .O(__7__)
  );
  INV __3691__ (
    .I(__1409__),
    .O(__8__)
  );
  INV __3692__ (
    .I(__1414__),
    .O(__9__)
  );
  INV __3693__ (
    .I(__1460__),
    .O(__10__)
  );
  INV __3694__ (
    .I(__1410__),
    .O(__11__)
  );
  INV __3695__ (
    .I(__1459__),
    .O(__12__)
  );
  INV __3696__ (
    .I(__1458__),
    .O(__13__)
  );
  INV __3697__ (
    .I(__1411__),
    .O(__14__)
  );
  INV __3698__ (
    .I(__1407__),
    .O(__15__)
  );
  INV __3699__ (
    .I(__1426__),
    .O(__16__)
  );
  INV __3700__ (
    .I(__1424__),
    .O(__17__)
  );
  INV __3701__ (
    .I(__1422__),
    .O(__18__)
  );
  INV __3702__ (
    .I(__1419__),
    .O(__19__)
  );
  INV __3703__ (
    .I(__1417__),
    .O(__20__)
  );
  INV __3704__ (
    .I(__1432__),
    .O(__21__)
  );
  INV __3705__ (
    .I(__1430__),
    .O(__22__)
  );
  INV __3706__ (
    .I(__1428__),
    .O(__23__)
  );
  INV __3707__ (
    .I(__1444__),
    .O(__24__)
  );
  INV __3708__ (
    .I(__1442__),
    .O(__25__)
  );
  INV __3709__ (
    .I(__1440__),
    .O(__26__)
  );
  INV __3710__ (
    .I(__1438__),
    .O(__27__)
  );
  INV __3711__ (
    .I(__1436__),
    .O(__28__)
  );
  INV __3712__ (
    .I(__1450__),
    .O(__29__)
  );
  INV __3713__ (
    .I(__1448__),
    .O(__30__)
  );
  INV __3714__ (
    .I(__1446__),
    .O(__31__)
  );
  INV __3715__ (
    .I(__1150__),
    .O(__32__)
  );
  INV __3716__ (
    .I(__1148__),
    .O(__33__)
  );
  INV __3717__ (
    .I(__1146__),
    .O(__34__)
  );
  INV __3718__ (
    .I(__1144__),
    .O(__35__)
  );
  INV __3719__ (
    .I(__1142__),
    .O(__36__)
  );
  INV __3720__ (
    .I(__1140__),
    .O(__37__)
  );
  INV __3721__ (
    .I(__1118__),
    .O(__38__)
  );
  INV __3722__ (
    .I(__1115__),
    .O(__39__)
  );
  INV __3723__ (
    .I(__1112__),
    .O(__40__)
  );
  INV __3724__ (
    .I(__402__),
    .O(__41__)
  );
  INV __3725__ (
    .I(__400__),
    .O(__42__)
  );
  INV __3726__ (
    .I(__398__),
    .O(__43__)
  );
  INV __3727__ (
    .I(__396__),
    .O(__44__)
  );
  INV __3728__ (
    .I(__394__),
    .O(__45__)
  );
  INV __3729__ (
    .I(__392__),
    .O(__46__)
  );
  INV __3730__ (
    .I(__388__),
    .O(__47__)
  );
  INV __3731__ (
    .I(__386__),
    .O(__48__)
  );
  INV __3732__ (
    .I(__384__),
    .O(__49__)
  );
  INV __3733__ (
    .I(__1071__),
    .O(__50__)
  );
  INV __3734__ (
    .I(__1068__),
    .O(__51__)
  );
  INV __3735__ (
    .I(__1066__),
    .O(__52__)
  );
  INV __3736__ (
    .I(__1064__),
    .O(__53__)
  );
  INV __3737__ (
    .I(__413__),
    .O(__54__)
  );
  INV __3738__ (
    .I(__1063__),
    .O(__55__)
  );
  INV __3739__ (
    .I(__1091__),
    .O(__56__)
  );
  INV __3740__ (
    .I(__1060__),
    .O(__57__)
  );
  INV __3741__ (
    .I(__1058__),
    .O(__58__)
  );
  INV __3742__ (
    .I(__468__),
    .O(__59__)
  );
  INV __3743__ (
    .I(__378__),
    .O(__60__)
  );
  INV __3744__ (
    .I(__410__),
    .O(__61__)
  );
  INV __3745__ (
    .I(__381__),
    .O(__62__)
  );
  INV __3746__ (
    .I(__358__),
    .O(__63__)
  );
  INV __3747__ (
    .I(__479__),
    .O(__64__)
  );
  INV __3748__ (
    .I(__419__),
    .O(__65__)
  );
  INV __3749__ (
    .I(__504__),
    .O(__66__)
  );
  INV __3750__ (
    .I(__502__),
    .O(__67__)
  );
  INV __3751__ (
    .I(__3498__),
    .O(__68__)
  );
  INV __3752__ (
    .I(__3243__),
    .O(__69__)
  );
  INV __3753__ (
    .I(__3452__),
    .O(__70__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3754__ (
    .D(__2471__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__71__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3755__ (
    .D(__49__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__72__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3756__ (
    .D(__3023__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__73__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3757__ (
    .D(__48__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__74__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3758__ (
    .D(__47__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__75__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3759__ (
    .D(__46__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__76__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3760__ (
    .D(__3463__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__77__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3761__ (
    .D(__3241__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__78__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3762__ (
    .D(__3556__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__79__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3763__ (
    .D(__3017__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__80__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3764__ (
    .D(__2712__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__81__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3765__ (
    .D(__3197__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__82__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3766__ (
    .D(__2768__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__83__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3767__ (
    .D(__45__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__84__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3768__ (
    .D(__44__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__85__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3769__ (
    .D(__3460__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__86__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3770__ (
    .D(__2554__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__87__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3771__ (
    .D(__3563__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__88__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3772__ (
    .D(__3355__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__89__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3773__ (
    .D(__43__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__90__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3774__ (
    .D(__42__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__91__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3775__ (
    .D(__41__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__92__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3776__ (
    .D(__94__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__93__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3777__ (
    .D(__2559__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__94__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3778__ (
    .D(__2895__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__95__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3779__ (
    .D(__2650__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__96__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3780__ (
    .D(__2486__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__97__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3781__ (
    .D(__142__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__98__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3782__ (
    .D(__3084__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__99__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3783__ (
    .D(__2704__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__100__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3784__ (
    .D(__3234__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__101__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3785__ (
    .D(__2671__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__102__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3786__ (
    .D(__56__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__103__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3787__ (
    .D(__2473__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__104__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3788__ (
    .D(__3109__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__105__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3789__ (
    .D(__3327__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__106__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3790__ (
    .D(__2352__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__107__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3791__ (
    .D(__2059__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__108__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3792__ (
    .D(__3573__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__109__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3793__ (
    .D(__2578__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__110__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3794__ (
    .D(__1954__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__111__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3795__ (
    .D(__3629__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__112__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3796__ (
    .D(__3215__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__113__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3797__ (
    .D(__1628__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__114__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3798__ (
    .D(__3136__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__115__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3799__ (
    .D(__3546__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__116__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3800__ (
    .D(__2349__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__117__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3801__ (
    .D(__3209__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__118__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3802__ (
    .D(__2826__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__119__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3803__ (
    .D(__2625__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__120__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3804__ (
    .D(__3114__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__121__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3805__ (
    .D(__2096__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__122__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3806__ (
    .D(__3042__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__123__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3807__ (
    .D(__3182__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__124__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3808__ (
    .D(__1803__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__125__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3809__ (
    .D(__2174__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__126__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3810__ (
    .D(__3614__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__127__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3811__ (
    .D(__3033__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__128__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3812__ (
    .D(__3644__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__129__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3813__ (
    .D(__2971__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__130__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3814__ (
    .D(__2604__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__131__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3815__ (
    .D(__3549__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__132__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3816__ (
    .D(__3094__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__133__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3817__ (
    .D(__3387__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__134__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3818__ (
    .D(__2505__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__135__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3819__ (
    .D(__2677__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__136__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3820__ (
    .D(__3147__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__137__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3821__ (
    .D(__3584__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__138__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3822__ (
    .D(__3250__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__139__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3823__ (
    .D(__141__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__140__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3824__ (
    .D(__3554__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__141__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3825__ (
    .D(__143__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__142__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3826__ (
    .D(__2293__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__143__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3827__ (
    .D(__2178__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__144__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3828__ (
    .D(__3592__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__145__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3829__ (
    .D(__2426__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__146__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3830__ (
    .D(__3601__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__147__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3831__ (
    .D(__3126__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__148__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3832__ (
    .D(__3026__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__149__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3833__ (
    .D(__2497__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__150__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3834__ (
    .D(__2855__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__151__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3835__ (
    .D(__3282__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__152__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3836__ (
    .D(__3433__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__153__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3837__ (
    .D(__3624__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__154__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3838__ (
    .D(__3289__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__155__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3839__ (
    .D(__2664__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__156__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3840__ (
    .D(__3478__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__157__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3841__ (
    .D(__163__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__158__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3842__ (
    .D(__3403__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__159__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3843__ (
    .D(__3079__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__160__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3844__ (
    .D(__3008__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__161__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3845__ (
    .D(__2215__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__162__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3846__ (
    .D(__3401__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__163__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3847__ (
    .D(__3124__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__164__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3848__ (
    .D(__2308__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__165__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3849__ (
    .D(__3146__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__166__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3850__ (
    .D(__173__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__167__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3851__ (
    .D(__2201__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__168__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3852__ (
    .D(__1660__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__169__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3853__ (
    .D(__3575__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__170__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3854__ (
    .D(__2907__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__171__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3855__ (
    .D(__2852__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__172__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3856__ (
    .D(__176__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__173__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3857__ (
    .D(__3414__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__174__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3858__ (
    .D(__3357__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__175__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3859__ (
    .D(__1625__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__176__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3860__ (
    .D(__3048__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__177__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3861__ (
    .D(__2073__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__178__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3862__ (
    .D(__2758__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__179__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3863__ (
    .D(__3302__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__180__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3864__ (
    .D(__3291__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__181__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3865__ (
    .D(__3202__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__182__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3866__ (
    .D(__2923__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__183__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3867__ (
    .D(__3212__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__184__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3868__ (
    .D(__3313__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__185__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3869__ (
    .D(__3625__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__186__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3870__ (
    .D(__3411__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__187__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3871__ (
    .D(__3493__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__188__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3872__ (
    .D(__3415__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__189__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3873__ (
    .D(__3430__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__190__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3874__ (
    .D(__3492__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__191__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3875__ (
    .D(__3427__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__192__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3876__ (
    .D(__3591__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__193__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3877__ (
    .D(__2302__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__194__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3878__ (
    .D(__3586__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__195__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3879__ (
    .D(__2688__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__196__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3880__ (
    .D(__3576__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__197__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3881__ (
    .D(__3128__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__198__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3882__ (
    .D(__2696__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__199__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3883__ (
    .D(__1607__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__200__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3884__ (
    .D(__3626__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__201__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3885__ (
    .D(__2414__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__202__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3886__ (
    .D(__2437__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__203__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3887__ (
    .D(__2434__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__204__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3888__ (
    .D(__2781__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__205__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3889__ (
    .D(__2481__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__206__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3890__ (
    .D(__2878__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__207__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3891__ (
    .D(__2638__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__208__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3892__ (
    .D(__3181__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__209__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3893__ (
    .D(__3185__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__210__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3894__ (
    .D(__3660__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__211__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3895__ (
    .D(__3204__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__212__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3896__ (
    .D(__3550__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__213__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3897__ (
    .D(__2081__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__214__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3898__ (
    .D(__3441__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__215__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3899__ (
    .D(__3583__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__216__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3900__ (
    .D(__2157__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__217__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3901__ (
    .D(__3631__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__218__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3902__ (
    .D(__3417__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__219__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3903__ (
    .D(__3131__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__220__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3904__ (
    .D(__2807__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__221__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3905__ (
    .D(__3135__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__222__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3906__ (
    .D(__230__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__223__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3907__ (
    .D(__3439__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__224__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3908__ (
    .D(__3458__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__225__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3909__ (
    .D(__3148__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__226__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3910__ (
    .D(__3122__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__227__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3911__ (
    .D(__3391__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__228__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3912__ (
    .D(__2324__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__229__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3913__ (
    .D(__178__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__230__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3914__ (
    .D(__2025__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__231__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3915__ (
    .D(__3413__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__232__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3916__ (
    .D(__3428__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__233__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3917__ (
    .D(__64__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__234__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3918__ (
    .D(__3536__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__235__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3919__ (
    .D(__63__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__236__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3920__ (
    .D(__241__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__237__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3921__ (
    .D(__62__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__238__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3922__ (
    .D(__61__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__239__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3923__ (
    .D(__59__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__240__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3924__ (
    .D(__179__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__241__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3925__ (
    .D(__244__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__242__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3926__ (
    .D(__426__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__243__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3927__ (
    .D(__2580__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__244__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3928__ (
    .D(__2735__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__245__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3929__ (
    .D(__247__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__246__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3930__ (
    .D(__181__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__247__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3931__ (
    .D(__3300__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__248__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3932__ (
    .D(__345__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__249__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3933__ (
    .D(__311__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__250__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3934__ (
    .D(__348__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__251__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3935__ (
    .D(__353__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__252__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3936__ (
    .D(__727__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__253__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3937__ (
    .D(__1975__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__254__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3938__ (
    .D(__2643__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__255__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3939__ (
    .D(__257__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__256__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3940__ (
    .D(__191__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__257__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3941__ (
    .D(__259__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__258__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3942__ (
    .D(__195__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__259__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3943__ (
    .D(__261__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__260__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3944__ (
    .D(__196__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__261__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3945__ (
    .D(__263__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__262__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3946__ (
    .D(__265__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__263__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3947__ (
    .D(__3610__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__264__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3948__ (
    .D(__1947__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__265__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3949__ (
    .D(__2567__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__266__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3950__ (
    .D(__300__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__267__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3951__ (
    .D(__2606__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__268__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3952__ (
    .D(__3540__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__269__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3953__ (
    .D(__2494__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__270__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3954__ (
    .D(__2532__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__271__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3955__ (
    .D(__2504__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__272__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3956__ (
    .D(__1971__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__273__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3957__ (
    .D(__2145__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__274__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3958__ (
    .D(__3347__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__275__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3959__ (
    .D(__2121__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__276__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3960__ (
    .D(__1845__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__277__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3961__ (
    .D(__3117__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__278__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3962__ (
    .D(__2172__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__279__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3963__ (
    .D(__2748__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__280__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3964__ (
    .D(__3395__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__281__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3965__ (
    .D(__3647__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__282__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3966__ (
    .D(__3437__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__283__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3967__ (
    .D(__3561__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__284__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3968__ (
    .D(__3495__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__285__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3969__ (
    .D(__2245__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__286__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3970__ (
    .D(__3050__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__287__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3971__ (
    .D(__3436__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__288__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3972__ (
    .D(__3011__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__289__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3973__ (
    .D(__3339__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__290__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3974__ (
    .D(__3539__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__291__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3975__ (
    .D(__3203__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__292__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3976__ (
    .D(__3617__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__293__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3977__ (
    .D(__3205__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__294__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3978__ (
    .D(__1984__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__295__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3979__ (
    .D(__3623__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__296__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3980__ (
    .D(__299__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__297__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3981__ (
    .D(__3661__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__298__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3982__ (
    .D(__2566__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__299__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3983__ (
    .D(__301__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__300__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3984__ (
    .D(__3213__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__301__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3985__ (
    .D(__1784__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__302__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3986__ (
    .D(__305__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__303__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3987__ (
    .D(__2985__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__304__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3988__ (
    .D(__3666__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__305__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3989__ (
    .D(__307__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__306__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3990__ (
    .D(__308__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__307__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3991__ (
    .D(__1842__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__308__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3992__ (
    .D(__3520__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__309__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3993__ (
    .D(__2323__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__310__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3994__ (
    .D(__3038__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__311__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3995__ (
    .D(__313__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__312__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3996__ (
    .D(__625__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__313__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3997__ (
    .D(__315__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__314__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3998__ (
    .D(__627__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__315__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3999__ (
    .D(__317__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__316__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4000__ (
    .D(__628__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__317__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4001__ (
    .D(__319__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__318__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4002__ (
    .D(__629__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__319__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4003__ (
    .D(__321__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__320__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4004__ (
    .D(__630__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__321__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4005__ (
    .D(__323__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__322__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4006__ (
    .D(__631__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__323__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4007__ (
    .D(__325__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__324__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4008__ (
    .D(__632__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__325__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4009__ (
    .D(__327__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__326__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4010__ (
    .D(__633__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__327__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4011__ (
    .D(__329__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__328__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4012__ (
    .D(__634__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__329__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4013__ (
    .D(__331__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__330__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4014__ (
    .D(__635__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__331__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4015__ (
    .D(__333__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__332__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4016__ (
    .D(__636__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__333__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4017__ (
    .D(__335__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__334__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4018__ (
    .D(__637__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__335__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4019__ (
    .D(__2067__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__336__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4020__ (
    .D(__2851__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__337__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4021__ (
    .D(__3589__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__338__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4022__ (
    .D(__2078__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__339__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4023__ (
    .D(__2339__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__340__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4024__ (
    .D(__1114__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__341__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4025__ (
    .D(__3552__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__342__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4026__ (
    .D(__2205__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__343__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4027__ (
    .D(__2892__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__344__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4028__ (
    .D(__389__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__345__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4029__ (
    .D(__347__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__346__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4030__ (
    .D(__309__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__347__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4031__ (
    .D(__482__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__348__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4032__ (
    .D(__2171__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__349__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4033__ (
    .D(__351__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__350__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4034__ (
    .D(__422__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__351__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4035__ (
    .D(__379__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__352__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4036__ (
    .D(__254__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__353__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4037__ (
    .D(__2564__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__354__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4038__ (
    .D(__3542__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__355__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4039__ (
    .D(__2928__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__356__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4040__ (
    .D(__2893__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__357__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4041__ (
    .D(__420__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__358__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4042__ (
    .D(__3__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__359__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4043__ (
    .D(__8__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__360__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4044__ (
    .D(__2547__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__361__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4045__ (
    .D(__2913__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__362__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4046__ (
    .D(__2991__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__363__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4047__ (
    .D(__557__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__364__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4048__ (
    .D(__3371__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__365__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4049__ (
    .D(__3453__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__366__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4050__ (
    .D(__2459__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__367__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4051__ (
    .D(__602__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__368__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4052__ (
    .D(__67__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__369__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4053__ (
    .D(__2740__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__370__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4054__ (
    .D(__66__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__371__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4055__ (
    .D(__65__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__372__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4056__ (
    .D(__518__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__373__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4057__ (
    .D(__3579__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__374__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4058__ (
    .D(__60__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__375__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4059__ (
    .D(__2969__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__376__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4060__ (
    .D(__2292__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__377__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4061__ (
    .D(__530__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__378__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4062__ (
    .D(__1876__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__379__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4063__ (
    .D(__2254__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__380__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4064__ (
    .D(__409__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__381__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4065__ (
    .D(__3378__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__382__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4066__ (
    .D(__2279__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__383__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4067__ (
    .D(__385__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__384__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4068__ (
    .D(__1434__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__385__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4069__ (
    .D(__387__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__386__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4070__ (
    .D(__28__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__387__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4071__ (
    .D(__390__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__388__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4072__ (
    .D(__2450__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__389__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4073__ (
    .D(__27__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__390__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4074__ (
    .D(__3207__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__391__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4075__ (
    .D(__393__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__392__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4076__ (
    .D(__26__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__393__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4077__ (
    .D(__395__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__394__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4078__ (
    .D(__25__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__395__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4079__ (
    .D(__397__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__396__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4080__ (
    .D(__24__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__397__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4081__ (
    .D(__399__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__398__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4082__ (
    .D(__31__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__399__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4083__ (
    .D(__401__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__400__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4084__ (
    .D(__30__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__401__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4085__ (
    .D(__403__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__402__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4086__ (
    .D(__29__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__403__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4087__ (
    .D(__3599__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__404__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4088__ (
    .D(__3650__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__405__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4089__ (
    .D(__3382__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__406__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4090__ (
    .D(__2316__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__407__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4091__ (
    .D(__3299__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__408__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4092__ (
    .D(__14__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__409__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4093__ (
    .D(__466__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__410__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4094__ (
    .D(__3245__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__411__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4095__ (
    .D(__957__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__412__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4096__ (
    .D(__1029__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__413__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4097__ (
    .D(__3217__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__414__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4098__ (
    .D(__3388__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__415__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4099__ (
    .D(__1620__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__416__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4100__ (
    .D(__2000__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__417__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4101__ (
    .D(__2734__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__418__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4102__ (
    .D(__359__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__419__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4103__ (
    .D(__11__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__420__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4104__ (
    .D(__2857__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__421__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4105__ (
    .D(__3465__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__422__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4106__ (
    .D(__1631__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__423__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4107__ (
    .D(__2401__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__424__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4108__ (
    .D(__3528__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__425__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4109__ (
    .D(__3572__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__426__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4110__ (
    .D(__3214__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__427__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4111__ (
    .D(__3510__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__428__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4112__ (
    .D(__3316__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__429__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4113__ (
    .D(__2579__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__430__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4114__ (
    .D(__3019__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__431__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4115__ (
    .D(__3227__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__432__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4116__ (
    .D(__2835__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__433__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4117__ (
    .D(__2204__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__434__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4118__ (
    .D(__3494__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__435__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4119__ (
    .D(__2480__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__436__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4120__ (
    .D(__3604__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__437__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4121__ (
    .D(__3564__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__438__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4122__ (
    .D(__2544__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__439__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4123__ (
    .D(__3537__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__440__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4124__ (
    .D(__2672__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__441__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4125__ (
    .D(__1604__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__442__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4126__ (
    .D(__352__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__443__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4127__ (
    .D(__2782__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__444__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4128__ (
    .D(__2805__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__445__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4129__ (
    .D(__2868__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__446__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4130__ (
    .D(__2549__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__447__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4131__ (
    .D(__1636__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__448__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4132__ (
    .D(__3396__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__449__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4133__ (
    .D(__3322__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__450__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4134__ (
    .D(__3634__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__451__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4135__ (
    .D(__2590__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__452__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4136__ (
    .D(__3480__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__453__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4137__ (
    .D(__1734__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__454__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4138__ (
    .D(__2673__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__455__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4139__ (
    .D(__2275__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__456__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4140__ (
    .D(__3059__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__457__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4141__ (
    .D(__2133__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__458__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4142__ (
    .D(__3374__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__459__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4143__ (
    .D(__3474__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__460__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4144__ (
    .D(__2891__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__461__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4145__ (
    .D(__970__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__462__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4146__ (
    .D(__3568__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__463__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4147__ (
    .D(__3593__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__464__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4148__ (
    .D(__872__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__465__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4149__ (
    .D(__6__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__466__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4150__ (
    .D(__3504__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__467__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4151__ (
    .D(__508__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__468__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4152__ (
    .D(__3020__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__469__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4153__ (
    .D(__2841__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__470__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4154__ (
    .D(__3607__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__471__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4155__ (
    .D(__3068__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__472__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4156__ (
    .D(__2681__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__473__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4157__ (
    .D(__3069__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__474__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4158__ (
    .D(__2793__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__475__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4159__ (
    .D(__2207__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__476__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4160__ (
    .D(__1958__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__477__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4161__ (
    .D(__364__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__478__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4162__ (
    .D(__360__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__479__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4163__ (
    .D(__1779__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__480__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4164__ (
    .D(__510__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__481__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4165__ (
    .D(__2301__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__482__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4166__ (
    .D(__484__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__483__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4167__ (
    .D(__600__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__484__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4168__ (
    .D(__2806__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__485__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4169__ (
    .D(__250__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__486__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4170__ (
    .D(__558__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__487__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4171__ (
    .D(__489__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__488__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4172__ (
    .D(__601__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__489__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4173__ (
    .D(__491__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__490__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4174__ (
    .D(__559__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__491__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4175__ (
    .D(__493__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__492__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4176__ (
    .D(__211__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__493__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4177__ (
    .D(__513__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__494__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4178__ (
    .D(__368__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__495__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4179__ (
    .D(__578__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__496__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4180__ (
    .D(__498__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__497__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4181__ (
    .D(__562__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__498__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4182__ (
    .D(__3172__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__499__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4183__ (
    .D(__3294__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__500__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4184__ (
    .D(__2211__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__501__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4185__ (
    .D(__503__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__502__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4186__ (
    .D(__1405__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__503__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4187__ (
    .D(__505__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__504__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4188__ (
    .D(__15__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__505__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4189__ (
    .D(__2707__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__506__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4190__ (
    .D(__3680__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__507__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4191__ (
    .D(__9__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__508__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4192__ (
    .D(__3553__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__509__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4193__ (
    .D(__599__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__510__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4194__ (
    .D(__487__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__511__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4195__ (
    .D(__2519__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__512__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4196__ (
    .D(__560__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__513__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4197__ (
    .D(__2993__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__514__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4198__ (
    .D(__496__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__515__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4199__ (
    .D(__2206__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__516__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4200__ (
    .D(__2936__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__517__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4201__ (
    .D(__563__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__518__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4202__ (
    .D(__2935__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__519__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4203__ (
    .D(__2538__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__520__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4204__ (
    .D(__3360__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__521__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4205__ (
    .D(__2144__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__522__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4206__ (
    .D(__3179__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__523__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4207__ (
    .D(__2156__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__524__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4208__ (
    .D(__2739__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__525__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4209__ (
    .D(__3404__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__526__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4210__ (
    .D(__3287__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__527__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4211__ (
    .D(__3380__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__528__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4212__ (
    .D(__3585__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__529__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4213__ (
    .D(__4__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__530__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4214__ (
    .D(__2413__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__531__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4215__ (
    .D(__2964__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__532__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4216__ (
    .D(__2163__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__533__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4217__ (
    .D(__2476__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__534__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4218__ (
    .D(__3432__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__535__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4219__ (
    .D(__2803__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__536__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4220__ (
    .D(__3134__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__537__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4221__ (
    .D(__3053__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__538__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4222__ (
    .D(__3402__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__539__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4223__ (
    .D(__2761__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__540__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4224__ (
    .D(__2265__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__541__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4225__ (
    .D(__2281__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__542__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4226__ (
    .D(__3484__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__543__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4227__ (
    .D(__3447__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__544__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4228__ (
    .D(__3581__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__545__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4229__ (
    .D(__3312__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__546__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4230__ (
    .D(__3455__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__547__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4231__ (
    .D(__3184__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__548__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4232__ (
    .D(__2321__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__549__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4233__ (
    .D(__3605__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__550__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4234__ (
    .D(__3259__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__551__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4235__ (
    .D(__3547__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__552__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4236__ (
    .D(__2467__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__553__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4237__ (
    .D(__2674__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__554__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4238__ (
    .D(__2463__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__555__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4239__ (
    .D(__3086__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__556__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4240__ (
    .D(__3481__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__557__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4241__ (
    .D(__2371__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__558__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4242__ (
    .D(__2771__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__559__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4243__ (
    .D(__2563__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__560__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4244__ (
    .D(__3052__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__561__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4245__ (
    .D(__3675__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__562__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4246__ (
    .D(__3120__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__563__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4247__ (
    .D(__3473__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__564__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4248__ (
    .D(__2282__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__565__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4249__ (
    .D(__1813__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__566__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4250__ (
    .D(__3571__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__567__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4251__ (
    .D(__2600__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__568__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4252__ (
    .D(__660__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__569__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4253__ (
    .D(__3483__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__570__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4254__ (
    .D(__3318__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__571__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4255__ (
    .D(__2331__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__572__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4256__ (
    .D(__2683__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__573__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4257__ (
    .D(__2770__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__574__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4258__ (
    .D(__3665__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__575__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4259__ (
    .D(__2291__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__576__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4260__ (
    .D(__3280__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__577__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4261__ (
    .D(__3435__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__578__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4262__ (
    .D(__2598__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__579__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4263__ (
    .D(__1138__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__580__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4264__ (
    .D(__565__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__581__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4265__ (
    .D(__2177__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__582__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4266__ (
    .D(__3141__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__583__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4267__ (
    .D(__3063__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__584__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4268__ (
    .D(__3582__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__585__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4269__ (
    .D(__3656__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__586__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4270__ (
    .D(__2744__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__587__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4271__ (
    .D(__1022__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__588__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4272__ (
    .D(__662__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__589__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4273__ (
    .D(__3538__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__590__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4274__ (
    .D(__3558__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__591__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4275__ (
    .D(__1956__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__592__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4276__ (
    .D(__3255__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__593__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4277__ (
    .D(__2091__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__594__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4278__ (
    .D(__2983__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__595__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4279__ (
    .D(__3340__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__596__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4280__ (
    .D(__2213__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__597__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4281__ (
    .D(__3383__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__598__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4282__ (
    .D(__3113__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__599__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4283__ (
    .D(__2289__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__600__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4284__ (
    .D(__2428__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__601__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4285__ (
    .D(__3663__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__602__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4286__ (
    .D(__581__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__603__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4287__ (
    .D(__2152__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__604__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4288__ (
    .D(__3256__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__605__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4289__ (
    .D(__3502__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__606__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4290__ (
    .D(__2170__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__607__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4291__ (
    .D(__2296__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__608__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4292__ (
    .D(__1963__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__609__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4293__ (
    .D(__3070__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__610__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4294__ (
    .D(__3560__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__611__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4295__ (
    .D(__2752__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__612__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4296__ (
    .D(__3674__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__613__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4297__ (
    .D(__3211__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__614__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4298__ (
    .D(__2933__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__615__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4299__ (
    .D(__2574__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__616__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4300__ (
    .D(__2557__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__617__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4301__ (
    .D(__2836__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__618__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4302__ (
    .D(__2283__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__619__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4303__ (
    .D(__919__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__620__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4304__ (
    .D(__2513__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__621__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4305__ (
    .D(__2299__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__622__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4306__ (
    .D(__2741__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__623__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4307__ (
    .D(__2755__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__624__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4308__ (
    .D(__2775__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__625__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4309__ (
    .D(__2083__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__626__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4310__ (
    .D(__2072__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__627__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4311__ (
    .D(__3652__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__628__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4312__ (
    .D(__3630__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__629__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4313__ (
    .D(__2989__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__630__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4314__ (
    .D(__2583__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__631__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4315__ (
    .D(__3165__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__632__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4316__ (
    .D(__2295__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__633__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4317__ (
    .D(__2990__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__634__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4318__ (
    .D(__3406__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__635__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4319__ (
    .D(__2789__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__636__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4320__ (
    .D(__3040__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__637__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4321__ (
    .D(__3228__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__638__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4322__ (
    .D(__3025__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__639__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4323__ (
    .D(__3570__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__640__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4324__ (
    .D(__3477__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__641__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4325__ (
    .D(__3574__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__642__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4326__ (
    .D(__2592__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__643__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4327__ (
    .D(__3132__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__644__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4328__ (
    .D(__2979__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__645__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4329__ (
    .D(__3673__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__646__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4330__ (
    .D(__3497__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__647__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4331__ (
    .D(__2988__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__648__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4332__ (
    .D(__2572__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__649__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4333__ (
    .D(__1018__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__650__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4334__ (
    .D(__2491__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__651__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4335__ (
    .D(__2794__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__652__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4336__ (
    .D(__1849__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__653__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4337__ (
    .D(__3111__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__654__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4338__ (
    .D(__3503__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__655__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4339__ (
    .D(__1848__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__656__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4340__ (
    .D(__3116__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__657__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4341__ (
    .D(__2854__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__658__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4342__ (
    .D(__3390__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__659__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4343__ (
    .D(__1137__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__660__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4344__ (
    .D(__2168__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__661__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4345__ (
    .D(__663__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__662__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4346__ (
    .D(__1494__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__663__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4347__ (
    .D(__2274__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__664__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4348__ (
    .D(__3279__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__665__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4349__ (
    .D(__3133__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__666__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4350__ (
    .D(__2910__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__667__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4351__ (
    .D(__2675__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__668__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4352__ (
    .D(__3345__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__669__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4353__ (
    .D(__2521__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__670__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4354__ (
    .D(__1840__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__671__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4355__ (
    .D(__2757__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__672__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4356__ (
    .D(__2575__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__673__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4357__ (
    .D(__3252__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__674__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4358__ (
    .D(__2310__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__675__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4359__ (
    .D(__3602__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__676__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4360__ (
    .D(__3200__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__677__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4361__ (
    .D(__2495__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__678__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4362__ (
    .D(__3129__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__679__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4363__ (
    .D(__3029__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__680__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4364__ (
    .D(__1988__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__681__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4365__ (
    .D(__3682__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__682__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4366__ (
    .D(__2330__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__683__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4367__ (
    .D(__2541__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__684__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4368__ (
    .D(__3359__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__685__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4369__ (
    .D(__2987__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__686__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4370__ (
    .D(__3105__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__687__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4371__ (
    .D(__2454__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__688__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4372__ (
    .D(__2531__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__689__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4373__ (
    .D(__3292__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__690__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4374__ (
    .D(__2615__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__691__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4375__ (
    .D(__2545__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__692__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4376__ (
    .D(__2693__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__693__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4377__ (
    .D(__2862__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__694__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4378__ (
    .D(__3679__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__695__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4379__ (
    .D(__3442__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__696__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4380__ (
    .D(__2786__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__697__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4381__ (
    .D(__3423__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__698__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4382__ (
    .D(__2273__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__699__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4383__ (
    .D(__1990__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__700__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4384__ (
    .D(__3468__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__701__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4385__ (
    .D(__2616__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__702__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4386__ (
    .D(__2356__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__703__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4387__ (
    .D(__2202__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__704__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4388__ (
    .D(__3092__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__705__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4389__ (
    .D(__3490__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__706__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4390__ (
    .D(__3190__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__707__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4391__ (
    .D(__2358__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__708__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4392__ (
    .D(__3543__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__709__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4393__ (
    .D(__3326__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__710__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4394__ (
    .D(__3594__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__711__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4395__ (
    .D(__2527__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__712__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4396__ (
    .D(__2745__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__713__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4397__ (
    .D(__3027__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__714__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4398__ (
    .D(__2996__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__715__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4399__ (
    .D(__2890__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__716__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4400__ (
    .D(__2802__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__717__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4401__ (
    .D(__2485__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__718__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4402__ (
    .D(__3051__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__719__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4403__ (
    .D(__3533__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__720__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4404__ (
    .D(__3475__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__721__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4405__ (
    .D(__2368__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__722__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4406__ (
    .D(__2588__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__723__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4407__ (
    .D(__1866__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__724__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4408__ (
    .D(__3323__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__725__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4409__ (
    .D(__2864__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__726__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4410__ (
    .D(__1131__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__727__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4411__ (
    .D(__2785__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__728__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4412__ (
    .D(__3206__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__729__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4413__ (
    .D(__2925__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__730__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4414__ (
    .D(__2294__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__731__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4415__ (
    .D(__2565__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__732__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4416__ (
    .D(__956__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__733__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4417__ (
    .D(__2773__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__734__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4418__ (
    .D(__3419__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__735__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4419__ (
    .D(__3389__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__736__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4420__ (
    .D(__3226__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__737__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4421__ (
    .D(__3344__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__738__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4422__ (
    .D(__2020__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__739__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4423__ (
    .D(__2760__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__740__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4424__ (
    .D(__1987__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__741__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4425__ (
    .D(__3551__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__742__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4426__ (
    .D(__3103__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__743__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4427__ (
    .D(__3464__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__744__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4428__ (
    .D(__2399__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__745__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4429__ (
    .D(__3309__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__746__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4430__ (
    .D(__2060__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__747__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4431__ (
    .D(__2624__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__748__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4432__ (
    .D(__3297__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__749__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4433__ (
    .D(__3093__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__750__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4434__ (
    .D(__2751__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__751__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4435__ (
    .D(__2093__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__752__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4436__ (
    .D(__2986__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__753__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4437__ (
    .D(__58__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__754__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4438__ (
    .D(__57__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__755__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4439__ (
    .D(__2449__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__756__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4440__ (
    .D(__2605__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__757__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4441__ (
    .D(__54__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__758__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4442__ (
    .D(__53__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__759__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4443__ (
    .D(__2466__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__760__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4444__ (
    .D(__52__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__761__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4445__ (
    .D(__51__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__762__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4446__ (
    .D(__50__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__763__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4447__ (
    .D(__771__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__764__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4448__ (
    .D(__2863__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__765__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4449__ (
    .D(__3527__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__766__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4450__ (
    .D(__2614__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__767__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4451__ (
    .D(__2253__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__768__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4452__ (
    .D(__55__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__769__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4453__ (
    .D(__2879__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__770__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4454__ (
    .D(__2560__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__771__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4455__ (
    .D(__3671__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__772__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4456__ (
    .D(__1026__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__773__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4457__ (
    .D(__2430__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__774__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4458__ (
    .D(__2611__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__775__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4459__ (
    .D(__3278__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__776__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4460__ (
    .D(__3397__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__777__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4461__ (
    .D(__3668__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__778__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4462__ (
    .D(__3446__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__779__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4463__ (
    .D(__2350__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__780__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4464__ (
    .D(__3628__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__781__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4465__ (
    .D(__2451__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__782__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4466__ (
    .D(__3511__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__783__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4467__ (
    .D(__2589__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__784__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4468__ (
    .D(__2911__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__785__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4469__ (
    .D(__3189__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__786__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4470__ (
    .D(__3112__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__787__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4471__ (
    .D(__2780__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__788__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4472__ (
    .D(__3578__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__789__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4473__ (
    .D(__2456__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__790__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4474__ (
    .D(__3531__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__791__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4475__ (
    .D(__3044__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__792__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4476__ (
    .D(__3627__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__793__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4477__ (
    .D(__3467__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__794__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4478__ (
    .D(__2496__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__795__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4479__ (
    .D(__2548__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__796__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4480__ (
    .D(__1847__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__797__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4481__ (
    .D(__3296__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__798__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4482__ (
    .D(__2798__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__799__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4483__ (
    .D(__3377__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__800__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4484__ (
    .D(__3530__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__801__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4485__ (
    .D(__3363__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__802__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4486__ (
    .D(__2561__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__803__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4487__ (
    .D(__3284__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__804__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4488__ (
    .D(__3180__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__805__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4489__ (
    .D(__2976__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__806__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4490__ (
    .D(__3192__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__807__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4491__ (
    .D(__2398__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__808__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4492__ (
    .D(__3615__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__809__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4493__ (
    .D(__3251__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__810__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4494__ (
    .D(__1666__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__811__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4495__ (
    .D(__1846__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__812__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4496__ (
    .D(__3281__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__813__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4497__ (
    .D(__3145__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__814__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4498__ (
    .D(__2452__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__815__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4499__ (
    .D(__1654__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__816__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4500__ (
    .D(__3580__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__817__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4501__ (
    .D(__3379__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__818__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4502__ (
    .D(__2917__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__819__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4503__ (
    .D(__2300__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__820__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4504__ (
    .D(__3422__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__821__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4505__ (
    .D(__3286__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__822__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4506__ (
    .D(__3426__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__823__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4507__ (
    .D(__2129__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__824__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4508__ (
    .D(__3021__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__825__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4509__ (
    .D(__3110__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__826__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4510__ (
    .D(__3664__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__827__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4511__ (
    .D(__2080__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__828__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4512__ (
    .D(__2329__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__829__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4513__ (
    .D(__2128__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__830__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4514__ (
    .D(__3434__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__831__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4515__ (
    .D(__3471__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__832__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4516__ (
    .D(__2562__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__833__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4517__ (
    .D(__2700__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__834__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4518__ (
    .D(__3535__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__835__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4519__ (
    .D(__3037__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__836__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4520__ (
    .D(__3443__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__837__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4521__ (
    .D(__3138__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__838__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4522__ (
    .D(__2457__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__839__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4523__ (
    .D(__2465__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__840__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4524__ (
    .D(__2252__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__841__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4525__ (
    .D(__3619__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__842__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4526__ (
    .D(__3041__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__843__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4527__ (
    .D(__3369__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__844__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4528__ (
    .D(__2599__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__845__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4529__ (
    .D(__2799__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__846__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4530__ (
    .D(__2433__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__847__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4531__ (
    .D(__868__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__848__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4532__ (
    .D(__2922__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__849__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4533__ (
    .D(__3001__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__850__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4534__ (
    .D(__3276__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__851__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4535__ (
    .D(__2997__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__852__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4536__ (
    .D(__3394__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__853__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4537__ (
    .D(__3277__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__854__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4538__ (
    .D(__3534__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__855__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4539__ (
    .D(__2242__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__856__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4540__ (
    .D(__2154__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__857__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4541__ (
    .D(__215__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__858__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4542__ (
    .D(__3407__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__859__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4543__ (
    .D(__1605__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__860__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4544__ (
    .D(__2750__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__861__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4545__ (
    .D(__870__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__862__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4546__ (
    .D(__2270__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__863__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4547__ (
    .D(__3608__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__864__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4548__ (
    .D(__2053__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__865__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4549__ (
    .D(__3004__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__866__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4550__ (
    .D(__860__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__867__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4551__ (
    .D(__377__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__868__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4552__ (
    .D(__1966__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__869__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4553__ (
    .D(__2869__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__870__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4554__ (
    .D(__3350__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__871__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4555__ (
    .D(__873__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__872__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4556__ (
    .D(__1663__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__873__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4557__ (
    .D(__2332__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__874__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4558__ (
    .D(__1630__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__875__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4559__ (
    .D(__3024__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__876__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4560__ (
    .D(__1675__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__877__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4561__ (
    .D(__3499__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__878__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4562__ (
    .D(__3022__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__879__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4563__ (
    .D(__3485__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__880__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4564__ (
    .D(__2980__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__881__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4565__ (
    .D(__2754__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__882__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4566__ (
    .D(__2656__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__883__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4567__ (
    .D(__2535__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__884__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4568__ (
    .D(__3137__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__885__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4569__ (
    .D(__2546__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__886__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4570__ (
    .D(__2492__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__887__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4571__ (
    .D(__1815__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__888__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4572__ (
    .D(__3544__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__889__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4573__ (
    .D(__2833__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__890__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4574__ (
    .D(__2340__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__891__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4575__ (
    .D(__2926__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__892__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4576__ (
    .D(__3655__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__893__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4577__ (
    .D(__3598__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__894__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4578__ (
    .D(__2533__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__895__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4579__ (
    .D(__2079__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__896__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4580__ (
    .D(__2266__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__897__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4581__ (
    .D(__3028__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__898__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4582__ (
    .D(__2403__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__899__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4583__ (
    .D(__3541__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__900__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4584__ (
    .D(__2284__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__901__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4585__ (
    .D(__3662__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__902__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4586__ (
    .D(__1676__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__903__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4587__ (
    .D(__2778__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__904__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4588__ (
    .D(__3431__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__905__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4589__ (
    .D(__1991__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__906__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4590__ (
    .D(__2966__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__907__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4591__ (
    .D(__3035__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__908__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4592__ (
    .D(__2872__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__909__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4593__ (
    .D(__3448__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__910__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4594__ (
    .D(__3080__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__911__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4595__ (
    .D(__1870__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__912__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4596__ (
    .D(__2320__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__913__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4597__ (
    .D(__1970__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__914__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4598__ (
    .D(__2777__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__915__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4599__ (
    .D(__2699__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__916__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4600__ (
    .D(__2747__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__917__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4601__ (
    .D(__3454__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__918__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4602__ (
    .D(__1130__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__919__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4603__ (
    .D(__2162__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__920__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4604__ (
    .D(__2603__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__921__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4605__ (
    .D(__948__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__922__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4606__ (
    .D(__1023__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__923__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4607__ (
    .D(__3288__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__924__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4608__ (
    .D(__3257__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__925__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4609__ (
    .D(__40__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__926__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4610__ (
    .D(__3506__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__927__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4611__ (
    .D(__39__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__928__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4612__ (
    .D(__38__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__929__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4613__ (
    .D(__37__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__930__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4614__ (
    .D(__36__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__931__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4615__ (
    .D(__35__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__932__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4616__ (
    .D(__34__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__933__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4617__ (
    .D(__33__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__934__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4618__ (
    .D(__32__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__935__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4619__ (
    .D(__937__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__936__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4620__ (
    .D(__2558__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__937__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4621__ (
    .D(__2429__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__938__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4622__ (
    .D(__988__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__939__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4623__ (
    .D(__3258__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__940__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4624__ (
    .D(__2968__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__941__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4625__ (
    .D(__2703__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__942__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4626__ (
    .D(__3559__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__943__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4627__ (
    .D(__954__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__944__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4628__ (
    .D(__2127__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__945__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4629__ (
    .D(__3095__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__946__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4630__ (
    .D(__2695__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__947__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4631__ (
    .D(__857__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__948__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4632__ (
    .D(__3361__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__949__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4633__ (
    .D(__2__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__950__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4634__ (
    .D(__2052__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__951__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4635__ (
    .D(__2024__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__952__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4636__ (
    .D(__2303__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__953__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4637__ (
    .D(__858__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__954__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4638__ (
    .D(__2796__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__955__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4639__ (
    .D(__1132__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__956__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4640__ (
    .D(__784__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__957__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4641__ (
    .D(__959__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__958__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4642__ (
    .D(__782__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__959__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4643__ (
    .D(__961__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__960__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4644__ (
    .D(__433__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__961__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4645__ (
    .D(__963__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__962__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4646__ (
    .D(__442__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__963__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4647__ (
    .D(__243__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__964__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4648__ (
    .D(__966__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__965__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4649__ (
    .D(__967__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__966__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4650__ (
    .D(__2392__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__967__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4651__ (
    .D(__1659__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__968__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4652__ (
    .D(__3399__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__969__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4653__ (
    .D(__1129__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__970__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4654__ (
    .D(__2577__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__971__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4655__ (
    .D(__2984__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__972__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4656__ (
    .D(__2530__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__973__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4657__ (
    .D(__2909__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__974__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4658__ (
    .D(__2694__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__975__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4659__ (
    .D(__2490__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__976__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4660__ (
    .D(__3368__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__977__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4661__ (
    .D(__3600__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__978__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4662__ (
    .D(__3065__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__979__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4663__ (
    .D(__2135__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__980__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4664__ (
    .D(__1811__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__981__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4665__ (
    .D(__3476__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__982__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4666__ (
    .D(__3125__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__983__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4667__ (
    .D(__3616__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__984__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4668__ (
    .D(__2963__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__985__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4669__ (
    .D(__987__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__986__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4670__ (
    .D(__2678__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__987__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4671__ (
    .D(__989__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__988__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4672__ (
    .D(__3032__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__989__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4673__ (
    .D(__1781__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__990__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4674__ (
    .D(__992__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__991__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4675__ (
    .D(__3014__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__992__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4676__ (
    .D(__994__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__993__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4677__ (
    .D(__995__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__994__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4678__ (
    .D(__2021__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__995__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4679__ (
    .D(__3409__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__996__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4680__ (
    .D(__3595__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__997__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4681__ (
    .D(__3246__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__998__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4682__ (
    .D(__1673__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__999__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4683__ (
    .D(__2074__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1000__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4684__ (
    .D(__3064__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1001__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4685__ (
    .D(__1814__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1002__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4686__ (
    .D(__2529__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1003__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4687__ (
    .D(__3587__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1004__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4688__ (
    .D(__2506__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1005__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4689__ (
    .D(__1661__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1006__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4690__ (
    .D(__3424__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1007__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4691__ (
    .D(__2432__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1008__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4692__ (
    .D(__2834__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1009__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4693__ (
    .D(__3526__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1010__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4694__ (
    .D(__1012__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1011__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4695__ (
    .D(__996__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1012__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4696__ (
    .D(__1014__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1013__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4697__ (
    .D(__997__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1014__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4698__ (
    .D(__1016__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1015__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4699__ (
    .D(__998__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1016__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4700__ (
    .D(__1021__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1017__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4701__ (
    .D(__1134__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1018__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4702__ (
    .D(__1020__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1019__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4703__ (
    .D(__1135__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1020__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4704__ (
    .D(__1005__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1021__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4705__ (
    .D(__1136__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1022__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4706__ (
    .D(__1133__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1023__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4707__ (
    .D(__1025__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1024__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4708__ (
    .D(__1006__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1025__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4709__ (
    .D(__1139__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1026__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4710__ (
    .D(__3519__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1027__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4711__ (
    .D(__1032__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1028__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4712__ (
    .D(__1__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1029__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4713__ (
    .D(__580__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1030__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4714__ (
    .D(__341__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1031__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4715__ (
    .D(__1007__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1032__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4716__ (
    .D(__1034__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1033__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4717__ (
    .D(__1035__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1034__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4718__ (
    .D(__2046__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1035__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4719__ (
    .D(__3343__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1036__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4720__ (
    .D(__3488__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1037__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4721__ (
    .D(__2077__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1038__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4722__ (
    .D(__1041__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1039__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4723__ (
    .D(__3392__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1040__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4724__ (
    .D(__1196__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1041__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4725__ (
    .D(__2458__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1042__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4726__ (
    .D(__2373__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1043__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4727__ (
    .D(__2017__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1044__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4728__ (
    .D(__3031__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1045__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4729__ (
    .D(__2479__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1046__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4730__ (
    .D(__1669__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1047__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4731__ (
    .D(__3532__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1048__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4732__ (
    .D(__1671__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1049__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4733__ (
    .D(__3367__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1050__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4734__ (
    .D(__3501__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1051__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4735__ (
    .D(__1053__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1052__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4736__ (
    .D(__1197__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1053__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4737__ (
    .D(__2776__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1054__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4738__ (
    .D(__3678__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1055__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4739__ (
    .D(__2914__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1056__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4740__ (
    .D(__2249__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1057__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4741__ (
    .D(__1090__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1058__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4742__ (
    .D(__1069__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1059__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4743__ (
    .D(__1061__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1060__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4744__ (
    .D(__7__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1061__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4745__ (
    .D(__5__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1062__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4746__ (
    .D(__950__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1063__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4747__ (
    .D(__1065__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1064__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4748__ (
    .D(__0__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1065__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4749__ (
    .D(__1067__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1066__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4750__ (
    .D(__13__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1067__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4751__ (
    .D(__1070__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1068__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4752__ (
    .D(__1199__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1069__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4753__ (
    .D(__12__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1070__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4754__ (
    .D(__1072__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1071__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4755__ (
    .D(__10__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1072__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4756__ (
    .D(__3039__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1073__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4757__ (
    .D(__1974__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1074__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4758__ (
    .D(__3676__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1075__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4759__ (
    .D(__1079__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1076__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4760__ (
    .D(__1924__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1077__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4761__ (
    .D(__2478__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1078__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4762__ (
    .D(__1206__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1079__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4763__ (
    .D(__3047__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1080__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4764__ (
    .D(__2766__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1081__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4765__ (
    .D(__1085__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1082__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4766__ (
    .D(__2787__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1083__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4767__ (
    .D(__3315__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1084__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4768__ (
    .D(__1208__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1085__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4769__ (
    .D(__3567__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1086__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4770__ (
    .D(__1089__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1087__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4771__ (
    .D(__3106__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1088__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4772__ (
    .D(__1209__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1089__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4773__ (
    .D(__1452__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1090__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4774__ (
    .D(__1062__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1091__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4775__ (
    .D(__1093__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1092__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4776__ (
    .D(__1210__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1093__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4777__ (
    .D(__1095__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1094__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4778__ (
    .D(__1211__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1095__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4779__ (
    .D(__1097__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1096__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4780__ (
    .D(__1212__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1097__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4781__ (
    .D(__1099__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1098__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4782__ (
    .D(__1214__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1099__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4783__ (
    .D(__1101__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1100__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4784__ (
    .D(__1215__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1101__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4785__ (
    .D(__1618__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1102__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4786__ (
    .D(__1104__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1103__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4787__ (
    .D(__1219__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1104__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4788__ (
    .D(__3225__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1105__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4789__ (
    .D(__2468__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1106__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4790__ (
    .D(__3164__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1107__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4791__ (
    .D(__2251__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1108__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4792__ (
    .D(__2487__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1109__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4793__ (
    .D(__2161__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1110__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4794__ (
    .D(__1672__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1111__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4795__ (
    .D(__1113__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1112__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4796__ (
    .D(__1415__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1113__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4797__ (
    .D(__2618__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1114__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4798__ (
    .D(__1116__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1115__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4799__ (
    .D(__20__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1116__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4800__ (
    .D(__3505__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1117__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4801__ (
    .D(__1121__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1118__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4802__ (
    .D(__2662__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1119__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4803__ (
    .D(__3261__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1120__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4804__ (
    .D(__19__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1121__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4805__ (
    .D(__2418__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1122__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4806__ (
    .D(__3487__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1123__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4807__ (
    .D(__2400__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1124__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4808__ (
    .D(__2493__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1125__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4809__ (
    .D(__3622__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1126__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4810__ (
    .D(__2772__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1127__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4811__ (
    .D(__3405__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1128__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4812__ (
    .D(__2169__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1129__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4813__ (
    .D(__3186__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1130__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4814__ (
    .D(__3645__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1131__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4815__ (
    .D(__3045__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1132__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4816__ (
    .D(__1634__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1133__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4817__ (
    .D(__3144__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1134__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4818__ (
    .D(__1603__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1135__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4819__ (
    .D(__3524__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1136__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4820__ (
    .D(__2871__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1137__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4821__ (
    .D(__3681__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1138__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4822__ (
    .D(__3646__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1139__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4823__ (
    .D(__1141__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1140__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4824__ (
    .D(__18__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1141__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4825__ (
    .D(__1143__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1142__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4826__ (
    .D(__17__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1143__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4827__ (
    .D(__1145__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1144__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4828__ (
    .D(__16__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1145__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4829__ (
    .D(__1147__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1146__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4830__ (
    .D(__23__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1147__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4831__ (
    .D(__1149__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1148__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4832__ (
    .D(__22__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1149__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4833__ (
    .D(__1151__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1150__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4834__ (
    .D(__21__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1151__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4835__ (
    .D(__2217__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1152__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4836__ (
    .D(__2659__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1153__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4837__ (
    .D(__2918__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1154__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4838__ (
    .D(__2448__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1155__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4839__ (
    .D(__2602__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1156__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4840__ (
    .D(__2698__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1157__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4841__ (
    .D(__2642__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1158__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4842__ (
    .D(__2853__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1159__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4843__ (
    .D(__3509__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1160__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4844__ (
    .D(__3293__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1161__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4845__ (
    .D(__3522__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1162__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4846__ (
    .D(__3523__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1163__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4847__ (
    .D(__1875__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1164__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4848__ (
    .D(__3253__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1165__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4849__ (
    .D(__3425__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1166__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4850__ (
    .D(__2726__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1167__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4851__ (
    .D(__2622__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1168__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4852__ (
    .D(__3260__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1169__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4853__ (
    .D(__3314__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1170__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4854__ (
    .D(__2967__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1171__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4855__ (
    .D(__2406__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1172__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4856__ (
    .D(__2982__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1173__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4857__ (
    .D(__3496__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1174__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4858__ (
    .D(__2800__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1175__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4859__ (
    .D(__2304__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1176__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4860__ (
    .D(__3249__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1177__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4861__ (
    .D(__2705__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1178__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4862__ (
    .D(__2542__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1179__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4863__ (
    .D(__3254__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1180__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4864__ (
    .D(__2453__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1181__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4865__ (
    .D(__2365__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1182__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4866__ (
    .D(__1645__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1183__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4867__ (
    .D(__3649__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1184__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4868__ (
    .D(__3545__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1185__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4869__ (
    .D(__3529__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1186__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4870__ (
    .D(__3472__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1187__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4871__ (
    .D(__2840__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1188__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4872__ (
    .D(__2861__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1189__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4873__ (
    .D(__3648__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1190__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4874__ (
    .D(__2511__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1191__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4875__ (
    .D(__2930__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1192__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4876__ (
    .D(__2663__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1193__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4877__ (
    .D(__2586__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1194__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4878__ (
    .D(__3194__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1195__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4879__ (
    .D(__3187__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1196__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4880__ (
    .D(__3071__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1197__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4881__ (
    .D(__3421__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1198__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4882__ (
    .D(__3486__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1199__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4883__ (
    .D(__3466__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1200__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4884__ (
    .D(__2792__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1201__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4885__ (
    .D(__3013__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1202__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4886__ (
    .D(__3348__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1203__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4887__ (
    .D(__3429__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1204__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4888__ (
    .D(__3054__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1205__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4889__ (
    .D(__3461__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1206__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4890__ (
    .D(__2517__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1207__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4891__ (
    .D(__2680__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1208__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4892__ (
    .D(__2702__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1209__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4893__ (
    .D(__2066__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1210__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4894__ (
    .D(__2569__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1211__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4895__ (
    .D(__3060__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1212__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4896__ (
    .D(__2328__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1213__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4897__ (
    .D(__2882__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1214__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4898__ (
    .D(__3290__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1215__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4899__ (
    .D(__3557__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1216__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4900__ (
    .D(__3139__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1217__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4901__ (
    .D(__3512__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1218__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4902__ (
    .D(__3410__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1219__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4903__ (
    .D(__2715__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1220__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4904__ (
    .D(__3613__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1221__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4905__ (
    .D(__3301__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1222__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4906__ (
    .D(__2311__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1223__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4907__ (
    .D(__2839__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1224__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4908__ (
    .D(__3590__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1225__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4909__ (
    .D(__3393__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1226__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4910__ (
    .D(__3365__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1227__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4911__ (
    .D(__3621__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1228__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4912__ (
    .D(__2837__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1229__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4913__ (
    .D(__3375__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1230__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4914__ (
    .D(__3606__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1231__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4915__ (
    .D(__2076__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1232__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4916__ (
    .D(__2408__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1233__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4917__ (
    .D(__3440__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1234__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4918__ (
    .D(__2998__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1235__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4919__ (
    .D(__2472__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1236__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4920__ (
    .D(__2880__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1237__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4921__ (
    .D(__3338__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1238__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4922__ (
    .D(__3670__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1239__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4923__ (
    .D(__2691__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1240__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4924__ (
    .D(__2716__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1241__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4925__ (
    .D(__1969__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1242__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4926__ (
    .D(__3321__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1243__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4927__ (
    .D(__2539__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1244__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4928__ (
    .D(__3199__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1245__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4929__ (
    .D(__2887__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1246__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4930__ (
    .D(__3308__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1247__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4931__ (
    .D(__2934__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1248__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4932__ (
    .D(__2338__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1249__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4933__ (
    .D(__1658__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1250__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4934__ (
    .D(__2844__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1251__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4935__ (
    .D(__3362__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1252__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4936__ (
    .D(__2654__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1253__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4937__ (
    .D(__2528__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1254__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4938__ (
    .D(__1594__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1255__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4939__ (
    .D(__3400__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1256__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4940__ (
    .D(__3376__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1257__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4941__ (
    .D(__3609__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1258__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4942__ (
    .D(__2804__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1259__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4943__ (
    .D(__2576__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1260__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4944__ (
    .D(__2995__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1261__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4945__ (
    .D(__3295__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1262__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4946__ (
    .D(__2147__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1263__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4947__ (
    .D(__3305__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1264__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4948__ (
    .D(__3372__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1265__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4949__ (
    .D(__1955__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1266__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4950__ (
    .D(__2710__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1267__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4951__ (
    .D(__3104__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1268__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4952__ (
    .D(__2932__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1269__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4953__ (
    .D(__2687__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1270__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4954__ (
    .D(__3358__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1271__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4955__ (
    .D(__3210__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1272__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4956__ (
    .D(__2609__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1273__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4957__ (
    .D(__1873__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1274__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4958__ (
    .D(__2717__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1275__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4959__ (
    .D(__1989__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1276__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4960__ (
    .D(__3479__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1277__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4961__ (
    .D(__2884__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1278__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4962__ (
    .D(__2587__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1279__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4963__ (
    .D(__2160__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1280__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4964__ (
    .D(__2858__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1281__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4965__ (
    .D(__2534__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1282__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4966__ (
    .D(__3036__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1283__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4967__ (
    .D(__3242__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1284__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4968__ (
    .D(__2416__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1285__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4969__ (
    .D(__1965__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1286__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4970__ (
    .D(__3230__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1287__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4971__ (
    .D(__3653__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1288__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4972__ (
    .D(__1841__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1289__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4973__ (
    .D(__2243__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1290__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4974__ (
    .D(__2123__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1291__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4975__ (
    .D(__2655__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1292__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4976__ (
    .D(__3325__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1293__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4977__ (
    .D(__2718__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1294__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4978__ (
    .D(__2351__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1295__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4979__ (
    .D(__3566__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1296__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4980__ (
    .D(__3009__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1297__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4981__ (
    .D(__3618__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1298__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4982__ (
    .D(__2061__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1299__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4983__ (
    .D(__2488__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1300__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4984__ (
    .D(__2920__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1301__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4985__ (
    .D(__3195__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1302__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4986__ (
    .D(__3030__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1303__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4987__ (
    .D(__2415__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1304__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4988__ (
    .D(__2097__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1305__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4989__ (
    .D(__3525__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1306__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4990__ (
    .D(__2843__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1307__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4991__ (
    .D(__3173__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1308__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4992__ (
    .D(__2122__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1309__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4993__ (
    .D(__2753__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1310__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4994__ (
    .D(__3085__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1311__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4995__ (
    .D(__3218__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1312__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4996__ (
    .D(__2464__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1313__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4997__ (
    .D(__2594__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1314__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4998__ (
    .D(__2842__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1315__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4999__ (
    .D(__3317__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1316__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5000__ (
    .D(__2523__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1317__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5001__ (
    .D(__2916__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1318__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5002__ (
    .D(__3508__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1319__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5003__ (
    .D(__2305__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1320__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5004__ (
    .D(__2268__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1321__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5005__ (
    .D(__2977__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1322__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5006__ (
    .D(__3193__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1323__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5007__ (
    .D(__2460__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1324__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5008__ (
    .D(__2927__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1325__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5009__ (
    .D(__2912__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1326__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5010__ (
    .D(__3183__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1327__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5011__ (
    .D(__2623__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1328__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5012__ (
    .D(__2054__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1329__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5013__ (
    .D(__2759__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1330__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5014__ (
    .D(__2692__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1331__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5015__ (
    .D(__3127__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1332__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5016__ (
    .D(__2298__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1333__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5017__ (
    .D(__2297__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1334__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5018__ (
    .D(__3418__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1335__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5019__ (
    .D(__3163__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1336__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5020__ (
    .D(__3384__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1337__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5021__ (
    .D(__3386__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1338__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5022__ (
    .D(__2130__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1339__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5023__ (
    .D(__3633__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1340__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5024__ (
    .D(__3248__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1341__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5025__ (
    .D(__1619__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1342__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5026__ (
    .D(__3677__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1343__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5027__ (
    .D(__3498__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1344__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5028__ (
    .D(__3243__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1345__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5029__ (
    .D(__3381__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1346__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5030__ (
    .D(__3452__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1347__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5031__ (
    .D(__3444__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1348__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5032__ (
    .D(__70__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1349__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5033__ (
    .D(__3275__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1350__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5034__ (
    .D(__2961__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1351__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5035__ (
    .D(__3337__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1352__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5036__ (
    .D(__2769__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1353__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5037__ (
    .D(__69__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1354__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5038__ (
    .D(__2769__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1355__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5039__ (
    .D(__68__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1356__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5040__ (
    .D(__3408__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1357__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5041__ (
    .D(__2706__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1358__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5042__ (
    .D(__2267__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1359__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5043__ (
    .D(__2573__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1360__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5044__ (
    .D(__2859__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1361__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5045__ (
    .D(__3597__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1362__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5046__ (
    .D(__2522__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1363__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5047__ (
    .D(__2738__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1364__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5048__ (
    .D(__3507__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1365__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5049__ (
    .D(__3521__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1366__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5050__ (
    .D(__2409__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1367__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5051__ (
    .D(__2540__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1368__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5052__ (
    .D(__2965__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1369__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5053__ (
    .D(__3366__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1370__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5054__ (
    .D(__2931__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1371__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5055__ (
    .D(__3577__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1372__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5056__ (
    .D(__2610__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1373__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5057__ (
    .D(__3654__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1374__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5058__ (
    .D(__3043__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1375__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5059__ (
    .D(__3651__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1376__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5060__ (
    .D(__3034__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1377__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5061__ (
    .D(__2500__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1378__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5062__ (
    .D(__2915__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1379__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5063__ (
    .D(__3285__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1380__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5064__ (
    .D(__3373__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1381__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5065__ (
    .D(__3658__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1382__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5066__ (
    .D(__2801__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1383__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5067__ (
    .D(__2795__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1384__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5068__ (
    .D(__3149__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1385__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5069__ (
    .D(__3565__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1386__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5070__ (
    .D(__1629__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1387__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5071__ (
    .D(__3489__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1388__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5072__ (
    .D(__3620__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1389__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5073__ (
    .D(__1670__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1390__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5074__ (
    .D(__3456__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1391__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5075__ (
    .D(__3191__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1392__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5076__ (
    .D(__2092__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1393__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5077__ (
    .D(__3588__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1394__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5078__ (
    .D(__3596__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1395__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5079__ (
    .D(__2461__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1396__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5080__ (
    .D(__3438__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1397__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5081__ (
    .D(__2873__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1398__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5082__ (
    .D(__2883__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1399__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5083__ (
    .D(__2322__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1400__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5084__ (
    .D(__2203__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1401__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5085__ (
    .D(__3216__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1402__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5086__ (
    .D(__3174__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1403__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5087__ (
    .D(__2214__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1404__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5088__ (
    .D(__3091__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1405__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5089__ (
    .D(__3118__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1406__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5090__ (
    .D(__3188__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1407__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5091__ (
    .D(__3659__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1408__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5092__ (
    .D(__2832__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1409__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5093__ (
    .D(__3470__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1410__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5094__ (
    .D(__3307__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1411__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5095__ (
    .D(__2994__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1412__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5096__ (
    .D(__2981__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1413__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5097__ (
    .D(__3669__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1414__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5098__ (
    .D(__1416__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1415__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5099__ (
    .D(__3306__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1416__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5100__ (
    .D(__1418__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1417__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5101__ (
    .D(__2435__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1418__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5102__ (
    .D(__1420__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1419__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5103__ (
    .D(__3010__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1420__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5104__ (
    .D(__2860__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1421__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5105__ (
    .D(__1423__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1422__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5106__ (
    .D(__2026__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1423__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5107__ (
    .D(__1425__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1424__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5108__ (
    .D(__2309__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1425__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5109__ (
    .D(__1427__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1426__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5110__ (
    .D(__2132__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1427__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5111__ (
    .D(__1429__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1428__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5112__ (
    .D(__3657__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1429__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5113__ (
    .D(__1431__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1430__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5114__ (
    .D(__2838__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1431__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5115__ (
    .D(__1433__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1432__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5116__ (
    .D(__3018__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1433__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5117__ (
    .D(__1435__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1434__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5118__ (
    .D(__2831__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1435__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5119__ (
    .D(__1437__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1436__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5120__ (
    .D(__2543__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1437__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5121__ (
    .D(__1439__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1438__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5122__ (
    .D(__2360__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1439__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5123__ (
    .D(__1441__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1440__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5124__ (
    .D(__3115__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1441__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5125__ (
    .D(__1443__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1442__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5126__ (
    .D(__1867__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1443__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5127__ (
    .D(__1445__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1444__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5128__ (
    .D(__2972__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1445__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5129__ (
    .D(__1447__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1446__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5130__ (
    .D(__3398__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1447__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5131__ (
    .D(__1449__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1448__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5132__ (
    .D(__2353__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1449__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5133__ (
    .D(__1451__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1450__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5134__ (
    .D(__2929__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1451__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5135__ (
    .D(__3090__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1452__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5136__ (
    .D(__2684__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1453__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5137__ (
    .D(__2159__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1454__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5138__ (
    .D(__3491__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1455__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5139__ (
    .D(__2436__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1456__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5140__ (
    .D(__2153__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1457__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5141__ (
    .D(__2359__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1458__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5142__ (
    .D(__3445__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1459__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5143__ (
    .D(__3283__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1460__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5144__ (
    .D(g3213),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1461__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5145__ (
    .D(g3214),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1462__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5146__ (
    .D(g3215),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1463__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5147__ (
    .D(g3216),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1464__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5148__ (
    .D(g3217),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1465__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5149__ (
    .D(g3218),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1466__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5150__ (
    .D(g3219),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1467__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5151__ (
    .D(g3220),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1468__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5152__ (
    .D(g3232),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1469__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5153__ (
    .D(g3221),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1470__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5154__ (
    .D(g3222),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1471__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5155__ (
    .D(g3223),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1472__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5156__ (
    .D(g3224),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1473__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5157__ (
    .D(g3225),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1474__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5158__ (
    .D(g3226),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1475__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5159__ (
    .D(g3227),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1476__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5160__ (
    .D(g3228),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1477__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5161__ (
    .D(g3212),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1478__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5162__ (
    .D(__1780__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1479__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5163__ (
    .D(__1497__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1480__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5164__ (
    .D(__3341__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1481__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5165__ (
    .D(__3198__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1482__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5166__ (
    .D(__3342__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1483__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5167__ (
    .D(__2318__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1484__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5168__ (
    .D(__2431__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1485__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5169__ (
    .D(__3612__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1486__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5170__ (
    .D(__1612__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1487__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5171__ (
    .D(__2921__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1488__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5172__ (
    .D(__2736__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1489__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5173__ (
    .D(__2499__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1490__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5174__ (
    .D(__2146__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1491__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5175__ (
    .D(__2737__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1492__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5176__ (
    .D(__3055__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1493__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5177__ (
    .D(__3235__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1494__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5178__ (
    .D(__3482__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1495__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5179__ (
    .D(__2682__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1496__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5180__ (
    .D(g51),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1497__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5181__ (
    .D(__3303__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1498__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5182__ (
    .D(__2337__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1499__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5183__ (
    .D(__3324__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1500__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5184__ (
    .D(__2470__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1501__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5185__ (
    .D(__3143__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1502__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5186__ (
    .D(__2908__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1503__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5187__ (
    .D(__2658__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1504__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5188__ (
    .D(__3352__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1505__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5189__ (
    .D(__3140__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1506__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5190__ (
    .D(__3420__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1507__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5191__ (
    .D(__3067__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1508__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5192__ (
    .D(g3234),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1509__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5193__ (
    .D(__1509__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1510__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5194__ (
    .D(__2584__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1511__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5195__ (
    .D(__2402__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1512__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5196__ (
    .D(__2131__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1513__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5197__ (
    .D(__3364__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1514__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5198__ (
    .D(__1804__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1515__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5199__ (
    .D(__3469__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1516__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5200__ (
    .D(__2612__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1517__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5201__ (
    .D(__2158__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1518__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5202__ (
    .D(__3667__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1519__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5203__ (
    .D(__3635__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1520__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5204__ (
    .D(__3247__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1521__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5205__ (
    .D(__2336__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1522__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5206__ (
    .D(__2827__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1523__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5207__ (
    .D(__2216__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1524__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5208__ (
    .D(__2919__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1525__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5209__ (
    .D(__2874__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1526__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5210__ (
    .D(__2626__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1527__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5211__ (
    .D(__2779__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1528__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5212__ (
    .D(__2593__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1529__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5213__ (
    .D(__1662__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1530__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5214__ (
    .D(__1621__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1531__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5215__ (
    .D(__3346__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1532__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5216__ (
    .D(__3178__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1533__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5219__ (
    .I5(__589__),
    .I4(__1241__),
    .I3(__663__),
    .I2(__1244__),
    .I1(__662__),
    .I0(__1242__),
    .O(__1536__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5220__ (
    .I5(__589__),
    .I4(__1257__),
    .I3(__663__),
    .I2(__1267__),
    .I1(__662__),
    .I0(__1265__),
    .O(__1537__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5221__ (
    .I5(__589__),
    .I4(__1271__),
    .I3(__663__),
    .I2(__1273__),
    .I1(__662__),
    .I0(__1272__),
    .O(__1538__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5222__ (
    .I5(__589__),
    .I4(__1268__),
    .I3(__663__),
    .I2(__1270__),
    .I1(__662__),
    .I0(__1269__),
    .O(__1539__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5223__ (
    .I5(__589__),
    .I4(__1238__),
    .I3(__663__),
    .I2(__1240__),
    .I1(__662__),
    .I0(__1239__),
    .O(__1540__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __5224__ (
    .I1(__1540__),
    .I0(__1539__),
    .O(__1541__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5225__ (
    .I5(__589__),
    .I4(__1158__),
    .I3(__663__),
    .I2(__1162__),
    .I1(__662__),
    .I0(__1159__),
    .O(__1542__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5226__ (
    .I5(__589__),
    .I4(__1168__),
    .I3(__663__),
    .I2(__1170__),
    .I1(__662__),
    .I0(__1169__),
    .O(__1543__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5227__ (
    .I5(__589__),
    .I4(__1163__),
    .I3(__663__),
    .I2(__1167__),
    .I1(__662__),
    .I0(__1166__),
    .O(__1544__)
  );
  LUT3 #(
    .INIT(8'h08)
  ) __5228__ (
    .I2(__1544__),
    .I1(__1543__),
    .I0(__1542__),
    .O(__1545__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5229__ (
    .I5(__589__),
    .I4(__1274__),
    .I3(__663__),
    .I2(__1276__),
    .I1(__662__),
    .I0(__1275__),
    .O(__1546__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5230__ (
    .I5(__589__),
    .I4(__1254__),
    .I3(__663__),
    .I2(__1256__),
    .I1(__662__),
    .I0(__1255__),
    .O(__1547__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5231__ (
    .I5(__589__),
    .I4(__1248__),
    .I3(__663__),
    .I2(__1250__),
    .I1(__662__),
    .I0(__1249__),
    .O(__1548__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5232__ (
    .I5(__589__),
    .I4(__1251__),
    .I3(__663__),
    .I2(__1253__),
    .I1(__662__),
    .I0(__1252__),
    .O(__1549__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5233__ (
    .I5(__589__),
    .I4(__1245__),
    .I3(__663__),
    .I2(__1247__),
    .I1(__662__),
    .I0(__1246__),
    .O(__1550__)
  );
  LUT5 #(
    .INIT(32'h80000000)
  ) __5234__ (
    .I4(__1550__),
    .I3(__1549__),
    .I2(__1548__),
    .I1(__1547__),
    .I0(__1546__),
    .O(__1551__)
  );
  LUT6 #(
    .INIT(64'h0100000000000000)
  ) __5235__ (
    .I5(__1551__),
    .I4(__1545__),
    .I3(__1541__),
    .I2(__1538__),
    .I1(__1537__),
    .I0(__1536__),
    .O(__1552__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5236__ (
    .I1(__1538__),
    .I0(__1537__),
    .O(__1553__)
  );
  LUT6 #(
    .INIT(64'h4000000000000000)
  ) __5237__ (
    .I5(__1540__),
    .I4(__1539__),
    .I3(__1536__),
    .I2(__1551__),
    .I1(__1553__),
    .I0(__1545__),
    .O(__1554__)
  );
  LUT4 #(
    .INIT(16'he000)
  ) __5238__ (
    .I3(__1543__),
    .I2(__1542__),
    .I1(__1554__),
    .I0(__1552__),
    .O(__1555__)
  );
  LUT6 #(
    .INIT(64'h8000010000000000)
  ) __5239__ (
    .I5(__1543__),
    .I4(__1544__),
    .I3(__1542__),
    .I2(__1538__),
    .I1(__1539__),
    .I0(__1546__),
    .O(__1556__)
  );
  LUT6 #(
    .INIT(64'h9393399393939393)
  ) __5240__ (
    .I5(__1543__),
    .I4(__1544__),
    .I3(__1542__),
    .I2(__1537__),
    .I1(__1547__),
    .I0(__1556__),
    .O(__1557__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5241__ (
    .I5(__589__),
    .I4(__1295__),
    .I3(__663__),
    .I2(__1297__),
    .I1(__662__),
    .I0(__1296__),
    .O(__1558__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5242__ (
    .I5(__589__),
    .I4(__1302__),
    .I3(__663__),
    .I2(__1305__),
    .I1(__662__),
    .I0(__1303__),
    .O(__1559__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5243__ (
    .I5(__589__),
    .I4(__1334__),
    .I3(__663__),
    .I2(__1342__),
    .I1(__662__),
    .I0(__1341__),
    .O(__1560__)
  );
  LUT6 #(
    .INIT(64'h0000066006600000)
  ) __5244__ (
    .I5(__1417__),
    .I4(__1560__),
    .I3(__1428__),
    .I2(__1559__),
    .I1(__1432__),
    .I0(__1558__),
    .O(__1561__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5245__ (
    .I5(__589__),
    .I4(__1313__),
    .I3(__663__),
    .I2(__1315__),
    .I1(__662__),
    .I0(__1314__),
    .O(__1562__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5246__ (
    .I5(__589__),
    .I4(__1319__),
    .I3(__663__),
    .I2(__1321__),
    .I1(__662__),
    .I0(__1320__),
    .O(__1563__)
  );
  LUT4 #(
    .INIT(16'h1428)
  ) __5247__ (
    .I3(__1426__),
    .I2(__1422__),
    .I1(__1563__),
    .I0(__1562__),
    .O(__1564__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5248__ (
    .I5(__589__),
    .I4(__1280__),
    .I3(__663__),
    .I2(__1282__),
    .I1(__662__),
    .I0(__1281__),
    .O(__1565__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5249__ (
    .I5(__589__),
    .I4(__1292__),
    .I3(__663__),
    .I2(__1294__),
    .I1(__662__),
    .I0(__1293__),
    .O(__1566__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5250__ (
    .I5(__589__),
    .I4(__1316__),
    .I3(__663__),
    .I2(__1318__),
    .I1(__662__),
    .I0(__1317__),
    .O(__1567__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5251__ (
    .I5(__589__),
    .I4(__1298__),
    .I3(__663__),
    .I2(__1300__),
    .I1(__662__),
    .I0(__1299__),
    .O(__1568__)
  );
  LUT6 #(
    .INIT(64'h0000099009900000)
  ) __5252__ (
    .I5(__1430__),
    .I4(__1568__),
    .I3(__1424__),
    .I2(__1567__),
    .I1(__1566__),
    .I0(__1565__),
    .O(__1569__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5253__ (
    .I5(__589__),
    .I4(__1286__),
    .I3(__663__),
    .I2(__1288__),
    .I1(__662__),
    .I0(__1287__),
    .O(__1570__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5254__ (
    .I5(__589__),
    .I4(__1289__),
    .I3(__663__),
    .I2(__1291__),
    .I1(__662__),
    .I0(__1290__),
    .O(__1571__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5255__ (
    .I5(__589__),
    .I4(__1283__),
    .I3(__663__),
    .I2(__1285__),
    .I1(__662__),
    .I0(__1284__),
    .O(__1572__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5256__ (
    .I5(__589__),
    .I4(__1322__),
    .I3(__663__),
    .I2(__1329__),
    .I1(__662__),
    .I0(__1323__),
    .O(__1573__)
  );
  LUT6 #(
    .INIT(64'h0041410000000000)
  ) __5257__ (
    .I5(__603__),
    .I4(__1419__),
    .I3(__1573__),
    .I2(__1572__),
    .I1(__1571__),
    .I0(__1570__),
    .O(__1574__)
  );
  LUT4 #(
    .INIT(16'h8000)
  ) __5258__ (
    .I3(__1574__),
    .I2(__1569__),
    .I1(__1564__),
    .I0(__1561__),
    .O(__1575__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __5259__ (
    .I1(__1417__),
    .I0(__1546__),
    .O(__1576__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __5260__ (
    .I1(__1426__),
    .I0(__1547__),
    .O(__1577__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __5261__ (
    .I1(__1430__),
    .I0(__1548__),
    .O(__1578__)
  );
  LUT2 #(
    .INIT(4'h9)
  ) __5262__ (
    .I1(__1565__),
    .I0(__1536__),
    .O(__1579__)
  );
  LUT6 #(
    .INIT(64'he880fee8fee8e880)
  ) __5263__ (
    .I5(__1422__),
    .I4(__1539__),
    .I3(__1579__),
    .I2(__1578__),
    .I1(__1577__),
    .I0(__1576__),
    .O(__1580__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __5264__ (
    .I1(__1428__),
    .I0(__1549__),
    .O(__1581__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __5265__ (
    .I1(__1432__),
    .I0(__1550__),
    .O(__1582__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __5266__ (
    .I1(__1572__),
    .I0(__1540__),
    .O(__1583__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __5267__ (
    .I1(__1424__),
    .I0(__1537__),
    .O(__1584__)
  );
  LUT6 #(
    .INIT(64'h8e08ef8eef8e8e08)
  ) __5268__ (
    .I5(__1419__),
    .I4(__1538__),
    .I3(__1584__),
    .I2(__1583__),
    .I1(__1582__),
    .I0(__1581__),
    .O(__1585__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5269__ (
    .I1(__1544__),
    .I0(__1542__),
    .O(__1586__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5270__ (
    .I5(__589__),
    .I4(__1155__),
    .I3(__663__),
    .I2(__1157__),
    .I1(__662__),
    .I0(__1156__),
    .O(__1587__)
  );
  LUT6 #(
    .INIT(64'h0000000000008000)
  ) __5271__ (
    .I5(__1543__),
    .I4(__1587__),
    .I3(__1586__),
    .I2(__1585__),
    .I1(__1580__),
    .I0(__1575__),
    .O(__1588__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5272__ (
    .I1(__1544__),
    .I0(__1542__),
    .O(__1589__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5273__ (
    .I1(__603__),
    .I0(__1570__),
    .O(__1590__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5274__ (
    .I5(__589__),
    .I4(__1152__),
    .I3(__663__),
    .I2(__1154__),
    .I1(__662__),
    .I0(__1153__),
    .O(__1591__)
  );
  LUT6 #(
    .INIT(64'hff00ffff0b000f0f)
  ) __5275__ (
    .I5(__1543__),
    .I4(__1575__),
    .I3(__1591__),
    .I2(__1590__),
    .I1(__1589__),
    .I0(__1587__),
    .O(__1592__)
  );
  LUT5 #(
    .INIT(32'h0fbb0f0f)
  ) __5276__ (
    .I4(__1592__),
    .I3(__1588__),
    .I2(__1426__),
    .I1(__1557__),
    .I0(__1555__),
    .O(__1593__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __5277__ (
    .I2(__662__),
    .I1(__1593__),
    .I0(__1255__),
    .O(__1594__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5278__ (
    .I5(__589__),
    .I4(__1081__),
    .I3(__663__),
    .I2(__1084__),
    .I1(__662__),
    .I0(__1083__),
    .O(__1595__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5279__ (
    .I5(__589__),
    .I4(__1086__),
    .I3(__663__),
    .I2(__743__),
    .I1(__662__),
    .I0(__1088__),
    .O(__1596__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5280__ (
    .I5(__589__),
    .I4(__850__),
    .I3(__663__),
    .I2(__791__),
    .I1(__662__),
    .I0(__787__),
    .O(__1597__)
  );
  LUT5 #(
    .INIT(32'h00000001)
  ) __5281__ (
    .I4(__1487__),
    .I3(__1488__),
    .I2(__1489__),
    .I1(__1490__),
    .I0(__1491__),
    .O(__1598__)
  );
  LUT5 #(
    .INIT(32'h80ef0000)
  ) __5282__ (
    .I4(__589__),
    .I3(__1598__),
    .I2(__1597__),
    .I1(__1596__),
    .I0(__1595__),
    .O(__1599__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5283__ (
    .I5(__589__),
    .I4(__1135__),
    .I3(__663__),
    .I2(__1137__),
    .I1(__662__),
    .I0(__1136__),
    .O(__1600__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5284__ (
    .I5(__589__),
    .I4(__1132__),
    .I3(__663__),
    .I2(__1134__),
    .I1(__662__),
    .I0(__1133__),
    .O(__1601__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5285__ (
    .I5(__589__),
    .I4(__1138__),
    .I3(__663__),
    .I2(__1139__),
    .I1(__662__),
    .I0(__1114__),
    .O(__1602__)
  );
  LUT6 #(
    .INIT(64'hd8fad850d850d8fa)
  ) __5286__ (
    .I5(g3229),
    .I4(__1602__),
    .I3(__1601__),
    .I2(__1135__),
    .I1(__1600__),
    .I0(__1599__),
    .O(__1603__)
  );
  LUT5 #(
    .INIT(32'h0030aaaa)
  ) __5287__ (
    .I4(__662__),
    .I3(__1596__),
    .I2(__1597__),
    .I1(__1595__),
    .I0(__442__),
    .O(__1604__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5288__ (
    .I5(__944__),
    .I4(__447__),
    .I3(__858__),
    .I2(__438__),
    .I1(__954__),
    .I0(__431__),
    .O(__1605__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5289__ (
    .I5(__589__),
    .I4(__523__),
    .I3(__663__),
    .I2(__525__),
    .I1(__662__),
    .I0(__524__),
    .O(__1606__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __5290__ (
    .I2(__662__),
    .I1(__1606__),
    .I0(__200__),
    .O(__1607__)
  );
  LUT5 #(
    .INIT(32'h80000000)
  ) __5291__ (
    .I4(__1490__),
    .I3(__1491__),
    .I2(__1493__),
    .I1(__1492__),
    .I0(__1494__),
    .O(__1608__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5292__ (
    .I1(__1492__),
    .I0(__1491__),
    .O(__1609__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5293__ (
    .I1(__1494__),
    .I0(__1493__),
    .O(__1610__)
  );
  LUT6 #(
    .INIT(64'h4000000000000000)
  ) __5294__ (
    .I5(__1487__),
    .I4(__1489__),
    .I3(__1490__),
    .I2(__1610__),
    .I1(__1609__),
    .I0(__1488__),
    .O(__1611__)
  );
  LUT6 #(
    .INIT(64'h00000000007f0080)
  ) __5295__ (
    .I5(__1497__),
    .I4(__1487__),
    .I3(__1611__),
    .I2(__1488__),
    .I1(__1489__),
    .I0(__1608__),
    .O(__1612__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5296__ (
    .I5(__589__),
    .I4(__1102__),
    .I3(__663__),
    .I2(__1107__),
    .I1(__662__),
    .I0(__1106__),
    .O(__1613__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5297__ (
    .I5(__589__),
    .I4(__1227__),
    .I3(__663__),
    .I2(__1262__),
    .I1(__662__),
    .I0(__1261__),
    .O(__1614__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5298__ (
    .I1(__1460__),
    .I0(__1457__),
    .O(__1615__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5299__ (
    .I1(__1455__),
    .I0(__1456__),
    .O(__1616__)
  );
  LUT6 #(
    .INIT(64'h8000000000000000)
  ) __5300__ (
    .I5(__1453__),
    .I4(__1458__),
    .I3(__1459__),
    .I2(__1454__),
    .I1(__1616__),
    .I0(__1615__),
    .O(__1617__)
  );
  LUT6 #(
    .INIT(64'h0f005555cccccccc)
  ) __5301__ (
    .I5(__589__),
    .I4(__603__),
    .I3(__1617__),
    .I2(__1614__),
    .I1(__1102__),
    .I0(__1613__),
    .O(__1618__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __5302__ (
    .I3(__663__),
    .I2(__603__),
    .I1(__1417__),
    .I0(__1342__),
    .O(__1619__)
  );
  LUT5 #(
    .INIT(32'h0030aaaa)
  ) __5303__ (
    .I4(__589__),
    .I3(__1597__),
    .I2(__1596__),
    .I1(__1595__),
    .I0(__416__),
    .O(__1620__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __5304__ (
    .I2(__1511__),
    .I1(__119__),
    .I0(__78__),
    .O(__1621__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5305__ (
    .I1(__1504__),
    .I0(__1501__),
    .O(__1622__)
  );
  LUT6 #(
    .INIT(64'h0100000000000000)
  ) __5306__ (
    .I5(__1622__),
    .I4(__1502__),
    .I3(__1499__),
    .I2(__1503__),
    .I1(__1500__),
    .I0(__1498__),
    .O(__1623__)
  );
  LUT5 #(
    .INIT(32'h00000080)
  ) __5307__ (
    .I4(__1508__),
    .I3(__1507__),
    .I2(__1623__),
    .I1(__1506__),
    .I0(__1505__),
    .O(__1624__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5308__ (
    .I5(__246__),
    .I4(__858__),
    .I3(__944__),
    .I2(__223__),
    .I1(__237__),
    .I0(__954__),
    .O(__1625__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5309__ (
    .I1(__954__),
    .I0(__114__),
    .O(__1626__)
  );
  LUT6 #(
    .INIT(64'h0000000000bfbfbf)
  ) __5310__ (
    .I5(__1626__),
    .I4(__944__),
    .I3(__113__),
    .I2(__1347__),
    .I1(__167__),
    .I0(__1625__),
    .O(__1627__)
  );
  LUT6 #(
    .INIT(64'h4545ff000505ff00)
  ) __5311__ (
    .I5(__858__),
    .I4(__954__),
    .I3(__114__),
    .I2(__1627__),
    .I1(__115__),
    .I0(__1624__),
    .O(__1628__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __5312__ (
    .I2(__858__),
    .I1(__867__),
    .I0(__1387__),
    .O(__1629__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __5313__ (
    .I2(__944__),
    .I1(__266__),
    .I0(__875__),
    .O(__1630__)
  );
  LUT5 #(
    .INIT(32'h0030aaaa)
  ) __5314__ (
    .I4(__663__),
    .I3(__1597__),
    .I2(__1596__),
    .I1(__1595__),
    .I0(__423__),
    .O(__1631__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5315__ (
    .I5(__589__),
    .I4(__1129__),
    .I3(__663__),
    .I2(__1131__),
    .I1(__662__),
    .I0(__1130__),
    .O(__1632__)
  );
  LUT5 #(
    .INIT(32'h80ef0000)
  ) __5316__ (
    .I4(__662__),
    .I3(__1598__),
    .I2(__1597__),
    .I1(__1596__),
    .I0(__1595__),
    .O(__1633__)
  );
  LUT6 #(
    .INIT(64'hcc77f0f077ccf0f0)
  ) __5317__ (
    .I5(g3229),
    .I4(__1633__),
    .I3(__1602__),
    .I2(__1133__),
    .I1(__1600__),
    .I0(__1632__),
    .O(__1634__)
  );
  LUT6 #(
    .INIT(64'h0000000000000008)
  ) __5318__ (
    .I5(__1492__),
    .I4(__1483__),
    .I3(__1485__),
    .I2(__1486__),
    .I1(__1484__),
    .I0(__1493__),
    .O(__1635__)
  );
  LUT5 #(
    .INIT(32'h4ecccccc)
  ) __5319__ (
    .I4(__663__),
    .I3(__1598__),
    .I2(__1408__),
    .I1(__448__),
    .I0(__1635__),
    .O(__1636__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5320__ (
    .I5(__589__),
    .I4(__1277__),
    .I3(__663__),
    .I2(__1279__),
    .I1(__662__),
    .I0(__1278__),
    .O(__1637__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5321__ (
    .I5(__589__),
    .I4(__1184__),
    .I3(__663__),
    .I2(__1186__),
    .I1(__662__),
    .I0(__1185__),
    .O(__1638__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5322__ (
    .I5(__589__),
    .I4(__1171__),
    .I3(__663__),
    .I2(__1177__),
    .I1(__662__),
    .I0(__1172__),
    .O(__1639__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5323__ (
    .I5(__589__),
    .I4(__1179__),
    .I3(__663__),
    .I2(__1183__),
    .I1(__662__),
    .I0(__1181__),
    .O(__1640__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5324__ (
    .I1(__1424__),
    .I0(__1422__),
    .O(__1641__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5325__ (
    .I1(__1426__),
    .I0(__1432__),
    .O(__1642__)
  );
  LUT6 #(
    .INIT(64'h8000000000000000)
  ) __5326__ (
    .I5(__1419__),
    .I4(__1430__),
    .I3(__1417__),
    .I2(__1428__),
    .I1(__1642__),
    .I0(__1641__),
    .O(__1643__)
  );
  LUT6 #(
    .INIT(64'h01f700f300ff00ff)
  ) __5327__ (
    .I5(__603__),
    .I4(__1643__),
    .I3(__1640__),
    .I2(__1639__),
    .I1(__1638__),
    .I0(__1637__),
    .O(__1644__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __5328__ (
    .I2(__663__),
    .I1(__1644__),
    .I0(__1183__),
    .O(__1645__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5329__ (
    .I5(__944__),
    .I4(__807__),
    .I3(__858__),
    .I2(__809__),
    .I1(__954__),
    .I0(__808__),
    .O(__1646__)
  );
  LUT5 #(
    .INIT(32'h00000001)
  ) __5330__ (
    .I4(__1504__),
    .I3(__1501__),
    .I2(__1502__),
    .I1(__1503__),
    .I0(__1500__),
    .O(__1647__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5331__ (
    .I5(__944__),
    .I4(__853__),
    .I3(__858__),
    .I2(__574__),
    .I1(__954__),
    .I0(__803__),
    .O(__1648__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5332__ (
    .I5(__944__),
    .I4(__804__),
    .I3(__858__),
    .I2(__806__),
    .I1(__954__),
    .I0(__805__),
    .O(__1649__)
  );
  LUT6 #(
    .INIT(64'h4f0f4f0000000000)
  ) __5333__ (
    .I5(__944__),
    .I4(__1649__),
    .I3(__1648__),
    .I2(__1647__),
    .I1(__968__),
    .I0(__1646__),
    .O(__1650__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5334__ (
    .I5(__944__),
    .I4(__564__),
    .I3(__858__),
    .I2(__821__),
    .I1(__954__),
    .I0(__863__),
    .O(__1651__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5335__ (
    .I5(__944__),
    .I4(__864__),
    .I3(__858__),
    .I2(__825__),
    .I1(__954__),
    .I0(__865__),
    .O(__1652__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5336__ (
    .I5(__944__),
    .I4(__577__),
    .I3(__858__),
    .I2(__866__),
    .I1(__954__),
    .I0(__859__),
    .O(__1653__)
  );
  LUT6 #(
    .INIT(64'h4eeeeeeeeeee4eee)
  ) __5337__ (
    .I5(g3229),
    .I4(__1653__),
    .I3(__1652__),
    .I2(__1651__),
    .I1(__816__),
    .I0(__1650__),
    .O(__1654__)
  );
  LUT5 #(
    .INIT(32'h81000000)
  ) __5338__ (
    .I4(__1543__),
    .I3(__1542__),
    .I2(__1544__),
    .I1(__1538__),
    .I0(__1546__),
    .O(__1655__)
  );
  LUT6 #(
    .INIT(64'h4000000200000000)
  ) __5339__ (
    .I5(__1655__),
    .I4(__1537__),
    .I3(__1549__),
    .I2(__1539__),
    .I1(__1547__),
    .I0(__1545__),
    .O(__1656__)
  );
  LUT6 #(
    .INIT(64'h5555cffc55555555)
  ) __5340__ (
    .I5(__1592__),
    .I4(__1588__),
    .I3(__1548__),
    .I2(__1656__),
    .I1(__1555__),
    .I0(__1430__),
    .O(__1657__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __5341__ (
    .I2(__663__),
    .I1(__1657__),
    .I0(__1250__),
    .O(__1658__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __5342__ (
    .I2(__944__),
    .I1(__969__),
    .I0(__968__),
    .O(__1659__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __5343__ (
    .I5(__858__),
    .I4(__242__),
    .I3(__370__),
    .I2(__229__),
    .I1(__169__),
    .I0(__220__),
    .O(__1660__)
  );
  LUT5 #(
    .INIT(32'h0030aaaa)
  ) __5344__ (
    .I4(__662__),
    .I3(__1544__),
    .I2(__1543__),
    .I1(__1542__),
    .I0(__1006__),
    .O(__1661__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __5345__ (
    .I2(__1511__),
    .I1(__79__),
    .I0(__102__),
    .O(__1662__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5346__ (
    .I5(__858__),
    .I4(__958__),
    .I3(__944__),
    .I2(__922__),
    .I1(__954__),
    .I0(__412__),
    .O(__1663__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5347__ (
    .I1(__954__),
    .I0(__811__),
    .O(__1664__)
  );
  LUT6 #(
    .INIT(64'h0000000000bfbfbf)
  ) __5348__ (
    .I5(__1664__),
    .I4(__944__),
    .I3(__810__),
    .I2(__1347__),
    .I1(__465__),
    .I0(__1663__),
    .O(__1665__)
  );
  LUT6 #(
    .INIT(64'h4545ff000505ff00)
  ) __5349__ (
    .I5(__858__),
    .I4(__954__),
    .I3(__811__),
    .I2(__1665__),
    .I1(__812__),
    .I0(__1624__),
    .O(__1666__)
  );
  LUT6 #(
    .INIT(64'h4000000000000000)
  ) __5350__ (
    .I5(__944__),
    .I4(__799__),
    .I3(__747__),
    .I2(__1051__),
    .I1(__802__),
    .I0(__748__),
    .O(__1667__)
  );
  LUT4 #(
    .INIT(16'h8000)
  ) __5351__ (
    .I3(__1055__),
    .I2(__788__),
    .I1(__796__),
    .I0(__1667__),
    .O(__1668__)
  );
  LUT5 #(
    .INIT(32'h12305af0)
  ) __5352__ (
    .I4(__954__),
    .I3(__737__),
    .I2(__1047__),
    .I1(__875__),
    .I0(__1668__),
    .O(__1669__)
  );
  LUT6 #(
    .INIT(64'haa3aaaaaaaaaaaaa)
  ) __5353__ (
    .I5(__858__),
    .I4(__93__),
    .I3(__748__),
    .I2(__73__),
    .I1(__788__),
    .I0(__1390__),
    .O(__1670__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __5354__ (
    .I3(__589__),
    .I2(__603__),
    .I1(__1460__),
    .I0(__1049__),
    .O(__1671__)
  );
  LUT6 #(
    .INIT(64'hfffff888f888f888)
  ) __5355__ (
    .I5(__589__),
    .I4(__1190__),
    .I3(__663__),
    .I2(__1192__),
    .I1(__662__),
    .I0(__1191__),
    .O(__1672__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __5356__ (
    .I2(__589__),
    .I1(__1672__),
    .I0(__999__),
    .O(__1673__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5357__ (
    .I5(__944__),
    .I4(__943__),
    .I3(__858__),
    .I2(__946__),
    .I1(__954__),
    .I0(__945__),
    .O(__1674__)
  );
  LUT4 #(
    .INIT(16'haccc)
  ) __5358__ (
    .I3(__858__),
    .I2(__925__),
    .I1(__877__),
    .I0(__1674__),
    .O(__1675__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __5359__ (
    .I5(__954__),
    .I4(__936__),
    .I3(__927__),
    .I2(__924__),
    .I1(__903__),
    .I0(__918__),
    .O(__1676__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5360__ (
    .I5(__589__),
    .I4(__617__),
    .I3(__663__),
    .I2(__618__),
    .I1(__662__),
    .I0(__441__),
    .O(__1677__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5361__ (
    .I5(__589__),
    .I4(__614__),
    .I3(__663__),
    .I2(__455__),
    .I1(__662__),
    .I0(__454__),
    .O(__1678__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5362__ (
    .I5(__589__),
    .I4(__452__),
    .I3(__663__),
    .I2(__616__),
    .I1(__662__),
    .I0(__520__),
    .O(__1679__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5363__ (
    .I5(__589__),
    .I4(__451__),
    .I3(__663__),
    .I2(__457__),
    .I1(__662__),
    .I0(__355__),
    .O(__1680__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5364__ (
    .I5(__589__),
    .I4(__583__),
    .I3(__663__),
    .I2(__160__),
    .I1(__662__),
    .I0(__159__),
    .O(__1681__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5365__ (
    .I5(__589__),
    .I4(__161__),
    .I3(__663__),
    .I2(__543__),
    .I1(__662__),
    .I0(__460__),
    .O(__1682__)
  );
  LUT6 #(
    .INIT(64'h9333363333333333)
  ) __5366__ (
    .I5(__1682__),
    .I4(__1681__),
    .I3(__1680__),
    .I2(__1679__),
    .I1(__1678__),
    .I0(__1677__),
    .O(__1683__)
  );
  LUT3 #(
    .INIT(8'h08)
  ) __5367__ (
    .I2(__1681__),
    .I1(__1682__),
    .I0(__1680__),
    .O(__1684__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5368__ (
    .I5(__589__),
    .I4(__439__),
    .I3(__663__),
    .I2(__609__),
    .I1(__662__),
    .I0(__516__),
    .O(__1685__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5369__ (
    .I5(__589__),
    .I4(__613__),
    .I3(__663__),
    .I2(__428__),
    .I1(__662__),
    .I0(__587__),
    .O(__1686__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5370__ (
    .I5(__589__),
    .I4(__582__),
    .I3(__663__),
    .I2(__444__),
    .I1(__662__),
    .I0(__572__),
    .O(__1687__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __5371__ (
    .I1(__1687__),
    .I0(__1678__),
    .O(__1688__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5372__ (
    .I5(__589__),
    .I4(__519__),
    .I3(__663__),
    .I2(__579__),
    .I1(__662__),
    .I0(__612__),
    .O(__1689__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5373__ (
    .I5(__589__),
    .I4(__576__),
    .I3(__663__),
    .I2(__611__),
    .I1(__662__),
    .I0(__517__),
    .O(__1690__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5374__ (
    .I5(__589__),
    .I4(__449__),
    .I3(__663__),
    .I2(__446__),
    .I1(__662__),
    .I0(__450__),
    .O(__1691__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5375__ (
    .I5(__589__),
    .I4(__575__),
    .I3(__663__),
    .I2(__584__),
    .I1(__662__),
    .I0(__610__),
    .O(__1692__)
  );
  LUT5 #(
    .INIT(32'h80000000)
  ) __5376__ (
    .I4(__1692__),
    .I3(__1691__),
    .I2(__1690__),
    .I1(__1689__),
    .I0(__1677__),
    .O(__1693__)
  );
  LUT6 #(
    .INIT(64'h0100000000000000)
  ) __5377__ (
    .I5(__1693__),
    .I4(__1684__),
    .I3(__1688__),
    .I2(__1679__),
    .I1(__1686__),
    .I0(__1685__),
    .O(__1694__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5378__ (
    .I1(__1679__),
    .I0(__1686__),
    .O(__1695__)
  );
  LUT6 #(
    .INIT(64'h4000000000000000)
  ) __5379__ (
    .I5(__1687__),
    .I4(__1678__),
    .I3(__1685__),
    .I2(__1693__),
    .I1(__1695__),
    .I0(__1684__),
    .O(__1696__)
  );
  LUT4 #(
    .INIT(16'he000)
  ) __5380__ (
    .I3(__1682__),
    .I2(__1680__),
    .I1(__1696__),
    .I0(__1694__),
    .O(__1697__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5381__ (
    .I5(__589__),
    .I4(__591__),
    .I3(__663__),
    .I2(__536__),
    .I1(__662__),
    .I0(__235__),
    .O(__1698__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5382__ (
    .I5(__589__),
    .I4(__340__),
    .I3(__663__),
    .I2(__638__),
    .I1(__662__),
    .I0(__344__),
    .O(__1699__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5383__ (
    .I5(__589__),
    .I4(__432__),
    .I3(__663__),
    .I2(__456__),
    .I1(__662__),
    .I0(__434__),
    .O(__1700__)
  );
  LUT6 #(
    .INIT(64'h0000066006600000)
  ) __5384__ (
    .I5(__1407__),
    .I4(__1700__),
    .I3(__1699__),
    .I2(__1412__),
    .I1(__1414__),
    .I0(__1698__),
    .O(__1701__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5385__ (
    .I5(__589__),
    .I4(__639__),
    .I3(__663__),
    .I2(__476__),
    .I1(__662__),
    .I0(__440__),
    .O(__1702__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5386__ (
    .I5(__589__),
    .I4(__471__),
    .I3(__663__),
    .I2(__538__),
    .I1(__662__),
    .I0(__485__),
    .O(__1703__)
  );
  LUT4 #(
    .INIT(16'h1428)
  ) __5387__ (
    .I3(__1411__),
    .I2(__1409__),
    .I1(__1703__),
    .I0(__1702__),
    .O(__1704__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5388__ (
    .I5(__589__),
    .I4(__622__),
    .I3(__663__),
    .I2(__623__),
    .I1(__662__),
    .I0(__437__),
    .O(__1705__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5389__ (
    .I5(__589__),
    .I4(__586__),
    .I3(__663__),
    .I2(__226__),
    .I1(__662__),
    .I0(__593__),
    .O(__1706__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5390__ (
    .I5(__589__),
    .I4(__665__),
    .I3(__663__),
    .I2(__655__),
    .I1(__662__),
    .I0(__453__),
    .O(__1707__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5391__ (
    .I5(__589__),
    .I4(__221__),
    .I3(__663__),
    .I2(__210__),
    .I1(__662__),
    .I0(__214__),
    .O(__1708__)
  );
  LUT6 #(
    .INIT(64'h0000099009900000)
  ) __5392__ (
    .I5(__1708__),
    .I4(__1413__),
    .I3(__1410__),
    .I2(__1707__),
    .I1(__1706__),
    .I0(__1705__),
    .O(__1709__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5393__ (
    .I5(__589__),
    .I4(__458__),
    .I3(__663__),
    .I2(__590__),
    .I1(__662__),
    .I0(__626__),
    .O(__1710__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5394__ (
    .I5(__589__),
    .I4(__374__),
    .I3(__663__),
    .I2(__376__),
    .I1(__662__),
    .I0(__592__),
    .O(__1711__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5395__ (
    .I5(__589__),
    .I4(__461__),
    .I3(__663__),
    .I2(__448__),
    .I1(__662__),
    .I0(__585__),
    .O(__1712__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5396__ (
    .I5(__589__),
    .I4(__425__),
    .I3(__663__),
    .I2(__430__),
    .I1(__662__),
    .I0(__427__),
    .O(__1713__)
  );
  LUT6 #(
    .INIT(64'h0041410000000000)
  ) __5397__ (
    .I5(__603__),
    .I4(__1408__),
    .I3(__1713__),
    .I2(__1712__),
    .I1(__1711__),
    .I0(__1710__),
    .O(__1714__)
  );
  LUT4 #(
    .INIT(16'h8000)
  ) __5398__ (
    .I3(__1714__),
    .I2(__1709__),
    .I1(__1704__),
    .I0(__1701__),
    .O(__1715__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __5399__ (
    .I1(__1407__),
    .I0(__1677__),
    .O(__1716__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __5400__ (
    .I1(__1411__),
    .I0(__1689__),
    .O(__1717__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __5401__ (
    .I1(__1413__),
    .I0(__1690__),
    .O(__1718__)
  );
  LUT2 #(
    .INIT(4'h9)
  ) __5402__ (
    .I1(__1705__),
    .I0(__1685__),
    .O(__1719__)
  );
  LUT6 #(
    .INIT(64'he880fee8fee8e880)
  ) __5403__ (
    .I5(__1409__),
    .I4(__1678__),
    .I3(__1719__),
    .I2(__1718__),
    .I1(__1717__),
    .I0(__1716__),
    .O(__1720__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __5404__ (
    .I1(__1412__),
    .I0(__1691__),
    .O(__1721__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __5405__ (
    .I1(__1414__),
    .I0(__1692__),
    .O(__1722__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __5406__ (
    .I1(__1712__),
    .I0(__1687__),
    .O(__1723__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __5407__ (
    .I1(__1410__),
    .I0(__1686__),
    .O(__1724__)
  );
  LUT6 #(
    .INIT(64'h8e08ef8eef8e8e08)
  ) __5408__ (
    .I5(__1408__),
    .I4(__1679__),
    .I3(__1724__),
    .I2(__1723__),
    .I1(__1722__),
    .I0(__1721__),
    .O(__1725__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5409__ (
    .I1(__1681__),
    .I0(__1680__),
    .O(__1726__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5410__ (
    .I5(__589__),
    .I4(__421__),
    .I3(__663__),
    .I2(__118__),
    .I1(__662__),
    .I0(__541__),
    .O(__1727__)
  );
  LUT6 #(
    .INIT(64'h0000000000008000)
  ) __5411__ (
    .I5(__1682__),
    .I4(__1727__),
    .I3(__1726__),
    .I2(__1725__),
    .I1(__1720__),
    .I0(__1715__),
    .O(__1728__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5412__ (
    .I1(__1681__),
    .I0(__1680__),
    .O(__1729__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5413__ (
    .I1(__603__),
    .I0(__1710__),
    .O(__1730__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5414__ (
    .I5(__589__),
    .I4(__467__),
    .I3(__663__),
    .I2(__533__),
    .I1(__662__),
    .I0(__470__),
    .O(__1731__)
  );
  LUT6 #(
    .INIT(64'hff00ffff0b000f0f)
  ) __5415__ (
    .I5(__1682__),
    .I4(__1715__),
    .I3(__1731__),
    .I2(__1730__),
    .I1(__1729__),
    .I0(__1727__),
    .O(__1732__)
  );
  LUT6 #(
    .INIT(64'hf0f033aaf0f0f0f0)
  ) __5416__ (
    .I5(__1732__),
    .I4(__1728__),
    .I3(__1697__),
    .I2(__1409__),
    .I1(__1684__),
    .I0(__1683__),
    .O(__1733__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __5417__ (
    .I2(__662__),
    .I1(__1733__),
    .I0(__454__),
    .O(__1734__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5418__ (
    .I5(__589__),
    .I4(__738__),
    .I3(__663__),
    .I2(__742__),
    .I1(__662__),
    .I0(__739__),
    .O(__1735__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __5419__ (
    .I1(__1436__),
    .I0(__1735__),
    .O(__1736__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5420__ (
    .I5(__589__),
    .I4(__714__),
    .I3(__663__),
    .I2(__716__),
    .I1(__662__),
    .I0(__715__),
    .O(__1737__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __5421__ (
    .I1(__1444__),
    .I0(__1737__),
    .O(__1738__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5422__ (
    .I5(__589__),
    .I4(__708__),
    .I3(__663__),
    .I2(__710__),
    .I1(__662__),
    .I0(__709__),
    .O(__1739__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __5423__ (
    .I1(__1448__),
    .I0(__1739__),
    .O(__1740__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5424__ (
    .I5(__589__),
    .I4(__687__),
    .I3(__663__),
    .I2(__699__),
    .I1(__662__),
    .I0(__695__),
    .O(__1741__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5425__ (
    .I5(__589__),
    .I4(__775__),
    .I3(__663__),
    .I2(__777__),
    .I1(__662__),
    .I0(__776__),
    .O(__1742__)
  );
  LUT2 #(
    .INIT(4'h9)
  ) __5426__ (
    .I1(__1742__),
    .I0(__1741__),
    .O(__1743__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5427__ (
    .I5(__589__),
    .I4(__720__),
    .I3(__663__),
    .I2(__722__),
    .I1(__662__),
    .I0(__721__),
    .O(__1744__)
  );
  LUT6 #(
    .INIT(64'he880fee8fee8e880)
  ) __5428__ (
    .I5(__1440__),
    .I4(__1744__),
    .I3(__1743__),
    .I2(__1740__),
    .I1(__1738__),
    .I0(__1736__),
    .O(__1745__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5429__ (
    .I5(__589__),
    .I4(__711__),
    .I3(__663__),
    .I2(__713__),
    .I1(__662__),
    .I0(__712__),
    .O(__1746__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __5430__ (
    .I1(__1446__),
    .I0(__1746__),
    .O(__1747__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5431__ (
    .I5(__589__),
    .I4(__702__),
    .I3(__663__),
    .I2(__707__),
    .I1(__662__),
    .I0(__703__),
    .O(__1748__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __5432__ (
    .I1(__1450__),
    .I0(__1748__),
    .O(__1749__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5433__ (
    .I5(__589__),
    .I4(__659__),
    .I3(__663__),
    .I2(__666__),
    .I1(__662__),
    .I0(__661__),
    .O(__1750__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5434__ (
    .I5(__589__),
    .I4(__778__),
    .I3(__663__),
    .I2(__780__),
    .I1(__662__),
    .I0(__779__),
    .O(__1751__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __5435__ (
    .I1(__1751__),
    .I0(__1750__),
    .O(__1752__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5436__ (
    .I5(__589__),
    .I4(__717__),
    .I3(__663__),
    .I2(__719__),
    .I1(__662__),
    .I0(__718__),
    .O(__1753__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __5437__ (
    .I1(__1442__),
    .I0(__1753__),
    .O(__1754__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5438__ (
    .I5(__589__),
    .I4(__723__),
    .I3(__663__),
    .I2(__725__),
    .I1(__662__),
    .I0(__724__),
    .O(__1755__)
  );
  LUT6 #(
    .INIT(64'h8e08ef8eef8e8e08)
  ) __5439__ (
    .I5(__1438__),
    .I4(__1755__),
    .I3(__1754__),
    .I2(__1752__),
    .I1(__1749__),
    .I0(__1747__),
    .O(__1756__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5440__ (
    .I5(__589__),
    .I4(__781__),
    .I3(__663__),
    .I2(__790__),
    .I1(__662__),
    .I0(__783__),
    .O(__1757__)
  );
  LUT4 #(
    .INIT(16'hf8ff)
  ) __5441__ (
    .I3(__603__),
    .I2(__1757__),
    .I1(__1756__),
    .I0(__1745__),
    .O(__1758__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5442__ (
    .I5(__589__),
    .I4(__414__),
    .I3(__663__),
    .I2(__417__),
    .I1(__662__),
    .I0(__415__),
    .O(__1759__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5443__ (
    .I5(__589__),
    .I4(__418__),
    .I3(__663__),
    .I2(__472__),
    .I1(__662__),
    .I0(__469__),
    .O(__1760__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5444__ (
    .I5(__589__),
    .I4(__473__),
    .I3(__663__),
    .I2(__480__),
    .I1(__662__),
    .I0(__475__),
    .O(__1761__)
  );
  LUT4 #(
    .INIT(16'hf3ba)
  ) __5445__ (
    .I3(__1761__),
    .I2(__1760__),
    .I1(__1759__),
    .I0(__1758__),
    .O(__1762__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5446__ (
    .I5(__589__),
    .I4(__824__),
    .I3(__663__),
    .I2(__827__),
    .I1(__662__),
    .I0(__826__),
    .O(__1763__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5447__ (
    .I5(__589__),
    .I4(__831__),
    .I3(__663__),
    .I2(__833__),
    .I1(__662__),
    .I0(__832__),
    .O(__1764__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5448__ (
    .I5(__589__),
    .I4(__846__),
    .I3(__663__),
    .I2(__849__),
    .I1(__662__),
    .I0(__847__),
    .O(__1765__)
  );
  LUT6 #(
    .INIT(64'h0000066006600000)
  ) __5449__ (
    .I5(__1436__),
    .I4(__1765__),
    .I3(__1446__),
    .I2(__1764__),
    .I1(__1450__),
    .I0(__1763__),
    .O(__1766__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5450__ (
    .I5(__589__),
    .I4(__834__),
    .I3(__663__),
    .I2(__836__),
    .I1(__662__),
    .I0(__835__),
    .O(__1767__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5451__ (
    .I5(__589__),
    .I4(__840__),
    .I3(__663__),
    .I2(__842__),
    .I1(__662__),
    .I0(__841__),
    .O(__1768__)
  );
  LUT4 #(
    .INIT(16'h1428)
  ) __5452__ (
    .I3(__1444__),
    .I2(__1440__),
    .I1(__1768__),
    .I0(__1767__),
    .O(__1769__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5453__ (
    .I5(__589__),
    .I4(__820__),
    .I3(__663__),
    .I2(__823__),
    .I1(__662__),
    .I0(__822__),
    .O(__1770__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5454__ (
    .I5(__589__),
    .I4(__837__),
    .I3(__663__),
    .I2(__839__),
    .I1(__662__),
    .I0(__838__),
    .O(__1771__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5455__ (
    .I5(__589__),
    .I4(__828__),
    .I3(__663__),
    .I2(__830__),
    .I1(__662__),
    .I0(__829__),
    .O(__1772__)
  );
  LUT6 #(
    .INIT(64'h0000099009900000)
  ) __5456__ (
    .I5(__1448__),
    .I4(__1772__),
    .I3(__1442__),
    .I2(__1771__),
    .I1(__1770__),
    .I0(__1742__),
    .O(__1773__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5457__ (
    .I5(__589__),
    .I4(__815__),
    .I3(__663__),
    .I2(__819__),
    .I1(__662__),
    .I0(__817__),
    .O(__1774__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5458__ (
    .I5(__589__),
    .I4(__843__),
    .I3(__663__),
    .I2(__845__),
    .I1(__662__),
    .I0(__844__),
    .O(__1775__)
  );
  LUT6 #(
    .INIT(64'h0041410000000000)
  ) __5459__ (
    .I5(__603__),
    .I4(__1438__),
    .I3(__1775__),
    .I2(__1751__),
    .I1(__1774__),
    .I0(__1757__),
    .O(__1776__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5460__ (
    .I5(__589__),
    .I4(__404__),
    .I3(__663__),
    .I2(__406__),
    .I1(__662__),
    .I0(__405__),
    .O(__1777__)
  );
  LUT5 #(
    .INIT(32'h00008000)
  ) __5461__ (
    .I4(__1777__),
    .I3(__1776__),
    .I2(__1773__),
    .I1(__1769__),
    .I0(__1766__),
    .O(__1778__)
  );
  LUT4 #(
    .INIT(16'h11f0)
  ) __5462__ (
    .I3(__663__),
    .I2(__480__),
    .I1(__1778__),
    .I0(__1762__),
    .O(__1779__)
  );
  LUT3 #(
    .INIT(8'h4f)
  ) __5463__ (
    .I2(__1479__),
    .I1(__1497__),
    .I0(__1480__),
    .O(__1780__)
  );
  LUT4 #(
    .INIT(16'hf044)
  ) __5464__ (
    .I3(__988__),
    .I2(__991__),
    .I1(__990__),
    .I0(__858__),
    .O(__1781__)
  );
  LUT6 #(
    .INIT(64'h00000000ccaaf0f0)
  ) __5465__ (
    .I5(__868__),
    .I4(__858__),
    .I3(__142__),
    .I2(__869__),
    .I1(__158__),
    .I0(__1781__),
    .O(__1782__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5466__ (
    .I1(__862__),
    .I0(__868__),
    .O(__1783__)
  );
  LUT6 #(
    .INIT(64'hff00ff00eeeef0f0)
  ) __5467__ (
    .I5(__300__),
    .I4(__858__),
    .I3(__303__),
    .I2(__302__),
    .I1(__1783__),
    .I0(__1782__),
    .O(__1784__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5468__ (
    .I5(__944__),
    .I4(__172__),
    .I3(__858__),
    .I2(__177__),
    .I1(__954__),
    .I0(__174__),
    .O(__1785__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5469__ (
    .I5(__944__),
    .I4(__180__),
    .I3(__858__),
    .I2(__189__),
    .I1(__954__),
    .I0(__186__),
    .O(__1786__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5470__ (
    .I5(__944__),
    .I4(__194__),
    .I3(__858__),
    .I2(__199__),
    .I1(__954__),
    .I0(__197__),
    .O(__1787__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5471__ (
    .I5(__944__),
    .I4(__153__),
    .I3(__858__),
    .I2(__154__),
    .I1(__954__),
    .I0(__336__),
    .O(__1788__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5472__ (
    .I5(__944__),
    .I4(__156__),
    .I3(__858__),
    .I2(__338__),
    .I1(__954__),
    .I0(__157__),
    .O(__1789__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5473__ (
    .I5(__944__),
    .I4(__285__),
    .I3(__858__),
    .I2(__298__),
    .I1(__954__),
    .I0(__292__),
    .O(__1790__)
  );
  LUT6 #(
    .INIT(64'h0000000000000008)
  ) __5474__ (
    .I5(__1790__),
    .I4(__1789__),
    .I3(__1788__),
    .I2(__1787__),
    .I1(__1786__),
    .I0(__1785__),
    .O(__1791__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5475__ (
    .I5(__944__),
    .I4(__201__),
    .I3(__858__),
    .I2(__204__),
    .I1(__954__),
    .I0(__202__),
    .O(__1792__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5476__ (
    .I5(__944__),
    .I4(__206__),
    .I3(__858__),
    .I2(__278__),
    .I1(__954__),
    .I0(__255__),
    .O(__1793__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5477__ (
    .I5(__944__),
    .I4(__245__),
    .I3(__858__),
    .I2(__213__),
    .I1(__954__),
    .I0(__228__),
    .O(__1794__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5478__ (
    .I5(__944__),
    .I4(__209__),
    .I3(__858__),
    .I2(__363__),
    .I1(__954__),
    .I0(__212__),
    .O(__1795__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5479__ (
    .I5(__944__),
    .I4(__170__),
    .I3(__858__),
    .I2(__169__),
    .I1(__954__),
    .I0(__166__),
    .O(__1796__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5480__ (
    .I5(__944__),
    .I4(__339__),
    .I3(__858__),
    .I2(__162__),
    .I1(__954__),
    .I0(__137__),
    .O(__1797__)
  );
  LUT6 #(
    .INIT(64'h0100000000000000)
  ) __5481__ (
    .I5(__1797__),
    .I4(__1796__),
    .I3(__1795__),
    .I2(__1794__),
    .I1(__1793__),
    .I0(__1792__),
    .O(__1798__)
  );
  LUT3 #(
    .INIT(8'h07)
  ) __5482__ (
    .I2(__1792__),
    .I1(__1798__),
    .I0(__1791__),
    .O(__1799__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5483__ (
    .I5(__944__),
    .I4(__274__),
    .I3(__858__),
    .I2(__276__),
    .I1(__954__),
    .I0(__275__),
    .O(__1800__)
  );
  LUT6 #(
    .INIT(64'h0001010000000000)
  ) __5484__ (
    .I5(__300__),
    .I4(__1800__),
    .I3(__1799__),
    .I2(__297__),
    .I1(g2637),
    .I0(__1784__),
    .O(__1801__)
  );
  LUT3 #(
    .INIT(8'h01)
  ) __5485__ (
    .I2(__297__),
    .I1(g2637),
    .I0(__1784__),
    .O(__1802__)
  );
  LUT6 #(
    .INIT(64'h000033330f0faf00)
  ) __5486__ (
    .I5(__354__),
    .I4(__356__),
    .I3(__242__),
    .I2(__1802__),
    .I1(__1801__),
    .I0(__234__),
    .O(__1803__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __5487__ (
    .I2(__1511__),
    .I1(__88__),
    .I0(__132__),
    .O(__1804__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5488__ (
    .I5(__944__),
    .I4(__947__),
    .I3(__858__),
    .I2(__951__),
    .I1(__954__),
    .I0(__949__),
    .O(__1805__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5489__ (
    .I5(__944__),
    .I4(__940__),
    .I3(__858__),
    .I2(__942__),
    .I1(__954__),
    .I0(__941__),
    .O(__1806__)
  );
  LUT6 #(
    .INIT(64'h4f0f4f0000000000)
  ) __5490__ (
    .I5(__954__),
    .I4(__1674__),
    .I3(__1806__),
    .I2(__1647__),
    .I1(__1036__),
    .I0(__1805__),
    .O(__1807__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5491__ (
    .I5(__944__),
    .I4(__980__),
    .I3(__858__),
    .I2(__982__),
    .I1(__954__),
    .I0(__981__),
    .O(__1808__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5492__ (
    .I5(__944__),
    .I4(__977__),
    .I3(__858__),
    .I2(__979__),
    .I1(__954__),
    .I0(__978__),
    .O(__1809__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5493__ (
    .I5(__944__),
    .I4(__983__),
    .I3(__858__),
    .I2(__985__),
    .I1(__954__),
    .I0(__984__),
    .O(__1810__)
  );
  LUT6 #(
    .INIT(64'hd8fad850d850d8fa)
  ) __5494__ (
    .I5(g3229),
    .I4(__1810__),
    .I3(__1809__),
    .I2(__981__),
    .I1(__1808__),
    .I0(__1807__),
    .O(__1811__)
  );
  LUT6 #(
    .INIT(64'h4f0f4f0000000000)
  ) __5495__ (
    .I5(__954__),
    .I4(__1649__),
    .I3(__1648__),
    .I2(__1647__),
    .I1(__968__),
    .I0(__1646__),
    .O(__1812__)
  );
  LUT6 #(
    .INIT(64'h4eeeeeeeeeee4eee)
  ) __5496__ (
    .I5(g3229),
    .I4(__1653__),
    .I3(__1652__),
    .I2(__1651__),
    .I1(__566__),
    .I0(__1812__),
    .O(__1813__)
  );
  LUT5 #(
    .INIT(32'h0030aaaa)
  ) __5497__ (
    .I4(__589__),
    .I3(__1543__),
    .I2(__1544__),
    .I1(__1542__),
    .I0(__1002__),
    .O(__1814__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __5498__ (
    .I5(__954__),
    .I4(__936__),
    .I3(__927__),
    .I2(__924__),
    .I1(__888__),
    .I0(__913__),
    .O(__1815__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5499__ (
    .I5(__944__),
    .I4(__682__),
    .I3(__858__),
    .I2(__684__),
    .I1(__954__),
    .I0(__683__),
    .O(__1816__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5500__ (
    .I5(__944__),
    .I4(__689__),
    .I3(__858__),
    .I2(__691__),
    .I1(__954__),
    .I0(__690__),
    .O(__1817__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5501__ (
    .I5(__944__),
    .I4(__679__),
    .I3(__858__),
    .I2(__681__),
    .I1(__954__),
    .I0(__680__),
    .O(__1818__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __5502__ (
    .I1(__1818__),
    .I0(__749__),
    .O(__1819__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5503__ (
    .I5(__944__),
    .I4(__692__),
    .I3(__858__),
    .I2(__694__),
    .I1(__954__),
    .I0(__693__),
    .O(__1820__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __5504__ (
    .I1(__765__),
    .I0(__1820__),
    .O(__1821__)
  );
  LUT6 #(
    .INIT(64'h1428000000000000)
  ) __5505__ (
    .I5(__1821__),
    .I4(__1819__),
    .I3(__770__),
    .I2(__772__),
    .I1(__1817__),
    .I0(__1816__),
    .O(__1822__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5506__ (
    .I5(__944__),
    .I4(__506__),
    .I3(__858__),
    .I2(__651__),
    .I1(__954__),
    .I0(__507__),
    .O(__1823__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5507__ (
    .I5(__944__),
    .I4(__696__),
    .I3(__858__),
    .I2(__698__),
    .I1(__954__),
    .I0(__697__),
    .O(__1824__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5508__ (
    .I1(__750__),
    .I0(__1824__),
    .O(__1825__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5509__ (
    .I5(__944__),
    .I4(__705__),
    .I3(__858__),
    .I2(__706__),
    .I1(__954__),
    .I0(__664__),
    .O(__1826__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __5510__ (
    .I1(__750__),
    .I0(__1824__),
    .O(__1827__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5511__ (
    .I5(__944__),
    .I4(__685__),
    .I3(__858__),
    .I2(__688__),
    .I1(__954__),
    .I0(__686__),
    .O(__1828__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __5512__ (
    .I1(__1828__),
    .I0(__741__),
    .O(__1829__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5513__ (
    .I5(__944__),
    .I4(__653__),
    .I3(__858__),
    .I2(__740__),
    .I1(__954__),
    .I0(__746__),
    .O(__1830__)
  );
  LUT4 #(
    .INIT(16'h7770)
  ) __5514__ (
    .I3(__768__),
    .I2(__1823__),
    .I1(__1828__),
    .I0(__741__),
    .O(__1831__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5515__ (
    .I5(__944__),
    .I4(__700__),
    .I3(__858__),
    .I2(__704__),
    .I1(__954__),
    .I0(__701__),
    .O(__1832__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __5516__ (
    .I1(__766__),
    .I0(__1832__),
    .O(__1833__)
  );
  LUT6 #(
    .INIT(64'h0110000000000000)
  ) __5517__ (
    .I5(__1833__),
    .I4(__1831__),
    .I3(__760__),
    .I2(__1830__),
    .I1(__1829__),
    .I0(__1827__),
    .O(__1834__)
  );
  LUT6 #(
    .INIT(64'h0007070000000000)
  ) __5518__ (
    .I5(__1834__),
    .I4(__767__),
    .I3(__1826__),
    .I2(__1825__),
    .I1(__768__),
    .I0(__1823__),
    .O(__1835__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5519__ (
    .I1(__944__),
    .I0(__676__),
    .O(__1836__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5520__ (
    .I5(__944__),
    .I4(__673__),
    .I3(__858__),
    .I2(__675__),
    .I1(__954__),
    .I0(__674__),
    .O(__1837__)
  );
  LUT6 #(
    .INIT(64'h00008acf00000000)
  ) __5521__ (
    .I5(__1837__),
    .I4(__1836__),
    .I3(__858__),
    .I2(__954__),
    .I1(__677__),
    .I0(__678__),
    .O(__1838__)
  );
  LUT4 #(
    .INIT(16'h0080)
  ) __5522__ (
    .I3(__745__),
    .I2(__764__),
    .I1(__573__),
    .I0(__954__),
    .O(__1839__)
  );
  LUT5 #(
    .INIT(32'h3f00aaaa)
  ) __5523__ (
    .I4(__1839__),
    .I3(__1838__),
    .I2(__1835__),
    .I1(__1822__),
    .I0(__671__),
    .O(__1840__)
  );
  LUT4 #(
    .INIT(16'haccc)
  ) __5524__ (
    .I3(__589__),
    .I2(__603__),
    .I1(__1289__),
    .I0(__1572__),
    .O(__1841__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5525__ (
    .I5(__858__),
    .I4(__486__),
    .I3(__944__),
    .I2(__249__),
    .I1(__954__),
    .I0(__346__),
    .O(__1842__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5526__ (
    .I1(__954__),
    .I0(__277__),
    .O(__1843__)
  );
  LUT6 #(
    .INIT(64'h0000000000bfbfbf)
  ) __5527__ (
    .I5(__1843__),
    .I4(__944__),
    .I3(__382__),
    .I2(__1347__),
    .I1(__306__),
    .I0(__1842__),
    .O(__1844__)
  );
  LUT6 #(
    .INIT(64'h4545ff000505ff00)
  ) __5528__ (
    .I5(__858__),
    .I4(__954__),
    .I3(__277__),
    .I2(__1844__),
    .I1(__279__),
    .I0(__1624__),
    .O(__1845__)
  );
  LUT4 #(
    .INIT(16'h0baa)
  ) __5529__ (
    .I3(__858__),
    .I2(__1624__),
    .I1(__1665__),
    .I0(__812__),
    .O(__1846__)
  );
  LUT6 #(
    .INIT(64'h132033005fa0ff00)
  ) __5530__ (
    .I5(__954__),
    .I4(__737__),
    .I3(__797__),
    .I2(__1047__),
    .I1(__875__),
    .I0(__1668__),
    .O(__1847__)
  );
  LUT6 #(
    .INIT(64'h00f07878f0f0f0f0)
  ) __5531__ (
    .I5(__589__),
    .I4(__1598__),
    .I3(__603__),
    .I2(__656__),
    .I1(__657__),
    .I0(__658__),
    .O(__1848__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __5532__ (
    .I5(__944__),
    .I4(__764__),
    .I3(__573__),
    .I2(__745__),
    .I1(__653__),
    .I0(__760__),
    .O(__1849__)
  );
  LUT5 #(
    .INIT(32'h6c9ccccc)
  ) __5533__ (
    .I4(__1761__),
    .I3(__1760__),
    .I2(__1759__),
    .I1(__1755__),
    .I0(__1735__),
    .O(__1850__)
  );
  LUT3 #(
    .INIT(8'h08)
  ) __5534__ (
    .I2(__1760__),
    .I1(__1761__),
    .I0(__1759__),
    .O(__1851__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __5535__ (
    .I1(__1750__),
    .I0(__1744__),
    .O(__1852__)
  );
  LUT5 #(
    .INIT(32'h80000000)
  ) __5536__ (
    .I4(__1748__),
    .I3(__1746__),
    .I2(__1739__),
    .I1(__1737__),
    .I0(__1735__),
    .O(__1853__)
  );
  LUT6 #(
    .INIT(64'h0100000000000000)
  ) __5537__ (
    .I5(__1853__),
    .I4(__1851__),
    .I3(__1852__),
    .I2(__1755__),
    .I1(__1753__),
    .I0(__1741__),
    .O(__1854__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5538__ (
    .I1(__1755__),
    .I0(__1753__),
    .O(__1855__)
  );
  LUT6 #(
    .INIT(64'h4000000000000000)
  ) __5539__ (
    .I5(__1750__),
    .I4(__1744__),
    .I3(__1741__),
    .I2(__1853__),
    .I1(__1855__),
    .I0(__1851__),
    .O(__1856__)
  );
  LUT4 #(
    .INIT(16'he000)
  ) __5540__ (
    .I3(__1761__),
    .I2(__1759__),
    .I1(__1856__),
    .I0(__1854__),
    .O(__1857__)
  );
  LUT4 #(
    .INIT(16'h8000)
  ) __5541__ (
    .I3(__1776__),
    .I2(__1773__),
    .I1(__1769__),
    .I0(__1766__),
    .O(__1858__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5542__ (
    .I1(__1760__),
    .I0(__1759__),
    .O(__1859__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5543__ (
    .I5(__589__),
    .I4(__407__),
    .I3(__663__),
    .I2(__411__),
    .I1(__662__),
    .I0(__408__),
    .O(__1860__)
  );
  LUT6 #(
    .INIT(64'h0000000000008000)
  ) __5544__ (
    .I5(__1761__),
    .I4(__1860__),
    .I3(__1859__),
    .I2(__1756__),
    .I1(__1745__),
    .I0(__1858__),
    .O(__1861__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5545__ (
    .I1(__1760__),
    .I0(__1759__),
    .O(__1862__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5546__ (
    .I1(__603__),
    .I0(__1757__),
    .O(__1863__)
  );
  LUT6 #(
    .INIT(64'hff00ffff0b000f0f)
  ) __5547__ (
    .I5(__1761__),
    .I4(__1858__),
    .I3(__1777__),
    .I2(__1863__),
    .I1(__1862__),
    .I0(__1860__),
    .O(__1864__)
  );
  LUT6 #(
    .INIT(64'hf0f03355f0f0f0f0)
  ) __5548__ (
    .I5(__1864__),
    .I4(__1861__),
    .I3(__1857__),
    .I2(__1438__),
    .I1(__1851__),
    .I0(__1850__),
    .O(__1865__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __5549__ (
    .I2(__662__),
    .I1(__1865__),
    .I0(__724__),
    .O(__1866__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __5550__ (
    .I2(__1479__),
    .I1(__1443__),
    .I0(__1465__),
    .O(__1867__)
  );
  LUT6 #(
    .INIT(64'h4000000000000000)
  ) __5551__ (
    .I5(__944__),
    .I4(__918__),
    .I3(__917__),
    .I2(__920__),
    .I1(__921__),
    .I0(__924__),
    .O(__1868__)
  );
  LUT4 #(
    .INIT(16'h8000)
  ) __5552__ (
    .I3(__915__),
    .I2(__916__),
    .I1(__914__),
    .I0(__1868__),
    .O(__1869__)
  );
  LUT5 #(
    .INIT(32'h12305af0)
  ) __5553__ (
    .I4(__954__),
    .I3(__913__),
    .I2(__912__),
    .I1(__925__),
    .I0(__1869__),
    .O(__1870__)
  );
  LUT2 #(
    .INIT(4'h7)
  ) __5554__ (
    .I1(__1543__),
    .I0(__1542__),
    .O(__1871__)
  );
  LUT6 #(
    .INIT(64'h5555fccf55555555)
  ) __5555__ (
    .I5(__1592__),
    .I4(__1588__),
    .I3(__1546__),
    .I2(__1871__),
    .I1(__1555__),
    .I0(__1417__),
    .O(__1872__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __5556__ (
    .I2(__589__),
    .I1(__1872__),
    .I0(__1274__),
    .O(__1873__)
  );
  LUT6 #(
    .INIT(64'h4000000000000000)
  ) __5557__ (
    .I5(__589__),
    .I4(__1178__),
    .I3(__1176__),
    .I2(__1180__),
    .I1(__1175__),
    .I0(__1598__),
    .O(__1874__)
  );
  LUT6 #(
    .INIT(64'h0078787878787878)
  ) __5558__ (
    .I5(__589__),
    .I4(__1598__),
    .I3(__603__),
    .I2(__1164__),
    .I1(__1174__),
    .I0(__1874__),
    .O(__1875__)
  );
  LUT5 #(
    .INIT(32'h0030aaaa)
  ) __5559__ (
    .I4(__663__),
    .I3(__1681__),
    .I2(__1682__),
    .I1(__1680__),
    .I0(__379__),
    .O(__1876__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5560__ (
    .I5(__589__),
    .I4(__1243__),
    .I3(__663__),
    .I2(__1226__),
    .I1(__662__),
    .I0(__1225__),
    .O(__1877__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __5561__ (
    .I1(__1453__),
    .I0(__1877__),
    .O(__1878__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5562__ (
    .I5(__589__),
    .I4(__1213__),
    .I3(__663__),
    .I2(__71__),
    .I1(__662__),
    .I0(__1218__),
    .O(__1879__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __5563__ (
    .I1(__1457__),
    .I0(__1879__),
    .O(__1880__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5564__ (
    .I5(__589__),
    .I4(__1202__),
    .I3(__663__),
    .I2(__1205__),
    .I1(__662__),
    .I0(__1203__),
    .O(__1881__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __5565__ (
    .I1(__1459__),
    .I0(__1881__),
    .O(__1882__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5566__ (
    .I5(__589__),
    .I4(__1160__),
    .I3(__663__),
    .I2(__1204__),
    .I1(__662__),
    .I0(__649__),
    .O(__1883__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5567__ (
    .I5(__589__),
    .I4(__1258__),
    .I3(__663__),
    .I2(__1259__),
    .I1(__662__),
    .I0(__1263__),
    .O(__1884__)
  );
  LUT2 #(
    .INIT(4'h9)
  ) __5568__ (
    .I1(__1884__),
    .I0(__1883__),
    .O(__1885__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5569__ (
    .I5(__589__),
    .I4(__793__),
    .I3(__663__),
    .I2(__736__),
    .I1(__662__),
    .I0(__1044__),
    .O(__1886__)
  );
  LUT6 #(
    .INIT(64'he880fee8fee8e880)
  ) __5570__ (
    .I5(__1455__),
    .I4(__1886__),
    .I3(__1885__),
    .I2(__1882__),
    .I1(__1880__),
    .I0(__1878__),
    .O(__1887__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5571__ (
    .I5(__589__),
    .I4(__1207__),
    .I3(__663__),
    .I2(__1217__),
    .I1(__662__),
    .I0(__1216__),
    .O(__1888__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __5572__ (
    .I1(__1458__),
    .I0(__1888__),
    .O(__1889__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5573__ (
    .I5(__589__),
    .I4(__1198__),
    .I3(__663__),
    .I2(__1201__),
    .I1(__662__),
    .I0(__1200__),
    .O(__1890__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __5574__ (
    .I1(__1460__),
    .I0(__1890__),
    .O(__1891__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5575__ (
    .I5(__589__),
    .I4(__1182__),
    .I3(__663__),
    .I2(__1165__),
    .I1(__662__),
    .I0(__1173__),
    .O(__1892__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5576__ (
    .I5(__589__),
    .I4(__1229__),
    .I3(__663__),
    .I2(__1230__),
    .I1(__662__),
    .I0(__1260__),
    .O(__1893__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __5577__ (
    .I1(__1893__),
    .I0(__1892__),
    .O(__1894__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5578__ (
    .I5(__589__),
    .I4(__1045__),
    .I3(__663__),
    .I2(__728__),
    .I1(__662__),
    .I0(__726__),
    .O(__1895__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __5579__ (
    .I1(__1456__),
    .I0(__1895__),
    .O(__1896__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5580__ (
    .I5(__589__),
    .I4(__534__),
    .I3(__663__),
    .I2(__1221__),
    .I1(__662__),
    .I0(__535__),
    .O(__1897__)
  );
  LUT6 #(
    .INIT(64'h8e08ef8eef8e8e08)
  ) __5581__ (
    .I5(__1454__),
    .I4(__1897__),
    .I3(__1896__),
    .I2(__1894__),
    .I1(__1891__),
    .I0(__1889__),
    .O(__1898__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5582__ (
    .I5(__589__),
    .I4(__1231__),
    .I3(__663__),
    .I2(__1233__),
    .I1(__662__),
    .I0(__1264__),
    .O(__1899__)
  );
  LUT4 #(
    .INIT(16'hf8ff)
  ) __5583__ (
    .I3(__603__),
    .I2(__1899__),
    .I1(__1898__),
    .I0(__1887__),
    .O(__1900__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5584__ (
    .I5(__589__),
    .I4(__1266__),
    .I3(__663__),
    .I2(__774__),
    .I1(__662__),
    .I0(__342__),
    .O(__1901__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5585__ (
    .I5(__589__),
    .I4(__1328__),
    .I3(__663__),
    .I2(__1331__),
    .I1(__662__),
    .I0(__1330__),
    .O(__1902__)
  );
  LUT6 #(
    .INIT(64'h0041410000000000)
  ) __5586__ (
    .I5(__603__),
    .I4(__1454__),
    .I3(__1902__),
    .I2(__1893__),
    .I1(__1901__),
    .I0(__1899__),
    .O(__1903__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5587__ (
    .I5(__589__),
    .I4(__785__),
    .I3(__663__),
    .I2(__792__),
    .I1(__662__),
    .I0(__800__),
    .O(__1904__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5588__ (
    .I5(__589__),
    .I4(__1312__),
    .I3(__663__),
    .I2(__1324__),
    .I1(__662__),
    .I0(__1117__),
    .O(__1905__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5589__ (
    .I5(__589__),
    .I4(__652__),
    .I3(__663__),
    .I2(__1304__),
    .I1(__662__),
    .I0(__1301__),
    .O(__1906__)
  );
  LUT6 #(
    .INIT(64'h0000099009900000)
  ) __5590__ (
    .I5(__1459__),
    .I4(__1906__),
    .I3(__1456__),
    .I2(__1905__),
    .I1(__1904__),
    .I0(__1884__),
    .O(__1907__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5591__ (
    .I5(__589__),
    .I4(__1309__),
    .I3(__663__),
    .I2(__1311__),
    .I1(__662__),
    .I0(__1310__),
    .O(__1908__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5592__ (
    .I5(__589__),
    .I4(__1325__),
    .I3(__663__),
    .I2(__1327__),
    .I1(__662__),
    .I0(__1326__),
    .O(__1909__)
  );
  LUT4 #(
    .INIT(16'h1428)
  ) __5593__ (
    .I3(__1457__),
    .I2(__1455__),
    .I1(__1909__),
    .I0(__1908__),
    .O(__1910__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5594__ (
    .I5(__589__),
    .I4(__1049__),
    .I3(__663__),
    .I2(__735__),
    .I1(__662__),
    .I0(__795__),
    .O(__1911__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5595__ (
    .I5(__589__),
    .I4(__1306__),
    .I3(__663__),
    .I2(__1308__),
    .I1(__662__),
    .I0(__1307__),
    .O(__1912__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5596__ (
    .I5(__589__),
    .I4(__1335__),
    .I3(__663__),
    .I2(__1339__),
    .I1(__662__),
    .I0(__1337__),
    .O(__1913__)
  );
  LUT6 #(
    .INIT(64'h0000066006600000)
  ) __5597__ (
    .I5(__1453__),
    .I4(__1913__),
    .I3(__1458__),
    .I2(__1912__),
    .I1(__1460__),
    .I0(__1911__),
    .O(__1914__)
  );
  LUT5 #(
    .INIT(32'h80000000)
  ) __5598__ (
    .I4(__1914__),
    .I3(__1910__),
    .I2(__1907__),
    .I1(__1903__),
    .I0(__1900__),
    .O(__1915__)
  );
  LUT6 #(
    .INIT(64'h4000000000000000)
  ) __5599__ (
    .I5(__1596__),
    .I4(__1914__),
    .I3(__1910__),
    .I2(__1907__),
    .I1(__1903__),
    .I0(__1595__),
    .O(__1916__)
  );
  LUT4 #(
    .INIT(16'h1428)
  ) __5600__ (
    .I3(__1453__),
    .I2(__1455__),
    .I1(__1886__),
    .I0(__1877__),
    .O(__1917__)
  );
  LUT4 #(
    .INIT(16'h0990)
  ) __5601__ (
    .I3(__1460__),
    .I2(__1890__),
    .I1(__1893__),
    .I0(__1892__),
    .O(__1918__)
  );
  LUT4 #(
    .INIT(16'h1428)
  ) __5602__ (
    .I3(__1456__),
    .I2(__1454__),
    .I1(__1897__),
    .I0(__1895__),
    .O(__1919__)
  );
  LUT4 #(
    .INIT(16'h0990)
  ) __5603__ (
    .I3(__1459__),
    .I2(__1881__),
    .I1(__1884__),
    .I0(__1883__),
    .O(__1920__)
  );
  LUT6 #(
    .INIT(64'h8000000000000000)
  ) __5604__ (
    .I5(__1889__),
    .I4(__1880__),
    .I3(__1920__),
    .I2(__1919__),
    .I1(__1918__),
    .I0(__1917__),
    .O(__1921__)
  );
  LUT3 #(
    .INIT(8'h10)
  ) __5605__ (
    .I2(__1596__),
    .I1(__1597__),
    .I0(__1595__),
    .O(__1922__)
  );
  LUT5 #(
    .INIT(32'hcd000000)
  ) __5606__ (
    .I4(__589__),
    .I3(__603__),
    .I2(__1899__),
    .I1(__1922__),
    .I0(__1921__),
    .O(__1923__)
  );
  LUT6 #(
    .INIT(64'hffff0707ff00ff00)
  ) __5607__ (
    .I5(__1923__),
    .I4(__1597__),
    .I3(__1077__),
    .I2(__1916__),
    .I1(__1595__),
    .I0(__1915__),
    .O(__1924__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5608__ (
    .I5(__858__),
    .I4(__316__),
    .I3(__944__),
    .I2(__312__),
    .I1(__954__),
    .I0(__314__),
    .O(__1925__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5609__ (
    .I5(__858__),
    .I4(__328__),
    .I3(__944__),
    .I2(__324__),
    .I1(__954__),
    .I0(__326__),
    .O(__1926__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5610__ (
    .I5(__858__),
    .I4(__322__),
    .I3(__944__),
    .I2(__318__),
    .I1(__954__),
    .I0(__320__),
    .O(__1927__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5611__ (
    .I5(__944__),
    .I4(__128__),
    .I3(__858__),
    .I2(__131__),
    .I1(__954__),
    .I0(__130__),
    .O(__1928__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5612__ (
    .I5(__944__),
    .I4(__122__),
    .I3(__858__),
    .I2(__126__),
    .I1(__954__),
    .I0(__124__),
    .O(__1929__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5613__ (
    .I5(__944__),
    .I4(__136__),
    .I3(__858__),
    .I2(__139__),
    .I1(__954__),
    .I0(__138__),
    .O(__1930__)
  );
  LUT6 #(
    .INIT(64'h0fff0fff88ccffff)
  ) __5614__ (
    .I5(__1930__),
    .I4(__1926__),
    .I3(__1929__),
    .I2(__1925__),
    .I1(__1928__),
    .I0(__1927__),
    .O(__1931__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5615__ (
    .I5(__944__),
    .I4(__133__),
    .I3(__858__),
    .I2(__135__),
    .I1(__954__),
    .I0(__134__),
    .O(__1932__)
  );
  LUT6 #(
    .INIT(64'hff000e00ff00ff00)
  ) __5616__ (
    .I5(__1928__),
    .I4(__1932__),
    .I3(__1931__),
    .I2(__1927__),
    .I1(__1926__),
    .I0(__1925__),
    .O(__1933__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5617__ (
    .I5(__858__),
    .I4(__334__),
    .I3(__944__),
    .I2(__330__),
    .I1(__954__),
    .I0(__332__),
    .O(__1934__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __5618__ (
    .I1(__1934__),
    .I0(__1933__),
    .O(__1935__)
  );
  LUT5 #(
    .INIT(32'h00000080)
  ) __5619__ (
    .I4(__1926__),
    .I3(__1927__),
    .I2(__1932__),
    .I1(__1934__),
    .I0(__1930__),
    .O(__1936__)
  );
  LUT6 #(
    .INIT(64'h00f000ff00ff00bb)
  ) __5620__ (
    .I5(__1930__),
    .I4(__1925__),
    .I3(__1936__),
    .I2(__1928__),
    .I1(__1934__),
    .I0(__1929__),
    .O(__1937__)
  );
  LUT6 #(
    .INIT(64'hfffffffc54fcffff)
  ) __5621__ (
    .I5(__1930__),
    .I4(__1926__),
    .I3(__1934__),
    .I2(__1927__),
    .I1(__1928__),
    .I0(__1932__),
    .O(__1938__)
  );
  LUT6 #(
    .INIT(64'h3b33000f00000000)
  ) __5622__ (
    .I5(__1927__),
    .I4(__1934__),
    .I3(__1932__),
    .I2(__1926__),
    .I1(__1929__),
    .I0(__1928__),
    .O(__1939__)
  );
  LUT3 #(
    .INIT(8'h08)
  ) __5623__ (
    .I2(__1939__),
    .I1(__1938__),
    .I0(__1937__),
    .O(__1940__)
  );
  LUT3 #(
    .INIT(8'h70)
  ) __5624__ (
    .I2(__1627__),
    .I1(__858__),
    .I0(__115__),
    .O(__1941__)
  );
  LUT6 #(
    .INIT(64'hf0f0fff3fff3ffa2)
  ) __5625__ (
    .I5(__1926__),
    .I4(__1928__),
    .I3(__1930__),
    .I2(__1932__),
    .I1(__1927__),
    .I0(__1925__),
    .O(__1942__)
  );
  LUT6 #(
    .INIT(64'h7f7f007fffffffff)
  ) __5626__ (
    .I5(__1930__),
    .I4(__1928__),
    .I3(__1926__),
    .I2(__1927__),
    .I1(__1932__),
    .I0(__1929__),
    .O(__1943__)
  );
  LUT6 #(
    .INIT(64'hfe0fffffffffffff)
  ) __5627__ (
    .I5(__1932__),
    .I4(__1928__),
    .I3(__1930__),
    .I2(__1925__),
    .I1(__1926__),
    .I0(__1934__),
    .O(__1944__)
  );
  LUT6 #(
    .INIT(64'hffffff55ffffbcfc)
  ) __5628__ (
    .I5(__1926__),
    .I4(__1927__),
    .I3(__1932__),
    .I2(__1934__),
    .I1(__1929__),
    .I0(__1930__),
    .O(__1945__)
  );
  LUT5 #(
    .INIT(32'hac000000)
  ) __5629__ (
    .I4(__1945__),
    .I3(__1944__),
    .I2(__1934__),
    .I1(__1943__),
    .I0(__1942__),
    .O(__1946__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5630__ (
    .I5(__858__),
    .I4(__260__),
    .I3(__944__),
    .I2(__256__),
    .I1(__954__),
    .I0(__258__),
    .O(__1947__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5631__ (
    .I1(__954__),
    .I0(__120__),
    .O(__1948__)
  );
  LUT6 #(
    .INIT(64'h0000000000bfbfbf)
  ) __5632__ (
    .I5(__1948__),
    .I4(__944__),
    .I3(__116__),
    .I2(__1347__),
    .I1(__262__),
    .I0(__1947__),
    .O(__1949__)
  );
  LUT6 #(
    .INIT(64'h4f440000ffcc0000)
  ) __5633__ (
    .I5(__858__),
    .I4(__1624__),
    .I3(__1949__),
    .I2(__121__),
    .I1(__1627__),
    .I0(__115__),
    .O(__1950__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5634__ (
    .I5(__944__),
    .I4(__110__),
    .I3(__858__),
    .I2(__112__),
    .I1(__954__),
    .I0(__111__),
    .O(__1951__)
  );
  LUT6 #(
    .INIT(64'h5455555555555555)
  ) __5635__ (
    .I5(__1623__),
    .I4(__1506__),
    .I3(__1505__),
    .I2(__1508__),
    .I1(__1507__),
    .I0(__1951__),
    .O(__1952__)
  );
  LUT6 #(
    .INIT(64'hffffffffbf000000)
  ) __5636__ (
    .I5(__1952__),
    .I4(__1950__),
    .I3(__1946__),
    .I2(__1941__),
    .I1(__1940__),
    .I0(__1935__),
    .O(__1953__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __5637__ (
    .I2(__954__),
    .I1(__1953__),
    .I0(__111__),
    .O(__1954__)
  );
  LUT4 #(
    .INIT(16'haccc)
  ) __5638__ (
    .I3(__589__),
    .I2(__603__),
    .I1(__1266__),
    .I0(__1893__),
    .O(__1955__)
  );
  LUT4 #(
    .INIT(16'haccc)
  ) __5639__ (
    .I3(__662__),
    .I2(__603__),
    .I1(__592__),
    .I0(__1712__),
    .O(__1956__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5640__ (
    .I5(__589__),
    .I4(__547__),
    .I3(__663__),
    .I2(__594__),
    .I1(__662__),
    .I0(__548__),
    .O(__1957__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __5641__ (
    .I2(__663__),
    .I1(__1957__),
    .I0(__477__),
    .O(__1958__)
  );
  LUT5 #(
    .INIT(32'h81000000)
  ) __5642__ (
    .I4(__1682__),
    .I3(__1680__),
    .I2(__1681__),
    .I1(__1679__),
    .I0(__1677__),
    .O(__1959__)
  );
  LUT6 #(
    .INIT(64'h4000000200000000)
  ) __5643__ (
    .I5(__1959__),
    .I4(__1686__),
    .I3(__1691__),
    .I2(__1678__),
    .I1(__1689__),
    .I0(__1684__),
    .O(__1960__)
  );
  LUT5 #(
    .INIT(32'hdff72008)
  ) __5644__ (
    .I4(__1685__),
    .I3(__1692__),
    .I2(__1690__),
    .I1(__1684__),
    .I0(__1960__),
    .O(__1961__)
  );
  LUT6 #(
    .INIT(64'h0f0f33550f0f0f0f)
  ) __5645__ (
    .I5(__1732__),
    .I4(__1728__),
    .I3(__1697__),
    .I2(__1705__),
    .I1(__1684__),
    .I0(__1961__),
    .O(__1962__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __5646__ (
    .I2(__663__),
    .I1(__1962__),
    .I0(__609__),
    .O(__1963__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __5647__ (
    .I2(__589__),
    .I1(__1598__),
    .I0(__1635__),
    .O(__1964__)
  );
  LUT6 #(
    .INIT(64'h55555d5500000800)
  ) __5648__ (
    .I5(__1286__),
    .I4(__1430__),
    .I3(__1426__),
    .I2(__1428__),
    .I1(__1432__),
    .I0(__1964__),
    .O(__1965__)
  );
  LUT3 #(
    .INIT(8'hea)
  ) __5649__ (
    .I2(__862__),
    .I1(__868__),
    .I0(__1782__),
    .O(__1966__)
  );
  LUT5 #(
    .INIT(32'hdff72008)
  ) __5650__ (
    .I4(__1536__),
    .I3(__1550__),
    .I2(__1548__),
    .I1(__1545__),
    .I0(__1656__),
    .O(__1967__)
  );
  LUT6 #(
    .INIT(64'h0f0f33550f0f0f0f)
  ) __5651__ (
    .I5(__1592__),
    .I4(__1588__),
    .I3(__1555__),
    .I2(__1565__),
    .I1(__1545__),
    .I0(__1967__),
    .O(__1968__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __5652__ (
    .I2(__662__),
    .I1(__1968__),
    .I0(__1242__),
    .O(__1969__)
  );
  LUT6 #(
    .INIT(64'h132033005fa0ff00)
  ) __5653__ (
    .I5(__954__),
    .I4(__915__),
    .I3(__914__),
    .I2(__916__),
    .I1(__925__),
    .I0(__1868__),
    .O(__1970__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __5654__ (
    .I2(__944__),
    .I1(__1624__),
    .I0(__273__),
    .O(__1971__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5655__ (
    .I5(__589__),
    .I4(__1073__),
    .I3(__663__),
    .I2(__1075__),
    .I1(__662__),
    .I0(__1074__),
    .O(__1972__)
  );
  LUT5 #(
    .INIT(32'h80000000)
  ) __5656__ (
    .I4(__1972__),
    .I3(__1914__),
    .I2(__1910__),
    .I1(__1907__),
    .I0(__1903__),
    .O(__1973__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __5657__ (
    .I3(__662__),
    .I2(__603__),
    .I1(__1973__),
    .I0(__1074__),
    .O(__1974__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5658__ (
    .I5(__858__),
    .I4(__443__),
    .I3(__944__),
    .I2(__251__),
    .I1(__954__),
    .I0(__350__),
    .O(__1975__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5659__ (
    .I5(__944__),
    .I4(__283__),
    .I3(__858__),
    .I2(__286__),
    .I1(__954__),
    .I0(__284__),
    .O(__1976__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5660__ (
    .I5(__944__),
    .I4(__290__),
    .I3(__858__),
    .I2(__293__),
    .I1(__954__),
    .I0(__291__),
    .O(__1977__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5661__ (
    .I5(__944__),
    .I4(__287__),
    .I3(__858__),
    .I2(__289__),
    .I1(__954__),
    .I0(__288__),
    .O(__1978__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5662__ (
    .I5(__944__),
    .I4(__294__),
    .I3(__858__),
    .I2(__296__),
    .I1(__954__),
    .I0(__295__),
    .O(__1979__)
  );
  LUT5 #(
    .INIT(32'haa20cf45)
  ) __5663__ (
    .I4(g3229),
    .I3(__1979__),
    .I2(__1978__),
    .I1(__1977__),
    .I0(__1976__),
    .O(__1980__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5664__ (
    .I5(__944__),
    .I4(__145__),
    .I3(__858__),
    .I2(__270__),
    .I1(__954__),
    .I0(__268__),
    .O(__1981__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5665__ (
    .I5(__944__),
    .I4(__271__),
    .I3(__858__),
    .I2(__272__),
    .I1(__954__),
    .I0(__205__),
    .O(__1982__)
  );
  LUT6 #(
    .INIT(64'h4f0f4f0000000000)
  ) __5666__ (
    .I5(__954__),
    .I4(__1982__),
    .I3(__1981__),
    .I2(__1647__),
    .I1(__354__),
    .I0(__1800__),
    .O(__1983__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __5667__ (
    .I2(__1983__),
    .I1(__1980__),
    .I0(__295__),
    .O(__1984__)
  );
  LUT6 #(
    .INIT(64'h4000000000000000)
  ) __5668__ (
    .I5(__944__),
    .I4(__768__),
    .I3(__767__),
    .I2(__760__),
    .I1(__766__),
    .I0(__745__),
    .O(__1985__)
  );
  LUT4 #(
    .INIT(16'h8000)
  ) __5669__ (
    .I3(__772__),
    .I2(__765__),
    .I1(__750__),
    .I0(__1985__),
    .O(__1986__)
  );
  LUT4 #(
    .INIT(16'h125a)
  ) __5670__ (
    .I3(__954__),
    .I2(__741__),
    .I1(__752__),
    .I0(__1986__),
    .O(__1987__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __5671__ (
    .I5(__764__),
    .I4(__573__),
    .I3(__858__),
    .I2(__745__),
    .I1(__681__),
    .I0(__749__),
    .O(__1988__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __5672__ (
    .I2(__663__),
    .I1(__1872__),
    .I0(__1276__),
    .O(__1989__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __5673__ (
    .I5(__944__),
    .I4(__764__),
    .I3(__573__),
    .I2(__745__),
    .I1(__700__),
    .I0(__766__),
    .O(__1990__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __5674__ (
    .I5(__954__),
    .I4(__936__),
    .I3(__927__),
    .I2(__924__),
    .I1(__906__),
    .I0(__920__),
    .O(__1991__)
  );
  LUT6 #(
    .INIT(64'h0f007f00ff00ff00)
  ) __5675__ (
    .I5(__603__),
    .I4(__1757__),
    .I3(__1760__),
    .I2(__1759__),
    .I1(__1756__),
    .I0(__1745__),
    .O(__1992__)
  );
  LUT4 #(
    .INIT(16'h1428)
  ) __5676__ (
    .I3(__1440__),
    .I2(__1436__),
    .I1(__1735__),
    .I0(__1744__),
    .O(__1993__)
  );
  LUT4 #(
    .INIT(16'h0990)
  ) __5677__ (
    .I3(__1450__),
    .I2(__1748__),
    .I1(__1751__),
    .I0(__1750__),
    .O(__1994__)
  );
  LUT4 #(
    .INIT(16'h1428)
  ) __5678__ (
    .I3(__1438__),
    .I2(__1442__),
    .I1(__1753__),
    .I0(__1755__),
    .O(__1995__)
  );
  LUT4 #(
    .INIT(16'h0990)
  ) __5679__ (
    .I3(__1448__),
    .I2(__1739__),
    .I1(__1742__),
    .I0(__1741__),
    .O(__1996__)
  );
  LUT6 #(
    .INIT(64'h8000000000000000)
  ) __5680__ (
    .I5(__1747__),
    .I4(__1738__),
    .I3(__1996__),
    .I2(__1995__),
    .I1(__1994__),
    .I0(__1993__),
    .O(__1997__)
  );
  LUT5 #(
    .INIT(32'hfcf9f0f0)
  ) __5681__ (
    .I4(__603__),
    .I3(__1757__),
    .I2(__1760__),
    .I1(__1759__),
    .I0(__1997__),
    .O(__1998__)
  );
  LUT6 #(
    .INIT(64'h00000000bfffffff)
  ) __5682__ (
    .I5(__1761__),
    .I4(__1776__),
    .I3(__1773__),
    .I2(__1769__),
    .I1(__1766__),
    .I0(__1777__),
    .O(__1999__)
  );
  LUT6 #(
    .INIT(64'hcf300000aaaaaaaa)
  ) __5683__ (
    .I5(__663__),
    .I4(__1999__),
    .I3(__1759__),
    .I2(__1998__),
    .I1(__1992__),
    .I0(__417__),
    .O(__2000__)
  );
  LUT6 #(
    .INIT(64'h9333363333333333)
  ) __5684__ (
    .I5(__1597__),
    .I4(__1596__),
    .I3(__1595__),
    .I2(__1897__),
    .I1(__1886__),
    .I0(__1877__),
    .O(__2001__)
  );
  LUT3 #(
    .INIT(8'h08)
  ) __5685__ (
    .I2(__1596__),
    .I1(__1597__),
    .I0(__1595__),
    .O(__2002__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __5686__ (
    .I1(__1892__),
    .I0(__1886__),
    .O(__2003__)
  );
  LUT5 #(
    .INIT(32'h80000000)
  ) __5687__ (
    .I4(__1890__),
    .I3(__1888__),
    .I2(__1881__),
    .I1(__1879__),
    .I0(__1877__),
    .O(__2004__)
  );
  LUT6 #(
    .INIT(64'h0100000000000000)
  ) __5688__ (
    .I5(__2004__),
    .I4(__2002__),
    .I3(__2003__),
    .I2(__1897__),
    .I1(__1895__),
    .I0(__1883__),
    .O(__2005__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5689__ (
    .I1(__1897__),
    .I0(__1895__),
    .O(__2006__)
  );
  LUT6 #(
    .INIT(64'h4000000000000000)
  ) __5690__ (
    .I5(__1892__),
    .I4(__1886__),
    .I3(__1883__),
    .I2(__2004__),
    .I1(__2006__),
    .I0(__2002__),
    .O(__2007__)
  );
  LUT4 #(
    .INIT(16'he000)
  ) __5691__ (
    .I3(__1597__),
    .I2(__1595__),
    .I1(__2007__),
    .I0(__2005__),
    .O(__2008__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5692__ (
    .I5(__589__),
    .I4(__1077__),
    .I3(__663__),
    .I2(__1080__),
    .I1(__662__),
    .I0(__1078__),
    .O(__2009__)
  );
  LUT3 #(
    .INIT(8'h08)
  ) __5693__ (
    .I2(__2009__),
    .I1(__1596__),
    .I0(__1595__),
    .O(__2010__)
  );
  LUT4 #(
    .INIT(16'h8000)
  ) __5694__ (
    .I3(__1914__),
    .I2(__1910__),
    .I1(__1907__),
    .I0(__1903__),
    .O(__2011__)
  );
  LUT5 #(
    .INIT(32'h00008000)
  ) __5695__ (
    .I4(__1597__),
    .I3(__2011__),
    .I2(__2010__),
    .I1(__1898__),
    .I0(__1887__),
    .O(__2012__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5696__ (
    .I1(__1596__),
    .I0(__1595__),
    .O(__2013__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5697__ (
    .I1(__603__),
    .I0(__1899__),
    .O(__2014__)
  );
  LUT6 #(
    .INIT(64'hff00ffff0b000f0f)
  ) __5698__ (
    .I5(__1597__),
    .I4(__2011__),
    .I3(__1972__),
    .I2(__2014__),
    .I1(__2013__),
    .I0(__2009__),
    .O(__2015__)
  );
  LUT6 #(
    .INIT(64'hf0f033aaf0f0f0f0)
  ) __5699__ (
    .I5(__2015__),
    .I4(__2012__),
    .I3(__2008__),
    .I2(__1455__),
    .I1(__2002__),
    .I0(__2001__),
    .O(__2016__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __5700__ (
    .I2(__662__),
    .I1(__2016__),
    .I0(__1044__),
    .O(__2017__)
  );
  LUT2 #(
    .INIT(4'h7)
  ) __5701__ (
    .I1(__1761__),
    .I0(__1759__),
    .O(__2018__)
  );
  LUT6 #(
    .INIT(64'h5555fccf55555555)
  ) __5702__ (
    .I5(__1864__),
    .I4(__1861__),
    .I3(__1735__),
    .I2(__2018__),
    .I1(__1857__),
    .I0(__1436__),
    .O(__2019__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __5703__ (
    .I2(__662__),
    .I1(__2019__),
    .I0(__739__),
    .O(__2020__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5704__ (
    .I5(__858__),
    .I4(__1015__),
    .I3(__944__),
    .I2(__1011__),
    .I1(__954__),
    .I0(__1013__),
    .O(__2021__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5705__ (
    .I1(__954__),
    .I0(__953__),
    .O(__2022__)
  );
  LUT6 #(
    .INIT(64'h0000000000bfbfbf)
  ) __5706__ (
    .I5(__2022__),
    .I4(__944__),
    .I3(__952__),
    .I2(__1347__),
    .I1(__993__),
    .I0(__2021__),
    .O(__2023__)
  );
  LUT6 #(
    .INIT(64'h4545ff000505ff00)
  ) __5707__ (
    .I5(__858__),
    .I4(__944__),
    .I3(__952__),
    .I2(__2023__),
    .I1(__955__),
    .I0(__1624__),
    .O(__2024__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __5708__ (
    .I2(__944__),
    .I1(__354__),
    .I0(__231__),
    .O(__2025__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __5709__ (
    .I2(__1479__),
    .I1(__1423__),
    .I0(__1475__),
    .O(__2026__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5710__ (
    .I5(__858__),
    .I4(__1059__),
    .I3(__944__),
    .I2(__1039__),
    .I1(__954__),
    .I0(__1052__),
    .O(__2027__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5711__ (
    .I5(__858__),
    .I4(__1096__),
    .I3(__944__),
    .I2(__1092__),
    .I1(__954__),
    .I0(__1094__),
    .O(__2028__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5712__ (
    .I5(__858__),
    .I4(__1087__),
    .I3(__944__),
    .I2(__1076__),
    .I1(__954__),
    .I0(__1082__),
    .O(__2029__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5713__ (
    .I5(__944__),
    .I4(__974__),
    .I3(__858__),
    .I2(__976__),
    .I1(__954__),
    .I0(__975__),
    .O(__2030__)
  );
  LUT6 #(
    .INIT(64'h0fff0fff88ccffff)
  ) __5714__ (
    .I5(__1810__),
    .I4(__2028__),
    .I3(__2030__),
    .I2(__2027__),
    .I1(__1809__),
    .I0(__2029__),
    .O(__2031__)
  );
  LUT6 #(
    .INIT(64'hff000e00ff00ff00)
  ) __5715__ (
    .I5(__1809__),
    .I4(__1808__),
    .I3(__2031__),
    .I2(__2029__),
    .I1(__2028__),
    .I0(__2027__),
    .O(__2032__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5716__ (
    .I5(__858__),
    .I4(__1103__),
    .I3(__944__),
    .I2(__1098__),
    .I1(__954__),
    .I0(__1100__),
    .O(__2033__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __5717__ (
    .I1(__2033__),
    .I0(__2032__),
    .O(__2034__)
  );
  LUT5 #(
    .INIT(32'h00000080)
  ) __5718__ (
    .I4(__2028__),
    .I3(__2029__),
    .I2(__1810__),
    .I1(__1808__),
    .I0(__2033__),
    .O(__2035__)
  );
  LUT6 #(
    .INIT(64'h00f000ff00ff00bb)
  ) __5719__ (
    .I5(__1810__),
    .I4(__2027__),
    .I3(__2035__),
    .I2(__1809__),
    .I1(__2033__),
    .I0(__2030__),
    .O(__2036__)
  );
  LUT6 #(
    .INIT(64'hfffffffc54fcffff)
  ) __5720__ (
    .I5(__1810__),
    .I4(__2028__),
    .I3(__2033__),
    .I2(__1809__),
    .I1(__2029__),
    .I0(__1808__),
    .O(__2037__)
  );
  LUT6 #(
    .INIT(64'h3b33000f00000000)
  ) __5721__ (
    .I5(__2029__),
    .I4(__2033__),
    .I3(__1808__),
    .I2(__2028__),
    .I1(__2030__),
    .I0(__1809__),
    .O(__2038__)
  );
  LUT3 #(
    .INIT(8'h08)
  ) __5722__ (
    .I2(__2038__),
    .I1(__2037__),
    .I0(__2036__),
    .O(__2039__)
  );
  LUT3 #(
    .INIT(8'h70)
  ) __5723__ (
    .I2(__2023__),
    .I1(__858__),
    .I0(__955__),
    .O(__2040__)
  );
  LUT6 #(
    .INIT(64'hf0f0fff3fff3ffa2)
  ) __5724__ (
    .I5(__1809__),
    .I4(__2028__),
    .I3(__1810__),
    .I2(__1808__),
    .I1(__2029__),
    .I0(__2027__),
    .O(__2041__)
  );
  LUT6 #(
    .INIT(64'h7f7f007fffffffff)
  ) __5725__ (
    .I5(__1810__),
    .I4(__1809__),
    .I3(__2028__),
    .I2(__1808__),
    .I1(__2030__),
    .I0(__2029__),
    .O(__2042__)
  );
  LUT6 #(
    .INIT(64'hfe0fffffffffffff)
  ) __5726__ (
    .I5(__1809__),
    .I4(__1808__),
    .I3(__1810__),
    .I2(__2027__),
    .I1(__2028__),
    .I0(__2033__),
    .O(__2043__)
  );
  LUT6 #(
    .INIT(64'hffffff55ffffbcfc)
  ) __5727__ (
    .I5(__2028__),
    .I4(__2029__),
    .I3(__1808__),
    .I2(__2030__),
    .I1(__2033__),
    .I0(__1810__),
    .O(__2044__)
  );
  LUT5 #(
    .INIT(32'hac000000)
  ) __5728__ (
    .I4(__2044__),
    .I3(__2043__),
    .I2(__2033__),
    .I1(__2042__),
    .I0(__2041__),
    .O(__2045__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5729__ (
    .I5(__858__),
    .I4(__1028__),
    .I3(__944__),
    .I2(__1017__),
    .I1(__954__),
    .I0(__1024__),
    .O(__2046__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5730__ (
    .I1(__954__),
    .I0(__972__),
    .O(__2047__)
  );
  LUT6 #(
    .INIT(64'h0000000000bfbfbf)
  ) __5731__ (
    .I5(__2047__),
    .I4(__944__),
    .I3(__971__),
    .I2(__1347__),
    .I1(__1033__),
    .I0(__2046__),
    .O(__2048__)
  );
  LUT6 #(
    .INIT(64'h4f440000ffcc0000)
  ) __5732__ (
    .I5(__858__),
    .I4(__1624__),
    .I3(__2048__),
    .I2(__973__),
    .I1(__2023__),
    .I0(__955__),
    .O(__2049__)
  );
  LUT6 #(
    .INIT(64'h5455555555555555)
  ) __5733__ (
    .I5(__1623__),
    .I4(__1506__),
    .I3(__1505__),
    .I2(__1508__),
    .I1(__1507__),
    .I0(__1805__),
    .O(__2050__)
  );
  LUT6 #(
    .INIT(64'hffffffffbf000000)
  ) __5734__ (
    .I5(__2050__),
    .I4(__2049__),
    .I3(__2045__),
    .I2(__2040__),
    .I1(__2039__),
    .I0(__2034__),
    .O(__2051__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __5735__ (
    .I2(__858__),
    .I1(__2051__),
    .I0(__951__),
    .O(__2052__)
  );
  LUT6 #(
    .INIT(64'hd8fad850d850d8fa)
  ) __5736__ (
    .I5(g3229),
    .I4(__1653__),
    .I3(__1651__),
    .I2(__865__),
    .I1(__1652__),
    .I0(__1812__),
    .O(__2053__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __5737__ (
    .I3(__663__),
    .I2(__603__),
    .I1(__1419__),
    .I0(__1329__),
    .O(__2054__)
  );
  LUT3 #(
    .INIT(8'h70)
  ) __5738__ (
    .I2(__1949__),
    .I1(__858__),
    .I0(__121__),
    .O(__2055__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5739__ (
    .I5(__944__),
    .I4(__107__),
    .I3(__858__),
    .I2(__109__),
    .I1(__954__),
    .I0(__108__),
    .O(__2056__)
  );
  LUT6 #(
    .INIT(64'h5455555555555555)
  ) __5740__ (
    .I5(__1623__),
    .I4(__1506__),
    .I3(__1505__),
    .I2(__1508__),
    .I1(__1507__),
    .I0(__2056__),
    .O(__2057__)
  );
  LUT6 #(
    .INIT(64'h0f080f0f0f0f0f0f)
  ) __5741__ (
    .I5(__1950__),
    .I4(__1940__),
    .I3(__1935__),
    .I2(__2057__),
    .I1(__2055__),
    .I0(__1946__),
    .O(__2058__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __5742__ (
    .I2(__954__),
    .I1(__2058__),
    .I0(__108__),
    .O(__2059__)
  );
  LUT5 #(
    .INIT(32'h21a522aa)
  ) __5743__ (
    .I4(__944__),
    .I3(__954__),
    .I2(__748__),
    .I1(__875__),
    .I0(__747__),
    .O(__2060__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __5744__ (
    .I3(__662__),
    .I2(__603__),
    .I1(__1430__),
    .I0(__1299__),
    .O(__2061__)
  );
  LUT5 #(
    .INIT(32'h80ef0000)
  ) __5745__ (
    .I4(__589__),
    .I3(__1598__),
    .I2(__1543__),
    .I1(__1544__),
    .I0(__1542__),
    .O(__2062__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5746__ (
    .I5(__589__),
    .I4(__1210__),
    .I3(__663__),
    .I2(__1212__),
    .I1(__662__),
    .I0(__1211__),
    .O(__2063__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5747__ (
    .I5(__589__),
    .I4(__1206__),
    .I3(__663__),
    .I2(__1209__),
    .I1(__662__),
    .I0(__1208__),
    .O(__2064__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5748__ (
    .I5(__589__),
    .I4(__1214__),
    .I3(__663__),
    .I2(__1219__),
    .I1(__662__),
    .I0(__1215__),
    .O(__2065__)
  );
  LUT6 #(
    .INIT(64'hd8fad850d850d8fa)
  ) __5749__ (
    .I5(g3229),
    .I4(__2065__),
    .I3(__2064__),
    .I2(__1210__),
    .I1(__2063__),
    .I0(__2062__),
    .O(__2066__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __5750__ (
    .I5(__954__),
    .I4(__242__),
    .I3(__370__),
    .I2(__229__),
    .I1(__336__),
    .I0(__216__),
    .O(__2067__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5751__ (
    .I5(__589__),
    .I4(__629__),
    .I3(__663__),
    .I2(__631__),
    .I1(__662__),
    .I0(__630__),
    .O(__2068__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5752__ (
    .I5(__589__),
    .I4(__632__),
    .I3(__663__),
    .I2(__634__),
    .I1(__662__),
    .I0(__633__),
    .O(__2069__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5753__ (
    .I5(__589__),
    .I4(__635__),
    .I3(__663__),
    .I2(__637__),
    .I1(__662__),
    .I0(__636__),
    .O(__2070__)
  );
  LUT5 #(
    .INIT(32'h80ef0000)
  ) __5754__ (
    .I4(__662__),
    .I3(__1598__),
    .I2(__1761__),
    .I1(__1760__),
    .I0(__1759__),
    .O(__2071__)
  );
  LUT6 #(
    .INIT(64'h3fffff3faaaaaaaa)
  ) __5755__ (
    .I5(__2071__),
    .I4(g3229),
    .I3(__2070__),
    .I2(__2069__),
    .I1(__2068__),
    .I0(__627__),
    .O(__2072__)
  );
  LUT5 #(
    .INIT(32'ha000cccc)
  ) __5756__ (
    .I4(__589__),
    .I3(__1761__),
    .I2(__1760__),
    .I1(__178__),
    .I0(__1759__),
    .O(__2073__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __5757__ (
    .I2(__662__),
    .I1(__1672__),
    .I0(__1000__),
    .O(__2074__)
  );
  LUT6 #(
    .INIT(64'h4000000000000000)
  ) __5758__ (
    .I5(__589__),
    .I4(__1236__),
    .I3(__1235__),
    .I2(__1237__),
    .I1(__1234__),
    .I0(__1598__),
    .O(__2075__)
  );
  LUT5 #(
    .INIT(32'h06666666)
  ) __5759__ (
    .I4(__589__),
    .I3(__1598__),
    .I2(__603__),
    .I1(__1232__),
    .I0(__2075__),
    .O(__2076__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __5760__ (
    .I2(__944__),
    .I1(__1624__),
    .I0(__1038__),
    .O(__2077__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __5761__ (
    .I5(__944__),
    .I4(__242__),
    .I3(__370__),
    .I2(__229__),
    .I1(__339__),
    .I0(__219__),
    .O(__2078__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __5762__ (
    .I5(__944__),
    .I4(__936__),
    .I3(__927__),
    .I2(__924__),
    .I1(__896__),
    .I0(__916__),
    .O(__2079__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __5763__ (
    .I3(__589__),
    .I2(__603__),
    .I1(__1448__),
    .I0(__828__),
    .O(__2080__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __5764__ (
    .I3(__662__),
    .I2(__603__),
    .I1(__1413__),
    .I0(__214__),
    .O(__2081__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __5765__ (
    .I2(__662__),
    .I1(__1598__),
    .I0(__1635__),
    .O(__2082__)
  );
  LUT6 #(
    .INIT(64'h55555d5500000800)
  ) __5766__ (
    .I5(__626__),
    .I4(__1413__),
    .I3(__1411__),
    .I2(__1412__),
    .I1(__1414__),
    .I0(__2082__),
    .O(__2083__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5767__ (
    .I5(__589__),
    .I4(__463__),
    .I3(__663__),
    .I2(__619__),
    .I1(__662__),
    .I0(__464__),
    .O(__2084__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5768__ (
    .I5(__589__),
    .I4(__549__),
    .I3(__663__),
    .I2(__551__),
    .I1(__662__),
    .I0(__550__),
    .O(__2085__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5769__ (
    .I5(__589__),
    .I4(__544__),
    .I3(__663__),
    .I2(__546__),
    .I1(__662__),
    .I0(__545__),
    .O(__2086__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5770__ (
    .I1(__1411__),
    .I0(__1414__),
    .O(__2087__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5771__ (
    .I1(__1408__),
    .I0(__1413__),
    .O(__2088__)
  );
  LUT6 #(
    .INIT(64'h8000000000000000)
  ) __5772__ (
    .I5(__1410__),
    .I4(__1409__),
    .I3(__1407__),
    .I2(__1412__),
    .I1(__2088__),
    .I0(__2087__),
    .O(__2089__)
  );
  LUT6 #(
    .INIT(64'h01f700f300ff00ff)
  ) __5773__ (
    .I5(__603__),
    .I4(__2089__),
    .I3(__1957__),
    .I2(__2086__),
    .I1(__2085__),
    .I0(__2084__),
    .O(__2090__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __5774__ (
    .I2(__663__),
    .I1(__2090__),
    .I0(__594__),
    .O(__2091__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __5775__ (
    .I5(__954__),
    .I4(__93__),
    .I3(__73__),
    .I2(__748__),
    .I1(__1393__),
    .I0(__737__),
    .O(__2092__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __5776__ (
    .I2(__944__),
    .I1(__968__),
    .I0(__752__),
    .O(__2093__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5777__ (
    .I5(__944__),
    .I4(__100__),
    .I3(__858__),
    .I2(__106__),
    .I1(__954__),
    .I0(__104__),
    .O(__2094__)
  );
  LUT6 #(
    .INIT(64'h4f0f4f0000000000)
  ) __5778__ (
    .I5(__944__),
    .I4(__2056__),
    .I3(__2094__),
    .I2(__1647__),
    .I1(__266__),
    .I0(__1951__),
    .O(__2095__)
  );
  LUT6 #(
    .INIT(64'h4eeeeeeeeeee4eee)
  ) __5779__ (
    .I5(g3229),
    .I4(__1930__),
    .I3(__1932__),
    .I2(__1928__),
    .I1(__122__),
    .I0(__2095__),
    .O(__2096__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __5780__ (
    .I3(__663__),
    .I2(__603__),
    .I1(__1428__),
    .I0(__1305__),
    .O(__2097__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5781__ (
    .I5(__858__),
    .I4(__483__),
    .I3(__944__),
    .I2(__478__),
    .I1(__954__),
    .I0(__481__),
    .O(__2098__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5782__ (
    .I5(__858__),
    .I4(__495__),
    .I3(__944__),
    .I2(__492__),
    .I1(__954__),
    .I0(__494__),
    .O(__2099__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5783__ (
    .I5(__858__),
    .I4(__490__),
    .I3(__944__),
    .I2(__511__),
    .I1(__954__),
    .I0(__488__),
    .O(__2100__)
  );
  LUT6 #(
    .INIT(64'h0fff0fff88ccffff)
  ) __5784__ (
    .I5(__1979__),
    .I4(__2099__),
    .I3(__1976__),
    .I2(__2098__),
    .I1(__1978__),
    .I0(__2100__),
    .O(__2101__)
  );
  LUT6 #(
    .INIT(64'hff000e00ff00ff00)
  ) __5785__ (
    .I5(__1978__),
    .I4(__1977__),
    .I3(__2101__),
    .I2(__2100__),
    .I1(__2099__),
    .I0(__2098__),
    .O(__2102__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5786__ (
    .I5(__858__),
    .I4(__373__),
    .I3(__944__),
    .I2(__515__),
    .I1(__954__),
    .I0(__497__),
    .O(__2103__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __5787__ (
    .I1(__2103__),
    .I0(__2102__),
    .O(__2104__)
  );
  LUT5 #(
    .INIT(32'h00000080)
  ) __5788__ (
    .I4(__2099__),
    .I3(__2100__),
    .I2(__1979__),
    .I1(__1977__),
    .I0(__2103__),
    .O(__2105__)
  );
  LUT6 #(
    .INIT(64'h00f000ff00ff00bb)
  ) __5789__ (
    .I5(__1979__),
    .I4(__2098__),
    .I3(__2105__),
    .I2(__1978__),
    .I1(__2103__),
    .I0(__1976__),
    .O(__2106__)
  );
  LUT6 #(
    .INIT(64'hfffffffc54fcffff)
  ) __5790__ (
    .I5(__1979__),
    .I4(__2099__),
    .I3(__2103__),
    .I2(__1978__),
    .I1(__2100__),
    .I0(__1977__),
    .O(__2107__)
  );
  LUT6 #(
    .INIT(64'h3b33000f00000000)
  ) __5791__ (
    .I5(__2100__),
    .I4(__2103__),
    .I3(__1977__),
    .I2(__2099__),
    .I1(__1976__),
    .I0(__1978__),
    .O(__2108__)
  );
  LUT3 #(
    .INIT(8'h08)
  ) __5792__ (
    .I2(__2108__),
    .I1(__2107__),
    .I0(__2106__),
    .O(__2109__)
  );
  LUT3 #(
    .INIT(8'h70)
  ) __5793__ (
    .I2(__1844__),
    .I1(__858__),
    .I0(__279__),
    .O(__2110__)
  );
  LUT6 #(
    .INIT(64'hf0f0fff3fff3ffa2)
  ) __5794__ (
    .I5(__1978__),
    .I4(__2099__),
    .I3(__1979__),
    .I2(__1977__),
    .I1(__2100__),
    .I0(__2098__),
    .O(__2111__)
  );
  LUT6 #(
    .INIT(64'h7f7f007fffffffff)
  ) __5795__ (
    .I5(__1979__),
    .I4(__1978__),
    .I3(__2099__),
    .I2(__1977__),
    .I1(__1976__),
    .I0(__2100__),
    .O(__2112__)
  );
  LUT6 #(
    .INIT(64'hfe0fffffffffffff)
  ) __5796__ (
    .I5(__1978__),
    .I4(__1977__),
    .I3(__1979__),
    .I2(__2098__),
    .I1(__2099__),
    .I0(__2103__),
    .O(__2113__)
  );
  LUT6 #(
    .INIT(64'hffffff55ffffbcfc)
  ) __5797__ (
    .I5(__2099__),
    .I4(__2100__),
    .I3(__1977__),
    .I2(__1976__),
    .I1(__2103__),
    .I0(__1979__),
    .O(__2114__)
  );
  LUT5 #(
    .INIT(32'hac000000)
  ) __5798__ (
    .I4(__2114__),
    .I3(__2113__),
    .I2(__2103__),
    .I1(__2112__),
    .I0(__2111__),
    .O(__2115__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5799__ (
    .I1(__954__),
    .I0(__281__),
    .O(__2116__)
  );
  LUT6 #(
    .INIT(64'h0000000000bfbfbf)
  ) __5800__ (
    .I5(__2116__),
    .I4(__944__),
    .I3(__280__),
    .I2(__252__),
    .I1(__1347__),
    .I0(__1975__),
    .O(__2117__)
  );
  LUT6 #(
    .INIT(64'h4f440000ffcc0000)
  ) __5801__ (
    .I5(__858__),
    .I4(__1624__),
    .I3(__2117__),
    .I2(__282__),
    .I1(__1844__),
    .I0(__279__),
    .O(__2118__)
  );
  LUT6 #(
    .INIT(64'h5455555555555555)
  ) __5802__ (
    .I5(__1623__),
    .I4(__1506__),
    .I3(__1505__),
    .I2(__1508__),
    .I1(__1507__),
    .I0(__1800__),
    .O(__2119__)
  );
  LUT6 #(
    .INIT(64'hffffffffbf000000)
  ) __5803__ (
    .I5(__2119__),
    .I4(__2118__),
    .I3(__2115__),
    .I2(__2110__),
    .I1(__2109__),
    .I0(__2104__),
    .O(__2120__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __5804__ (
    .I2(__858__),
    .I1(__2120__),
    .I0(__276__),
    .O(__2121__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __5805__ (
    .I3(__589__),
    .I2(__603__),
    .I1(__1457__),
    .I0(__1309__),
    .O(__2122__)
  );
  LUT4 #(
    .INIT(16'haccc)
  ) __5806__ (
    .I3(__663__),
    .I2(__603__),
    .I1(__1291__),
    .I0(__1572__),
    .O(__2123__)
  );
  LUT3 #(
    .INIT(8'h70)
  ) __5807__ (
    .I2(__2048__),
    .I1(__858__),
    .I0(__973__),
    .O(__2124__)
  );
  LUT6 #(
    .INIT(64'h5455555555555555)
  ) __5808__ (
    .I5(__1623__),
    .I4(__1506__),
    .I3(__1505__),
    .I2(__1508__),
    .I1(__1507__),
    .I0(__1674__),
    .O(__2125__)
  );
  LUT6 #(
    .INIT(64'h0f080f0f0f0f0f0f)
  ) __5809__ (
    .I5(__2049__),
    .I4(__2039__),
    .I3(__2034__),
    .I2(__2125__),
    .I1(__2124__),
    .I0(__2045__),
    .O(__2126__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __5810__ (
    .I2(__954__),
    .I1(__2126__),
    .I0(__945__),
    .O(__2127__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __5811__ (
    .I3(__663__),
    .I2(__603__),
    .I1(__1448__),
    .I0(__830__),
    .O(__2128__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __5812__ (
    .I3(__589__),
    .I2(__603__),
    .I1(__1450__),
    .I0(__824__),
    .O(__2129__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __5813__ (
    .I3(__663__),
    .I2(__603__),
    .I1(__1453__),
    .I0(__1339__),
    .O(__2130__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __5814__ (
    .I2(__1511__),
    .I1(__87__),
    .I0(__208__),
    .O(__2131__)
  );
  LUT3 #(
    .INIT(8'he2)
  ) __5815__ (
    .I2(__1427__),
    .I1(__1479__),
    .I0(__1473__),
    .O(__2132__)
  );
  LUT6 #(
    .INIT(64'h55555d5500000800)
  ) __5816__ (
    .I5(__458__),
    .I4(__1413__),
    .I3(__1411__),
    .I2(__1412__),
    .I1(__1414__),
    .I0(__1964__),
    .O(__2133__)
  );
  LUT6 #(
    .INIT(64'h4f0f4f0000000000)
  ) __5817__ (
    .I5(__944__),
    .I4(__1674__),
    .I3(__1806__),
    .I2(__1647__),
    .I1(__1036__),
    .I0(__1805__),
    .O(__2134__)
  );
  LUT6 #(
    .INIT(64'hd8fad850d850d8fa)
  ) __5818__ (
    .I5(g3229),
    .I4(__1810__),
    .I3(__1809__),
    .I2(__980__),
    .I1(__1808__),
    .I0(__2134__),
    .O(__2135__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5819__ (
    .I5(__589__),
    .I4(__526__),
    .I3(__663__),
    .I2(__528__),
    .I1(__662__),
    .I0(__527__),
    .O(__2136__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5820__ (
    .I5(__589__),
    .I4(__751__),
    .I3(__663__),
    .I2(__756__),
    .I1(__662__),
    .I0(__753__),
    .O(__2137__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5821__ (
    .I1(__1442__),
    .I0(__1440__),
    .O(__2138__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5822__ (
    .I1(__1444__),
    .I0(__1450__),
    .O(__2139__)
  );
  LUT6 #(
    .INIT(64'h8000000000000000)
  ) __5823__ (
    .I5(__1438__),
    .I4(__1448__),
    .I3(__1436__),
    .I2(__1446__),
    .I1(__2139__),
    .I0(__2138__),
    .O(__2140__)
  );
  LUT4 #(
    .INIT(16'he7ee)
  ) __5824__ (
    .I3(__2140__),
    .I2(__2137__),
    .I1(__2136__),
    .I0(__1606__),
    .O(__2141__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5825__ (
    .I5(__589__),
    .I4(__509__),
    .I3(__663__),
    .I2(__522__),
    .I1(__662__),
    .I0(__521__),
    .O(__2142__)
  );
  LUT6 #(
    .INIT(64'h108000c000000000)
  ) __5826__ (
    .I5(__603__),
    .I4(__2140__),
    .I3(__1606__),
    .I2(__2142__),
    .I1(__2136__),
    .I0(__2137__),
    .O(__2143__)
  );
  LUT5 #(
    .INIT(32'h00f4f0f0)
  ) __5827__ (
    .I4(__663__),
    .I3(__2143__),
    .I2(__522__),
    .I1(__603__),
    .I0(__2141__),
    .O(__2144__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __5828__ (
    .I2(__944__),
    .I1(__2120__),
    .I0(__274__),
    .O(__2145__)
  );
  LUT6 #(
    .INIT(64'h00000000007f0080)
  ) __5829__ (
    .I5(__1497__),
    .I4(__1491__),
    .I3(__1611__),
    .I2(__1493__),
    .I1(__1492__),
    .I0(__1494__),
    .O(__2146__)
  );
  LUT5 #(
    .INIT(32'h4ecccccc)
  ) __5830__ (
    .I4(__662__),
    .I3(__1598__),
    .I2(__1453__),
    .I1(__1263__),
    .I0(__1635__),
    .O(__2147__)
  );
  LUT6 #(
    .INIT(64'hfffffffe00000000)
  ) __5831__ (
    .I5(__589__),
    .I4(__1487__),
    .I3(__1488__),
    .I2(__1489__),
    .I1(__1490__),
    .I0(__1491__),
    .O(__2148__)
  );
  LUT6 #(
    .INIT(64'h8000000000000000)
  ) __5832__ (
    .I5(__2148__),
    .I4(__514__),
    .I3(__571__),
    .I2(__606__),
    .I1(__607__),
    .I0(__570__),
    .O(__2149__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5833__ (
    .I1(__589__),
    .I0(__603__),
    .O(__2150__)
  );
  LUT6 #(
    .INIT(64'h0000000000000010)
  ) __5834__ (
    .I5(__1487__),
    .I4(__1488__),
    .I3(__1489__),
    .I2(__2150__),
    .I1(__1490__),
    .I0(__1491__),
    .O(__2151__)
  );
  LUT5 #(
    .INIT(32'h007f0080)
  ) __5835__ (
    .I4(__604__),
    .I3(__2151__),
    .I2(__605__),
    .I1(__568__),
    .I0(__2149__),
    .O(__2152__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __5836__ (
    .I2(__1479__),
    .I1(__1473__),
    .I0(__1457__),
    .O(__2153__)
  );
  LUT5 #(
    .INIT(32'ha000cccc)
  ) __5837__ (
    .I4(__589__),
    .I3(__1597__),
    .I2(__1596__),
    .I1(__857__),
    .I0(__1595__),
    .O(__2154__)
  );
  LUT6 #(
    .INIT(64'h01f700f300ff00ff)
  ) __5838__ (
    .I5(__603__),
    .I4(__2140__),
    .I3(__1606__),
    .I2(__2142__),
    .I1(__2136__),
    .I0(__2137__),
    .O(__2155__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __5839__ (
    .I2(__662__),
    .I1(__2155__),
    .I0(__524__),
    .O(__2156__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5840__ (
    .I1(__215__),
    .I0(g3234),
    .O(__2157__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __5841__ (
    .I2(__1511__),
    .I1(__101__),
    .I0(__182__),
    .O(__2158__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __5842__ (
    .I2(__1479__),
    .I1(__1476__),
    .I0(__1454__),
    .O(__2159__)
  );
  LUT5 #(
    .INIT(32'h4ecccccc)
  ) __5843__ (
    .I4(__589__),
    .I3(__1598__),
    .I2(__1417__),
    .I1(__1280__),
    .I0(__1635__),
    .O(__2160__)
  );
  LUT4 #(
    .INIT(16'h440f)
  ) __5844__ (
    .I3(__1111__),
    .I2(__1105__),
    .I1(__1110__),
    .I0(__662__),
    .O(__2161__)
  );
  LUT6 #(
    .INIT(64'h4150c3f05050f0f0)
  ) __5845__ (
    .I5(__944__),
    .I4(__954__),
    .I3(__921__),
    .I2(__920__),
    .I1(__924__),
    .I0(__925__),
    .O(__2162__)
  );
  LUT5 #(
    .INIT(32'h77f0f0f0)
  ) __5846__ (
    .I4(__663__),
    .I3(__603__),
    .I2(__533__),
    .I1(__1731__),
    .I0(__1715__),
    .O(__2163__)
  );
  LUT5 #(
    .INIT(32'h81000000)
  ) __5847__ (
    .I4(__1761__),
    .I3(__1759__),
    .I2(__1760__),
    .I1(__1755__),
    .I0(__1735__),
    .O(__2164__)
  );
  LUT6 #(
    .INIT(64'h4000000200000000)
  ) __5848__ (
    .I5(__2164__),
    .I4(__1753__),
    .I3(__1746__),
    .I2(__1744__),
    .I1(__1737__),
    .I0(__1851__),
    .O(__2165__)
  );
  LUT6 #(
    .INIT(64'hdffffff720000008)
  ) __5849__ (
    .I5(__1750__),
    .I4(__1748__),
    .I3(__1741__),
    .I2(__1739__),
    .I1(__1851__),
    .I0(__2165__),
    .O(__2166__)
  );
  LUT6 #(
    .INIT(64'h0f0f33550f0f0f0f)
  ) __5850__ (
    .I5(__1864__),
    .I4(__1861__),
    .I3(__1857__),
    .I2(__1751__),
    .I1(__1851__),
    .I0(__2166__),
    .O(__2167__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __5851__ (
    .I2(__662__),
    .I1(__2167__),
    .I0(__661__),
    .O(__2168__)
  );
  LUT6 #(
    .INIT(64'h3fffff3faaaaaaaa)
  ) __5852__ (
    .I5(__1599__),
    .I4(g3229),
    .I3(__1602__),
    .I2(__1601__),
    .I1(__1600__),
    .I0(__1129__),
    .O(__2169__)
  );
  LUT4 #(
    .INIT(16'h25aa)
  ) __5853__ (
    .I3(__589__),
    .I2(__1598__),
    .I1(__603__),
    .I0(__607__),
    .O(__2170__)
  );
  LUT4 #(
    .INIT(16'haccc)
  ) __5854__ (
    .I3(__858__),
    .I2(__875__),
    .I1(__349__),
    .I0(__1951__),
    .O(__2171__)
  );
  LUT4 #(
    .INIT(16'h0baa)
  ) __5855__ (
    .I3(__858__),
    .I2(__1624__),
    .I1(__1844__),
    .I0(__279__),
    .O(__2172__)
  );
  LUT6 #(
    .INIT(64'h4f0f4f0000000000)
  ) __5856__ (
    .I5(__858__),
    .I4(__2056__),
    .I3(__2094__),
    .I2(__1647__),
    .I1(__266__),
    .I0(__1951__),
    .O(__2173__)
  );
  LUT6 #(
    .INIT(64'h4eeeeeeeeeee4eee)
  ) __5857__ (
    .I5(g3229),
    .I4(__1930__),
    .I3(__1932__),
    .I2(__1928__),
    .I1(__126__),
    .I0(__2173__),
    .O(__2174__)
  );
  LUT6 #(
    .INIT(64'hdffffff720000008)
  ) __5858__ (
    .I5(__1687__),
    .I4(__1692__),
    .I3(__1685__),
    .I2(__1690__),
    .I1(__1684__),
    .I0(__1960__),
    .O(__2175__)
  );
  LUT6 #(
    .INIT(64'h0f0f33550f0f0f0f)
  ) __5859__ (
    .I5(__1732__),
    .I4(__1728__),
    .I3(__1697__),
    .I2(__1712__),
    .I1(__1684__),
    .I0(__2175__),
    .O(__2176__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __5860__ (
    .I2(__589__),
    .I1(__2176__),
    .I0(__582__),
    .O(__2177__)
  );
  LUT5 #(
    .INIT(32'hf0f0ccaa)
  ) __5861__ (
    .I4(__142__),
    .I3(__858__),
    .I2(__158__),
    .I1(__1781__),
    .I0(__144__),
    .O(__2178__)
  );
  LUT3 #(
    .INIT(8'h01)
  ) __5862__ (
    .I2(__2178__),
    .I1(__140__),
    .I0(g1249),
    .O(__2179__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5863__ (
    .I5(__944__),
    .I4(__1392__),
    .I3(__858__),
    .I2(__459__),
    .I1(__954__),
    .I0(__1393__),
    .O(__2180__)
  );
  LUT6 #(
    .INIT(64'h0100000100000000)
  ) __5864__ (
    .I5(__142__),
    .I4(__2056__),
    .I3(__2180__),
    .I2(__2178__),
    .I1(__140__),
    .I0(g1249),
    .O(__2181__)
  );
  LUT3 #(
    .INIT(8'hf1)
  ) __5865__ (
    .I2(__269__),
    .I1(__93__),
    .I0(__266__),
    .O(__2182__)
  );
  LUT3 #(
    .INIT(8'hf1)
  ) __5866__ (
    .I2(__266__),
    .I1(__93__),
    .I0(__269__),
    .O(__2183__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5867__ (
    .I5(__944__),
    .I4(__1054__),
    .I3(__858__),
    .I2(__1390__),
    .I1(__954__),
    .I0(__801__),
    .O(__2184__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5868__ (
    .I5(__944__),
    .I4(__1391__),
    .I3(__858__),
    .I2(__1398__),
    .I1(__954__),
    .I0(__786__),
    .O(__2185__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5869__ (
    .I1(__2185__),
    .I0(__2184__),
    .O(__2186__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5870__ (
    .I5(__944__),
    .I4(__1399__),
    .I3(__858__),
    .I2(__1406__),
    .I1(__954__),
    .I0(__1404__),
    .O(__2187__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5871__ (
    .I5(__944__),
    .I4(__1348__),
    .I3(__858__),
    .I2(__1364__),
    .I1(__954__),
    .I0(__1343__),
    .O(__2188__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __5872__ (
    .I1(__2188__),
    .I0(__2187__),
    .O(__2189__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5873__ (
    .I5(__944__),
    .I4(__789__),
    .I3(__858__),
    .I2(__734__),
    .I1(__954__),
    .I0(__1050__),
    .O(__2190__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5874__ (
    .I5(__944__),
    .I4(__794__),
    .I3(__858__),
    .I2(__732__),
    .I1(__954__),
    .I0(__729__),
    .O(__2191__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5875__ (
    .I5(__944__),
    .I4(__1400__),
    .I3(__858__),
    .I2(__1402__),
    .I1(__954__),
    .I0(__1401__),
    .O(__2192__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5876__ (
    .I5(__944__),
    .I4(__1403__),
    .I3(__858__),
    .I2(__192__),
    .I1(__954__),
    .I0(__1421__),
    .O(__2193__)
  );
  LUT6 #(
    .INIT(64'h0000000000008000)
  ) __5877__ (
    .I5(__2193__),
    .I4(__2192__),
    .I3(__2191__),
    .I2(__2190__),
    .I1(__2189__),
    .I0(__2186__),
    .O(__2194__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5878__ (
    .I5(__944__),
    .I4(__757__),
    .I3(__858__),
    .I2(__1333__),
    .I1(__954__),
    .I0(__1332__),
    .O(__2195__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5879__ (
    .I5(__944__),
    .I4(__1042__),
    .I3(__858__),
    .I2(__1040__),
    .I1(__954__),
    .I0(__343__),
    .O(__2196__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5880__ (
    .I5(__944__),
    .I4(__1046__),
    .I3(__858__),
    .I2(__798__),
    .I1(__954__),
    .I0(__731__),
    .O(__2197__)
  );
  LUT5 #(
    .INIT(32'h00000008)
  ) __5881__ (
    .I4(__2197__),
    .I3(__2196__),
    .I2(__2195__),
    .I1(__2180__),
    .I0(__2194__),
    .O(__2198__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5882__ (
    .I5(__944__),
    .I4(__1336__),
    .I3(__858__),
    .I2(__1340__),
    .I1(__954__),
    .I0(__1338__),
    .O(__2199__)
  );
  LUT6 #(
    .INIT(64'h000000004fff0000)
  ) __5883__ (
    .I5(__266__),
    .I4(__269__),
    .I3(__142__),
    .I2(__2179__),
    .I1(__2199__),
    .I0(__2198__),
    .O(__2200__)
  );
  LUT6 #(
    .INIT(64'hffffffff000f00bb)
  ) __5884__ (
    .I5(__2200__),
    .I4(__2183__),
    .I3(__2182__),
    .I2(__2181__),
    .I1(__2179__),
    .I0(__92__),
    .O(__2201__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __5885__ (
    .I5(__764__),
    .I4(__573__),
    .I3(__858__),
    .I2(__745__),
    .I1(__704__),
    .I0(__766__),
    .O(__2202__)
  );
  LUT6 #(
    .INIT(64'haa3aaaaaaaaaaaaa)
  ) __5886__ (
    .I5(__954__),
    .I4(__93__),
    .I3(__748__),
    .I2(__73__),
    .I1(__799__),
    .I0(__1401__),
    .O(__2203__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __5887__ (
    .I3(__662__),
    .I2(__603__),
    .I1(__1407__),
    .I0(__434__),
    .O(__2204__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __5888__ (
    .I5(__954__),
    .I4(__93__),
    .I3(__73__),
    .I2(__748__),
    .I1(__343__),
    .I0(__1047__),
    .O(__2205__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __5889__ (
    .I2(__662__),
    .I1(__1962__),
    .I0(__516__),
    .O(__2206__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __5890__ (
    .I3(__663__),
    .I2(__603__),
    .I1(__1411__),
    .I0(__476__),
    .O(__2207__)
  );
  LUT3 #(
    .INIT(8'h10)
  ) __5891__ (
    .I2(__2089__),
    .I1(__1712__),
    .I0(__1705__),
    .O(__2208__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5892__ (
    .I5(__589__),
    .I4(__598__),
    .I3(__663__),
    .I2(__556__),
    .I1(__662__),
    .I0(__555__),
    .O(__2209__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5893__ (
    .I5(__589__),
    .I4(__595__),
    .I3(__663__),
    .I2(__552__),
    .I1(__662__),
    .I0(__596__),
    .O(__2210__)
  );
  LUT6 #(
    .INIT(64'hfffff888f888f888)
  ) __5894__ (
    .I5(__589__),
    .I4(__553__),
    .I3(__663__),
    .I2(__554__),
    .I1(__662__),
    .I0(__597__),
    .O(__2211__)
  );
  LUT6 #(
    .INIT(64'h000377730000ffff)
  ) __5895__ (
    .I5(__603__),
    .I4(__2211__),
    .I3(__2210__),
    .I2(__2209__),
    .I1(__2208__),
    .I0(__1710__),
    .O(__2212__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __5896__ (
    .I2(__662__),
    .I1(__2212__),
    .I0(__597__),
    .O(__2213__)
  );
  LUT6 #(
    .INIT(64'haa3aaaaaaaaaaaaa)
  ) __5897__ (
    .I5(__954__),
    .I4(__93__),
    .I3(__748__),
    .I2(__73__),
    .I1(__1051__),
    .I0(__1404__),
    .O(__2214__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __5898__ (
    .I5(__858__),
    .I4(__242__),
    .I3(__370__),
    .I2(__229__),
    .I1(__162__),
    .I0(__219__),
    .O(__2215__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __5899__ (
    .I2(__1511__),
    .I1(__95__),
    .I0(__165__),
    .O(__2216__)
  );
  LUT5 #(
    .INIT(32'h77f0f0f0)
  ) __5900__ (
    .I4(__589__),
    .I3(__603__),
    .I2(__1152__),
    .I1(__1591__),
    .I0(__1575__),
    .O(__2217__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5901__ (
    .I5(__944__),
    .I4(__884__),
    .I3(__858__),
    .I2(__886__),
    .I1(__954__),
    .I0(__885__),
    .O(__2218__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5902__ (
    .I5(__944__),
    .I4(__890__),
    .I3(__858__),
    .I2(__892__),
    .I1(__954__),
    .I0(__891__),
    .O(__2219__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5903__ (
    .I5(__944__),
    .I4(__881__),
    .I3(__858__),
    .I2(__883__),
    .I1(__954__),
    .I0(__882__),
    .O(__2220__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __5904__ (
    .I1(__2220__),
    .I0(__911__),
    .O(__2221__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5905__ (
    .I5(__944__),
    .I4(__893__),
    .I3(__858__),
    .I2(__895__),
    .I1(__954__),
    .I0(__894__),
    .O(__2222__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __5906__ (
    .I1(__915__),
    .I0(__2222__),
    .O(__2223__)
  );
  LUT6 #(
    .INIT(64'h1428000000000000)
  ) __5907__ (
    .I5(__2223__),
    .I4(__2221__),
    .I3(__2219__),
    .I2(__2218__),
    .I1(__912__),
    .I0(__914__),
    .O(__2224__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5908__ (
    .I5(__944__),
    .I4(__905__),
    .I3(__858__),
    .I2(__907__),
    .I1(__954__),
    .I0(__906__),
    .O(__2225__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5909__ (
    .I5(__944__),
    .I4(__896__),
    .I3(__858__),
    .I2(__898__),
    .I1(__954__),
    .I0(__897__),
    .O(__2226__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5910__ (
    .I1(__2226__),
    .I0(__916__),
    .O(__2227__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5911__ (
    .I5(__944__),
    .I4(__902__),
    .I3(__858__),
    .I2(__904__),
    .I1(__954__),
    .I0(__903__),
    .O(__2228__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __5912__ (
    .I1(__2226__),
    .I0(__916__),
    .O(__2229__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5913__ (
    .I5(__944__),
    .I4(__887__),
    .I3(__858__),
    .I2(__889__),
    .I1(__954__),
    .I0(__888__),
    .O(__2230__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __5914__ (
    .I1(__2230__),
    .I0(__913__),
    .O(__2231__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5915__ (
    .I5(__944__),
    .I4(__908__),
    .I3(__858__),
    .I2(__910__),
    .I1(__954__),
    .I0(__909__),
    .O(__2232__)
  );
  LUT4 #(
    .INIT(16'h7770)
  ) __5916__ (
    .I3(__2225__),
    .I2(__920__),
    .I1(__2230__),
    .I0(__913__),
    .O(__2233__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5917__ (
    .I5(__944__),
    .I4(__899__),
    .I3(__858__),
    .I2(__901__),
    .I1(__954__),
    .I0(__900__),
    .O(__2234__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __5918__ (
    .I1(__2234__),
    .I0(__917__),
    .O(__2235__)
  );
  LUT6 #(
    .INIT(64'h0110000000000000)
  ) __5919__ (
    .I5(__2235__),
    .I4(__2233__),
    .I3(__2232__),
    .I2(__921__),
    .I1(__2231__),
    .I0(__2229__),
    .O(__2236__)
  );
  LUT6 #(
    .INIT(64'h0007070000000000)
  ) __5920__ (
    .I5(__2236__),
    .I4(__918__),
    .I3(__2228__),
    .I2(__2227__),
    .I1(__2225__),
    .I0(__920__),
    .O(__2237__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5921__ (
    .I1(__944__),
    .I0(__878__),
    .O(__2238__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5922__ (
    .I5(__944__),
    .I4(__874__),
    .I3(__858__),
    .I2(__877__),
    .I1(__954__),
    .I0(__876__),
    .O(__2239__)
  );
  LUT6 #(
    .INIT(64'h00008acf00000000)
  ) __5923__ (
    .I5(__2239__),
    .I4(__2238__),
    .I3(__858__),
    .I2(__954__),
    .I1(__879__),
    .I0(__880__),
    .O(__2240__)
  );
  LUT4 #(
    .INIT(16'h0080)
  ) __5924__ (
    .I3(__924__),
    .I2(__944__),
    .I1(__936__),
    .I0(__927__),
    .O(__2241__)
  );
  LUT5 #(
    .INIT(32'h3f00aaaa)
  ) __5925__ (
    .I4(__2241__),
    .I3(__2240__),
    .I2(__2237__),
    .I1(__2224__),
    .I0(__856__),
    .O(__2242__)
  );
  LUT4 #(
    .INIT(16'haccc)
  ) __5926__ (
    .I3(__662__),
    .I2(__603__),
    .I1(__1290__),
    .I0(__1572__),
    .O(__2243__)
  );
  LUT6 #(
    .INIT(64'h4f0f4f0000000000)
  ) __5927__ (
    .I5(__858__),
    .I4(__1982__),
    .I3(__1981__),
    .I2(__1647__),
    .I1(__354__),
    .I0(__1800__),
    .O(__2244__)
  );
  LUT6 #(
    .INIT(64'h3fffff3faaaaaaaa)
  ) __5928__ (
    .I5(__2244__),
    .I4(g3229),
    .I3(__1979__),
    .I2(__1978__),
    .I1(__1977__),
    .I0(__286__),
    .O(__2245__)
  );
  LUT3 #(
    .INIT(8'h10)
  ) __5929__ (
    .I2(__1617__),
    .I1(__1884__),
    .I0(__1893__),
    .O(__2246__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5930__ (
    .I5(__589__),
    .I4(__1120__),
    .I3(__663__),
    .I2(__1123__),
    .I1(__662__),
    .I0(__1122__),
    .O(__2247__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5931__ (
    .I5(__589__),
    .I4(__1126__),
    .I3(__663__),
    .I2(__1128__),
    .I1(__662__),
    .I0(__1127__),
    .O(__2248__)
  );
  LUT6 #(
    .INIT(64'hfffff888f888f888)
  ) __5932__ (
    .I5(__589__),
    .I4(__1108__),
    .I3(__663__),
    .I2(__1125__),
    .I1(__662__),
    .I0(__1124__),
    .O(__2249__)
  );
  LUT6 #(
    .INIT(64'h000377730000ffff)
  ) __5933__ (
    .I5(__603__),
    .I4(__2249__),
    .I3(__2248__),
    .I2(__2247__),
    .I1(__2246__),
    .I0(__1899__),
    .O(__2250__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __5934__ (
    .I2(__589__),
    .I1(__2250__),
    .I0(__1108__),
    .O(__2251__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __5935__ (
    .I3(__662__),
    .I2(__603__),
    .I1(__1440__),
    .I0(__841__),
    .O(__2252__)
  );
  LUT6 #(
    .INIT(64'h4150c3f05050f0f0)
  ) __5936__ (
    .I5(__944__),
    .I4(__954__),
    .I3(__760__),
    .I2(__768__),
    .I1(__745__),
    .I0(__752__),
    .O(__2253__)
  );
  LUT5 #(
    .INIT(32'h0030aaaa)
  ) __5937__ (
    .I4(__663__),
    .I3(__1682__),
    .I2(__1681__),
    .I1(__1680__),
    .I0(__380__),
    .O(__2254__)
  );
  LUT4 #(
    .INIT(16'hf8ff)
  ) __5938__ (
    .I3(__603__),
    .I2(__1710__),
    .I1(__1725__),
    .I0(__1720__),
    .O(__2255__)
  );
  LUT5 #(
    .INIT(32'h80000000)
  ) __5939__ (
    .I4(__1714__),
    .I3(__1709__),
    .I2(__1704__),
    .I1(__1701__),
    .I0(__2255__),
    .O(__2256__)
  );
  LUT6 #(
    .INIT(64'h4000000000000000)
  ) __5940__ (
    .I5(__1681__),
    .I4(__1714__),
    .I3(__1709__),
    .I2(__1704__),
    .I1(__1701__),
    .I0(__1680__),
    .O(__2257__)
  );
  LUT4 #(
    .INIT(16'h1428)
  ) __5941__ (
    .I3(__1409__),
    .I2(__1407__),
    .I1(__1677__),
    .I0(__1678__),
    .O(__2258__)
  );
  LUT4 #(
    .INIT(16'h0990)
  ) __5942__ (
    .I3(__1414__),
    .I2(__1692__),
    .I1(__1712__),
    .I0(__1687__),
    .O(__2259__)
  );
  LUT4 #(
    .INIT(16'h1428)
  ) __5943__ (
    .I3(__1408__),
    .I2(__1410__),
    .I1(__1686__),
    .I0(__1679__),
    .O(__2260__)
  );
  LUT4 #(
    .INIT(16'h0990)
  ) __5944__ (
    .I3(__1413__),
    .I2(__1690__),
    .I1(__1705__),
    .I0(__1685__),
    .O(__2261__)
  );
  LUT6 #(
    .INIT(64'h8000000000000000)
  ) __5945__ (
    .I5(__1721__),
    .I4(__1717__),
    .I3(__2261__),
    .I2(__2260__),
    .I1(__2259__),
    .I0(__2258__),
    .O(__2262__)
  );
  LUT3 #(
    .INIT(8'h10)
  ) __5946__ (
    .I2(__1681__),
    .I1(__1682__),
    .I0(__1680__),
    .O(__2263__)
  );
  LUT5 #(
    .INIT(32'hcd000000)
  ) __5947__ (
    .I4(__662__),
    .I3(__603__),
    .I2(__1710__),
    .I1(__2263__),
    .I0(__2262__),
    .O(__2264__)
  );
  LUT6 #(
    .INIT(64'hffff0707ff00ff00)
  ) __5948__ (
    .I5(__2264__),
    .I4(__1682__),
    .I3(__541__),
    .I2(__2257__),
    .I1(__1680__),
    .I0(__2256__),
    .O(__2265__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __5949__ (
    .I5(__954__),
    .I4(__936__),
    .I3(__927__),
    .I2(__924__),
    .I1(__897__),
    .I0(__916__),
    .O(__2266__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __5950__ (
    .I2(__858__),
    .I1(__300__),
    .I0(__1359__),
    .O(__2267__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __5951__ (
    .I3(__663__),
    .I2(__603__),
    .I1(__1422__),
    .I0(__1321__),
    .O(__2268__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5952__ (
    .I5(__944__),
    .I4(__816__),
    .I3(__858__),
    .I2(__818__),
    .I1(__954__),
    .I0(__566__),
    .O(__2269__)
  );
  LUT6 #(
    .INIT(64'he4ee4e4e4eeee4e4)
  ) __5953__ (
    .I5(g3229),
    .I4(__1652__),
    .I3(__2269__),
    .I2(__1653__),
    .I1(__863__),
    .I0(__1812__),
    .O(__2270__)
  );
  LUT5 #(
    .INIT(32'hdff72008)
  ) __5954__ (
    .I4(__1741__),
    .I3(__1748__),
    .I2(__1739__),
    .I1(__1851__),
    .I0(__2165__),
    .O(__2271__)
  );
  LUT6 #(
    .INIT(64'h0f0f33550f0f0f0f)
  ) __5955__ (
    .I5(__1864__),
    .I4(__1861__),
    .I3(__1857__),
    .I2(__1742__),
    .I1(__1851__),
    .I0(__2271__),
    .O(__2272__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __5956__ (
    .I2(__663__),
    .I1(__2272__),
    .I0(__699__),
    .O(__2273__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __5957__ (
    .I5(__764__),
    .I4(__573__),
    .I3(__954__),
    .I2(__745__),
    .I1(__664__),
    .I0(__767__),
    .O(__2274__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __5958__ (
    .I3(__663__),
    .I2(__603__),
    .I1(__1407__),
    .I0(__456__),
    .O(__2275__)
  );
  LUT3 #(
    .INIT(8'h10)
  ) __5959__ (
    .I2(__2140__),
    .I1(__1751__),
    .I0(__1742__),
    .O(__2276__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5960__ (
    .I5(__589__),
    .I4(__615__),
    .I3(__663__),
    .I2(__624__),
    .I1(__662__),
    .I0(__621__),
    .O(__2277__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5961__ (
    .I5(__589__),
    .I4(__529__),
    .I3(__663__),
    .I2(__539__),
    .I1(__662__),
    .I0(__537__),
    .O(__2278__)
  );
  LUT6 #(
    .INIT(64'hfffff888f888f888)
  ) __5962__ (
    .I5(__589__),
    .I4(__540__),
    .I3(__663__),
    .I2(__608__),
    .I1(__662__),
    .I0(__542__),
    .O(__2279__)
  );
  LUT6 #(
    .INIT(64'h000377730000ffff)
  ) __5963__ (
    .I5(__603__),
    .I4(__2279__),
    .I3(__2278__),
    .I2(__2277__),
    .I1(__2276__),
    .I0(__1757__),
    .O(__2280__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __5964__ (
    .I2(__662__),
    .I1(__2280__),
    .I0(__542__),
    .O(__2281__)
  );
  LUT6 #(
    .INIT(64'h0000000000000010)
  ) __5965__ (
    .I5(__1487__),
    .I4(__1488__),
    .I3(__1489__),
    .I2(__1635__),
    .I1(__1490__),
    .I0(__1491__),
    .O(__2282__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __5966__ (
    .I3(__663__),
    .I2(__2282__),
    .I1(__2089__),
    .I0(__619__),
    .O(__2283__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __5967__ (
    .I5(__858__),
    .I4(__936__),
    .I3(__927__),
    .I2(__924__),
    .I1(__901__),
    .I0(__917__),
    .O(__2284__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5968__ (
    .I5(__589__),
    .I4(__211__),
    .I3(__663__),
    .I2(__602__),
    .I1(__662__),
    .I0(__560__),
    .O(__2285__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5969__ (
    .I5(__589__),
    .I4(__558__),
    .I3(__663__),
    .I2(__559__),
    .I1(__662__),
    .I0(__601__),
    .O(__2286__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5970__ (
    .I5(__589__),
    .I4(__578__),
    .I3(__663__),
    .I2(__563__),
    .I1(__662__),
    .I0(__562__),
    .O(__2287__)
  );
  LUT5 #(
    .INIT(32'h80ef0000)
  ) __5971__ (
    .I4(__663__),
    .I3(__1598__),
    .I2(__1682__),
    .I1(__1681__),
    .I0(__1680__),
    .O(__2288__)
  );
  LUT6 #(
    .INIT(64'h3fffff3faaaaaaaa)
  ) __5972__ (
    .I5(__2288__),
    .I4(g3229),
    .I3(__2287__),
    .I2(__2286__),
    .I1(__2285__),
    .I0(__600__),
    .O(__2289__)
  );
  LUT6 #(
    .INIT(64'h5555cffc55555555)
  ) __5973__ (
    .I5(__1732__),
    .I4(__1728__),
    .I3(__1690__),
    .I2(__1960__),
    .I1(__1697__),
    .I0(__1413__),
    .O(__2290__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __5974__ (
    .I2(__589__),
    .I1(__2290__),
    .I0(__576__),
    .O(__2291__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5975__ (
    .I5(__944__),
    .I4(__436__),
    .I3(__858__),
    .I2(__429__),
    .I1(__954__),
    .I0(__424__),
    .O(__2292__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __5976__ (
    .I5(__944__),
    .I4(__184__),
    .I3(__858__),
    .I2(__183__),
    .I1(__954__),
    .I0(__185__),
    .O(__2293__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __5977__ (
    .I5(__954__),
    .I4(__93__),
    .I3(__73__),
    .I2(__748__),
    .I1(__731__),
    .I0(__797__),
    .O(__2294__)
  );
  LUT6 #(
    .INIT(64'hd8fad850d850d8fa)
  ) __5978__ (
    .I5(g3229),
    .I4(__2070__),
    .I3(__2068__),
    .I2(__633__),
    .I1(__2069__),
    .I0(__2071__),
    .O(__2295__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __5979__ (
    .I2(__663__),
    .I1(__2280__),
    .I0(__608__),
    .O(__2296__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __5980__ (
    .I3(__589__),
    .I2(__603__),
    .I1(__1417__),
    .I0(__1334__),
    .O(__2297__)
  );
  LUT6 #(
    .INIT(64'h0000baaaaaaaaaaa)
  ) __5981__ (
    .I5(__858__),
    .I4(__875__),
    .I3(__93__),
    .I2(__73__),
    .I1(__748__),
    .I0(__1333__),
    .O(__2298__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __5982__ (
    .I3(__589__),
    .I2(__2282__),
    .I1(__1407__),
    .I0(__622__),
    .O(__2299__)
  );
  LUT4 #(
    .INIT(16'haccc)
  ) __5983__ (
    .I3(__589__),
    .I2(__603__),
    .I1(__820__),
    .I0(__1742__),
    .O(__2300__)
  );
  LUT5 #(
    .INIT(32'h0030aaaa)
  ) __5984__ (
    .I4(__589__),
    .I3(__1681__),
    .I2(__1682__),
    .I1(__1680__),
    .I0(__482__),
    .O(__2301__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __5985__ (
    .I5(__944__),
    .I4(__242__),
    .I3(__370__),
    .I2(__229__),
    .I1(__194__),
    .I0(__225__),
    .O(__2302__)
  );
  LUT6 #(
    .INIT(64'h4545ff000505ff00)
  ) __5986__ (
    .I5(__858__),
    .I4(__954__),
    .I3(__953__),
    .I2(__2023__),
    .I1(__955__),
    .I0(__1624__),
    .O(__2303__)
  );
  LUT6 #(
    .INIT(64'h00f07878f0f0f0f0)
  ) __5987__ (
    .I5(__589__),
    .I4(__1598__),
    .I3(__603__),
    .I2(__1176__),
    .I1(__1178__),
    .I0(__1180__),
    .O(__2304__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __5988__ (
    .I3(__662__),
    .I2(__603__),
    .I1(__1422__),
    .I0(__1320__),
    .O(__2305__)
  );
  LUT6 #(
    .INIT(64'h0100000100000000)
  ) __5989__ (
    .I5(__142__),
    .I4(__2191__),
    .I3(__1951__),
    .I2(__2178__),
    .I1(__140__),
    .I0(g1249),
    .O(__2306__)
  );
  LUT6 #(
    .INIT(64'h0000df0f00000000)
  ) __5990__ (
    .I5(__269__),
    .I4(__266__),
    .I3(__142__),
    .I2(__2179__),
    .I1(__2198__),
    .I0(__2199__),
    .O(__2307__)
  );
  LUT6 #(
    .INIT(64'hffffffff000f00bb)
  ) __5991__ (
    .I5(__2307__),
    .I4(__2183__),
    .I3(__2182__),
    .I2(__2306__),
    .I1(__2179__),
    .I0(__91__),
    .O(__2308__)
  );
  LUT3 #(
    .INIT(8'he2)
  ) __5992__ (
    .I2(__1425__),
    .I1(__1479__),
    .I0(__1474__),
    .O(__2309__)
  );
  LUT4 #(
    .INIT(16'haccc)
  ) __5993__ (
    .I3(__858__),
    .I2(__752__),
    .I1(__675__),
    .I0(__1649__),
    .O(__2310__)
  );
  LUT6 #(
    .INIT(64'h00007fff00008000)
  ) __5994__ (
    .I5(__1223__),
    .I4(__2151__),
    .I3(__1228__),
    .I2(__1232__),
    .I1(__2075__),
    .I0(__1224__),
    .O(__2311__)
  );
  LUT5 #(
    .INIT(32'h80000000)
  ) __5995__ (
    .I4(__1776__),
    .I3(__1773__),
    .I2(__1769__),
    .I1(__1766__),
    .I0(__1758__),
    .O(__2312__)
  );
  LUT6 #(
    .INIT(64'h4000000000000000)
  ) __5996__ (
    .I5(__1776__),
    .I4(__1773__),
    .I3(__1769__),
    .I2(__1766__),
    .I1(__1760__),
    .I0(__1759__),
    .O(__2313__)
  );
  LUT3 #(
    .INIT(8'h10)
  ) __5997__ (
    .I2(__1760__),
    .I1(__1761__),
    .I0(__1759__),
    .O(__2314__)
  );
  LUT5 #(
    .INIT(32'hcd000000)
  ) __5998__ (
    .I4(__589__),
    .I3(__603__),
    .I2(__1757__),
    .I1(__2314__),
    .I0(__1997__),
    .O(__2315__)
  );
  LUT6 #(
    .INIT(64'hffff0707ff00ff00)
  ) __5999__ (
    .I5(__2315__),
    .I4(__1761__),
    .I3(__407__),
    .I2(__2313__),
    .I1(__1759__),
    .I0(__2312__),
    .O(__2316__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6000__ (
    .I1(__1486__),
    .I0(__1611__),
    .O(__2317__)
  );
  LUT5 #(
    .INIT(32'h13132020)
  ) __6001__ (
    .I4(__1484__),
    .I3(__1483__),
    .I2(__1485__),
    .I1(__1497__),
    .I0(__2317__),
    .O(__2318__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6002__ (
    .I1(__954__),
    .I0(__925__),
    .O(__2319__)
  );
  LUT6 #(
    .INIT(64'h00007fff00008000)
  ) __6003__ (
    .I5(__913__),
    .I4(__2319__),
    .I3(__915__),
    .I2(__916__),
    .I1(__914__),
    .I0(__1868__),
    .O(__2320__)
  );
  LUT6 #(
    .INIT(64'h0f005555cccccccc)
  ) __6004__ (
    .I5(__589__),
    .I4(__603__),
    .I3(__2089__),
    .I2(__2084__),
    .I1(__549__),
    .I0(__2085__),
    .O(__2321__)
  );
  LUT6 #(
    .INIT(64'haa3aaaaaaaaaaaaa)
  ) __6005__ (
    .I5(__944__),
    .I4(__93__),
    .I3(__748__),
    .I2(__73__),
    .I1(__799__),
    .I0(__1400__),
    .O(__2322__)
  );
  LUT4 #(
    .INIT(16'haccc)
  ) __6006__ (
    .I3(__954__),
    .I2(__231__),
    .I1(__310__),
    .I0(__1800__),
    .O(__2323__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6007__ (
    .I2(__944__),
    .I1(__1647__),
    .I0(__229__),
    .O(__2324__)
  );
  LUT6 #(
    .INIT(64'h8000010000000000)
  ) __6008__ (
    .I5(__1597__),
    .I4(__1596__),
    .I3(__1595__),
    .I2(__1897__),
    .I1(__1886__),
    .I0(__1877__),
    .O(__2325__)
  );
  LUT6 #(
    .INIT(64'h9393399393939393)
  ) __6009__ (
    .I5(__1597__),
    .I4(__1596__),
    .I3(__1595__),
    .I2(__1895__),
    .I1(__1879__),
    .I0(__2325__),
    .O(__2326__)
  );
  LUT5 #(
    .INIT(32'h0fbb0f0f)
  ) __6010__ (
    .I4(__2015__),
    .I3(__2012__),
    .I2(__1457__),
    .I1(__2326__),
    .I0(__2008__),
    .O(__2327__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __6011__ (
    .I2(__589__),
    .I1(__2327__),
    .I0(__1213__),
    .O(__2328__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __6012__ (
    .I3(__662__),
    .I2(__603__),
    .I1(__1448__),
    .I0(__829__),
    .O(__2329__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __6013__ (
    .I5(__764__),
    .I4(__573__),
    .I3(__954__),
    .I2(__745__),
    .I1(__683__),
    .I0(__770__),
    .O(__2330__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6014__ (
    .I2(__662__),
    .I1(__2176__),
    .I0(__572__),
    .O(__2331__)
  );
  LUT4 #(
    .INIT(16'haccc)
  ) __6015__ (
    .I3(__944__),
    .I2(__925__),
    .I1(__874__),
    .I0(__1674__),
    .O(__2332__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __6016__ (
    .I1(__1514__),
    .I0(__1513__),
    .O(__2333__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __6017__ (
    .I1(__1512__),
    .I0(__1515__),
    .O(__2334__)
  );
  LUT6 #(
    .INIT(64'h6996966996696996)
  ) __6018__ (
    .I5(__1516__),
    .I4(__1517__),
    .I3(__1519__),
    .I2(__1518__),
    .I1(__2334__),
    .I0(__2333__),
    .O(__2335__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __6019__ (
    .I1(__2335__),
    .I0(__1520__),
    .O(__2336__)
  );
  LUT5 #(
    .INIT(32'hafbfbaaa)
  ) __6020__ (
    .I4(__1499__),
    .I3(__1498__),
    .I2(__215__),
    .I1(__1623__),
    .I0(g3234),
    .O(__2337__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __6021__ (
    .I2(__662__),
    .I1(__1657__),
    .I0(__1249__),
    .O(__2338__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __6022__ (
    .I3(__589__),
    .I2(__603__),
    .I1(__1412__),
    .I0(__340__),
    .O(__2339__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __6023__ (
    .I5(__954__),
    .I4(__936__),
    .I3(__927__),
    .I2(__924__),
    .I1(__891__),
    .I0(__914__),
    .O(__2340__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __6024__ (
    .I5(__944__),
    .I4(__667__),
    .I3(__858__),
    .I2(__669__),
    .I1(__954__),
    .I0(__668__),
    .O(__2341__)
  );
  LUT6 #(
    .INIT(64'h0100000000000000)
  ) __6025__ (
    .I5(__1817__),
    .I4(__1828__),
    .I3(__1830__),
    .I2(__1826__),
    .I1(__2341__),
    .I0(__1823__),
    .O(__2342__)
  );
  LUT6 #(
    .INIT(64'h0000000000000008)
  ) __6026__ (
    .I5(__1837__),
    .I4(__1816__),
    .I3(__1818__),
    .I2(__1832__),
    .I1(__1824__),
    .I0(__1820__),
    .O(__2343__)
  );
  LUT5 #(
    .INIT(32'h00000010)
  ) __6027__ (
    .I4(__862__),
    .I3(__1782__),
    .I2(__868__),
    .I1(g1943),
    .I0(__867__),
    .O(__2344__)
  );
  LUT5 #(
    .INIT(32'hf8070000)
  ) __6028__ (
    .I4(__2344__),
    .I3(__1646__),
    .I2(__1826__),
    .I1(__2343__),
    .I0(__2342__),
    .O(__2345__)
  );
  LUT5 #(
    .INIT(32'h00000007)
  ) __6029__ (
    .I4(__1782__),
    .I3(g1943),
    .I2(__867__),
    .I1(__862__),
    .I0(__868__),
    .O(__2346__)
  );
  LUT3 #(
    .INIT(8'hf1)
  ) __6030__ (
    .I2(__969__),
    .I1(__764__),
    .I0(__968__),
    .O(__2347__)
  );
  LUT3 #(
    .INIT(8'hf1)
  ) __6031__ (
    .I2(__968__),
    .I1(__764__),
    .I0(__969__),
    .O(__2348__)
  );
  LUT5 #(
    .INIT(32'h00330fab)
  ) __6032__ (
    .I4(__2348__),
    .I3(__2347__),
    .I2(__2346__),
    .I1(__2345__),
    .I0(__769__),
    .O(__2349__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __6033__ (
    .I3(__663__),
    .I2(__2282__),
    .I1(__1438__),
    .I0(__780__),
    .O(__2350__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __6034__ (
    .I3(__589__),
    .I2(__603__),
    .I1(__1432__),
    .I0(__1295__),
    .O(__2351__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __6035__ (
    .I2(__944__),
    .I1(__2058__),
    .I0(__107__),
    .O(__2352__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6036__ (
    .I2(__1479__),
    .I1(__1449__),
    .I0(__1462__),
    .O(__2353__)
  );
  LUT6 #(
    .INIT(64'h7878d27878787878)
  ) __6037__ (
    .I5(__1761__),
    .I4(__1760__),
    .I3(__1759__),
    .I2(__1748__),
    .I1(__1739__),
    .I0(__2165__),
    .O(__2354__)
  );
  LUT5 #(
    .INIT(32'hf011f0f0)
  ) __6038__ (
    .I4(__1864__),
    .I3(__1861__),
    .I2(__1450__),
    .I1(__1857__),
    .I0(__2354__),
    .O(__2355__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6039__ (
    .I2(__662__),
    .I1(__2355__),
    .I0(__703__),
    .O(__2356__)
  );
  LUT6 #(
    .INIT(64'h5555cffc55555555)
  ) __6040__ (
    .I5(__1864__),
    .I4(__1861__),
    .I3(__1739__),
    .I2(__2165__),
    .I1(__1857__),
    .I0(__1448__),
    .O(__2357__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __6041__ (
    .I2(__589__),
    .I1(__2357__),
    .I0(__708__),
    .O(__2358__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6042__ (
    .I2(__1479__),
    .I1(__1472__),
    .I0(__1458__),
    .O(__2359__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6043__ (
    .I2(__1479__),
    .I1(__1439__),
    .I0(__1467__),
    .O(__2360__)
  );
  LUT5 #(
    .INIT(32'h81000000)
  ) __6044__ (
    .I4(__1597__),
    .I3(__1595__),
    .I2(__1596__),
    .I1(__1897__),
    .I0(__1877__),
    .O(__2361__)
  );
  LUT6 #(
    .INIT(64'h4000000200000000)
  ) __6045__ (
    .I5(__2361__),
    .I4(__1895__),
    .I3(__1888__),
    .I2(__1886__),
    .I1(__1879__),
    .I0(__2002__),
    .O(__2362__)
  );
  LUT6 #(
    .INIT(64'hdffffff720000008)
  ) __6046__ (
    .I5(__1892__),
    .I4(__1890__),
    .I3(__1883__),
    .I2(__1881__),
    .I1(__2002__),
    .I0(__2362__),
    .O(__2363__)
  );
  LUT6 #(
    .INIT(64'h0f0f33550f0f0f0f)
  ) __6047__ (
    .I5(__2015__),
    .I4(__2012__),
    .I3(__2008__),
    .I2(__1893__),
    .I1(__2002__),
    .I0(__2363__),
    .O(__2364__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6048__ (
    .I2(__589__),
    .I1(__2364__),
    .I0(__1182__),
    .O(__2365__)
  );
  LUT6 #(
    .INIT(64'h9333363333333333)
  ) __6049__ (
    .I5(__1761__),
    .I4(__1760__),
    .I3(__1759__),
    .I2(__1755__),
    .I1(__1744__),
    .I0(__1735__),
    .O(__2366__)
  );
  LUT6 #(
    .INIT(64'hf0f033aaf0f0f0f0)
  ) __6050__ (
    .I5(__1864__),
    .I4(__1861__),
    .I3(__1857__),
    .I2(__1440__),
    .I1(__1851__),
    .I0(__2366__),
    .O(__2367__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6051__ (
    .I2(__663__),
    .I1(__2367__),
    .I0(__722__),
    .O(__2368__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __6052__ (
    .I5(__589__),
    .I4(__557__),
    .I3(__663__),
    .I2(__600__),
    .I1(__662__),
    .I0(__599__),
    .O(__2369__)
  );
  LUT5 #(
    .INIT(32'h80ef0000)
  ) __6053__ (
    .I4(__589__),
    .I3(__1598__),
    .I2(__1682__),
    .I1(__1681__),
    .I0(__1680__),
    .O(__2370__)
  );
  LUT6 #(
    .INIT(64'hcc77f0f077ccf0f0)
  ) __6054__ (
    .I5(g3229),
    .I4(__2370__),
    .I3(__2287__),
    .I2(__558__),
    .I1(__2285__),
    .I0(__2369__),
    .O(__2371__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __6055__ (
    .I2(__1164__),
    .I1(__1174__),
    .I0(__1874__),
    .O(__2372__)
  );
  LUT6 #(
    .INIT(64'h00007fff00008000)
  ) __6056__ (
    .I5(__1043__),
    .I4(__2151__),
    .I3(__1048__),
    .I2(__730__),
    .I1(__1161__),
    .I0(__2372__),
    .O(__2373__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __6057__ (
    .I5(__858__),
    .I4(__253__),
    .I3(__944__),
    .I2(__462__),
    .I1(__954__),
    .I0(__620__),
    .O(__2374__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __6058__ (
    .I5(__858__),
    .I4(__569__),
    .I3(__944__),
    .I2(__1019__),
    .I1(__954__),
    .I0(__588__),
    .O(__2375__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __6059__ (
    .I5(__858__),
    .I4(__650__),
    .I3(__944__),
    .I2(__733__),
    .I1(__954__),
    .I0(__923__),
    .O(__2376__)
  );
  LUT6 #(
    .INIT(64'h0fff0fff88ccffff)
  ) __6060__ (
    .I5(__1653__),
    .I4(__2375__),
    .I3(__2269__),
    .I2(__2374__),
    .I1(__1651__),
    .I0(__2376__),
    .O(__2377__)
  );
  LUT6 #(
    .INIT(64'hff000e00ff00ff00)
  ) __6061__ (
    .I5(__1651__),
    .I4(__1652__),
    .I3(__2377__),
    .I2(__2376__),
    .I1(__2375__),
    .I0(__2374__),
    .O(__2378__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __6062__ (
    .I5(__858__),
    .I4(__773__),
    .I3(__944__),
    .I2(__1030__),
    .I1(__954__),
    .I0(__1031__),
    .O(__2379__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __6063__ (
    .I1(__2379__),
    .I0(__2378__),
    .O(__2380__)
  );
  LUT5 #(
    .INIT(32'h00000080)
  ) __6064__ (
    .I4(__2375__),
    .I3(__2376__),
    .I2(__1652__),
    .I1(__2379__),
    .I0(__1653__),
    .O(__2381__)
  );
  LUT6 #(
    .INIT(64'h00f000ff00ff00bb)
  ) __6065__ (
    .I5(__1653__),
    .I4(__2374__),
    .I3(__2381__),
    .I2(__1651__),
    .I1(__2379__),
    .I0(__2269__),
    .O(__2382__)
  );
  LUT6 #(
    .INIT(64'hfffffffc54fcffff)
  ) __6066__ (
    .I5(__1653__),
    .I4(__2375__),
    .I3(__2379__),
    .I2(__2376__),
    .I1(__1651__),
    .I0(__1652__),
    .O(__2383__)
  );
  LUT6 #(
    .INIT(64'h3b33000f00000000)
  ) __6067__ (
    .I5(__2376__),
    .I4(__2379__),
    .I3(__1652__),
    .I2(__2375__),
    .I1(__2269__),
    .I0(__1651__),
    .O(__2384__)
  );
  LUT3 #(
    .INIT(8'h08)
  ) __6068__ (
    .I2(__2384__),
    .I1(__2383__),
    .I0(__2382__),
    .O(__2385__)
  );
  LUT3 #(
    .INIT(8'h70)
  ) __6069__ (
    .I2(__1665__),
    .I1(__858__),
    .I0(__812__),
    .O(__2386__)
  );
  LUT6 #(
    .INIT(64'hf0f0fff3fff3ffa2)
  ) __6070__ (
    .I5(__2375__),
    .I4(__1651__),
    .I3(__1653__),
    .I2(__1652__),
    .I1(__2376__),
    .I0(__2374__),
    .O(__2387__)
  );
  LUT6 #(
    .INIT(64'h7f7f007fffffffff)
  ) __6071__ (
    .I5(__1653__),
    .I4(__1651__),
    .I3(__2375__),
    .I2(__2376__),
    .I1(__1652__),
    .I0(__2269__),
    .O(__2388__)
  );
  LUT6 #(
    .INIT(64'hfe0fffffffffffff)
  ) __6072__ (
    .I5(__1652__),
    .I4(__1651__),
    .I3(__1653__),
    .I2(__2374__),
    .I1(__2375__),
    .I0(__2379__),
    .O(__2389__)
  );
  LUT6 #(
    .INIT(64'hffffff55ffffbcfc)
  ) __6073__ (
    .I5(__2375__),
    .I4(__2376__),
    .I3(__1652__),
    .I2(__2379__),
    .I1(__2269__),
    .I0(__1653__),
    .O(__2390__)
  );
  LUT5 #(
    .INIT(32'hac000000)
  ) __6074__ (
    .I4(__2390__),
    .I3(__2389__),
    .I2(__2379__),
    .I1(__2388__),
    .I0(__2387__),
    .O(__2391__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __6075__ (
    .I5(__858__),
    .I4(__964__),
    .I3(__944__),
    .I2(__960__),
    .I1(__954__),
    .I0(__962__),
    .O(__2392__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6076__ (
    .I1(__954__),
    .I0(__813__),
    .O(__2393__)
  );
  LUT6 #(
    .INIT(64'h0000000000bfbfbf)
  ) __6077__ (
    .I5(__2393__),
    .I4(__944__),
    .I3(__561__),
    .I2(__1347__),
    .I1(__965__),
    .I0(__2392__),
    .O(__2394__)
  );
  LUT6 #(
    .INIT(64'h4f440000ffcc0000)
  ) __6078__ (
    .I5(__858__),
    .I4(__1624__),
    .I3(__2394__),
    .I2(__814__),
    .I1(__1665__),
    .I0(__812__),
    .O(__2395__)
  );
  LUT6 #(
    .INIT(64'h5455555555555555)
  ) __6079__ (
    .I5(__1623__),
    .I4(__1506__),
    .I3(__1505__),
    .I2(__1508__),
    .I1(__1507__),
    .I0(__1646__),
    .O(__2396__)
  );
  LUT6 #(
    .INIT(64'hffffffffbf000000)
  ) __6080__ (
    .I5(__2396__),
    .I4(__2395__),
    .I3(__2391__),
    .I2(__2386__),
    .I1(__2385__),
    .I0(__2380__),
    .O(__2397__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6081__ (
    .I2(__954__),
    .I1(__2397__),
    .I0(__808__),
    .O(__2398__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6082__ (
    .I2(__944__),
    .I1(__1647__),
    .I0(__745__),
    .O(__2399__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __6083__ (
    .I2(__662__),
    .I1(__2250__),
    .I0(__1124__),
    .O(__2400__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __6084__ (
    .I2(__663__),
    .I1(__2249__),
    .I0(__424__),
    .O(__2401__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6085__ (
    .I2(__1511__),
    .I1(__89__),
    .I0(__232__),
    .O(__2402__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __6086__ (
    .I5(__944__),
    .I4(__936__),
    .I3(__927__),
    .I2(__924__),
    .I1(__899__),
    .I0(__917__),
    .O(__2403__)
  );
  LUT4 #(
    .INIT(16'he7ee)
  ) __6087__ (
    .I3(__1643__),
    .I2(__1637__),
    .I1(__1638__),
    .I0(__1640__),
    .O(__2404__)
  );
  LUT6 #(
    .INIT(64'h108000c000000000)
  ) __6088__ (
    .I5(__603__),
    .I4(__1643__),
    .I3(__1640__),
    .I2(__1639__),
    .I1(__1638__),
    .I0(__1637__),
    .O(__2405__)
  );
  LUT5 #(
    .INIT(32'h00f4f0f0)
  ) __6089__ (
    .I4(__662__),
    .I3(__2405__),
    .I2(__1172__),
    .I1(__603__),
    .I0(__2404__),
    .O(__2406__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __6090__ (
    .I2(__663__),
    .I1(__1598__),
    .I0(__1635__),
    .O(__2407__)
  );
  LUT6 #(
    .INIT(64'h55555d5500000800)
  ) __6091__ (
    .I5(__1233__),
    .I4(__1458__),
    .I3(__1460__),
    .I2(__1459__),
    .I1(__1457__),
    .I0(__2407__),
    .O(__2408__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6092__ (
    .I2(__944__),
    .I1(__988__),
    .I0(__1367__),
    .O(__2409__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __6093__ (
    .I5(__589__),
    .I4(__1119__),
    .I3(__663__),
    .I2(__648__),
    .I1(__662__),
    .I0(__647__),
    .O(__2410__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __6094__ (
    .I5(__589__),
    .I4(__531__),
    .I3(__663__),
    .I2(__1109__),
    .I1(__662__),
    .I0(__532__),
    .O(__2411__)
  );
  LUT6 #(
    .INIT(64'h01f700f300ff00ff)
  ) __6095__ (
    .I5(__603__),
    .I4(__1617__),
    .I3(__2411__),
    .I2(__2410__),
    .I1(__1613__),
    .I0(__1614__),
    .O(__2412__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6096__ (
    .I2(__589__),
    .I1(__2412__),
    .I0(__531__),
    .O(__2413__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __6097__ (
    .I5(__954__),
    .I4(__242__),
    .I3(__370__),
    .I2(__229__),
    .I1(__202__),
    .I0(__227__),
    .O(__2414__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __6098__ (
    .I3(__663__),
    .I2(__603__),
    .I1(__1459__),
    .I0(__1304__),
    .O(__2415__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __6099__ (
    .I3(__663__),
    .I2(__2282__),
    .I1(__1419__),
    .I0(__1285__),
    .O(__2416__)
  );
  LUT6 #(
    .INIT(64'haaaaa2a6aaaaa6a6)
  ) __6100__ (
    .I5(__603__),
    .I4(__1884__),
    .I3(__1899__),
    .I2(__1893__),
    .I1(__1617__),
    .I0(__2249__),
    .O(__2417__)
  );
  LUT6 #(
    .INIT(64'hbfffffffa0000000)
  ) __6101__ (
    .I5(__1122__),
    .I4(__662__),
    .I3(__603__),
    .I2(__2417__),
    .I1(__2247__),
    .I0(__2248__),
    .O(__2418__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __6102__ (
    .I5(__944__),
    .I4(__304__),
    .I3(__858__),
    .I2(__152__),
    .I1(__954__),
    .I0(__310__),
    .O(__2419__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6103__ (
    .I1(__1790__),
    .I0(__2419__),
    .O(__2420__)
  );
  LUT6 #(
    .INIT(64'h00000ee00ee00000)
  ) __6104__ (
    .I5(__1795__),
    .I4(__367__),
    .I3(__1785__),
    .I2(__222__),
    .I1(__224__),
    .I0(__1786__),
    .O(__2421__)
  );
  LUT5 #(
    .INIT(32'h0ee00000)
  ) __6105__ (
    .I4(__2421__),
    .I3(__1787__),
    .I2(__225__),
    .I1(__1797__),
    .I0(__219__),
    .O(__2422__)
  );
  LUT6 #(
    .INIT(64'h0000077007700000)
  ) __6106__ (
    .I5(__227__),
    .I4(__1792__),
    .I3(__1793__),
    .I2(__366__),
    .I1(__1797__),
    .I0(__219__),
    .O(__2423__)
  );
  LUT6 #(
    .INIT(64'h0000077007700000)
  ) __6107__ (
    .I5(__1796__),
    .I4(__220__),
    .I3(__1789__),
    .I2(__365__),
    .I1(__224__),
    .I0(__1786__),
    .O(__2424__)
  );
  LUT6 #(
    .INIT(64'h82aaaaaaaaaaaaaa)
  ) __6108__ (
    .I5(__2424__),
    .I4(__2423__),
    .I3(__2422__),
    .I2(__216__),
    .I1(__1788__),
    .I0(__2420__),
    .O(__2425__)
  );
  LUT6 #(
    .INIT(64'haaaacaaaaaaaaaaa)
  ) __6109__ (
    .I5(__858__),
    .I4(__229__),
    .I3(__242__),
    .I2(__370__),
    .I1(__2425__),
    .I0(__146__),
    .O(__2426__)
  );
  LUT5 #(
    .INIT(32'h80ef0000)
  ) __6110__ (
    .I4(__662__),
    .I3(__1598__),
    .I2(__1682__),
    .I1(__1681__),
    .I0(__1680__),
    .O(__2427__)
  );
  LUT6 #(
    .INIT(64'hcc77f0f077ccf0f0)
  ) __6111__ (
    .I5(g3229),
    .I4(__2427__),
    .I3(__2287__),
    .I2(__601__),
    .I1(__2285__),
    .I0(__2369__),
    .O(__2428__)
  );
  LUT5 #(
    .INIT(32'h44ff00f0)
  ) __6112__ (
    .I4(__1806__),
    .I3(__1647__),
    .I2(__1674__),
    .I1(__1036__),
    .I0(__1805__),
    .O(__2429__)
  );
  LUT4 #(
    .INIT(16'haccc)
  ) __6113__ (
    .I3(__663__),
    .I2(__603__),
    .I1(__774__),
    .I0(__1893__),
    .O(__2430__)
  );
  LUT6 #(
    .INIT(64'h1320132013001320)
  ) __6114__ (
    .I5(__1484__),
    .I4(__1483__),
    .I3(__1485__),
    .I2(__1486__),
    .I1(__1497__),
    .I0(__1611__),
    .O(__2431__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __6115__ (
    .I2(__589__),
    .I1(__1640__),
    .I0(__1008__),
    .O(__2432__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __6116__ (
    .I3(__662__),
    .I2(__603__),
    .I1(__1436__),
    .I0(__847__),
    .O(__2433__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __6117__ (
    .I5(__858__),
    .I4(__242__),
    .I3(__370__),
    .I2(__229__),
    .I1(__204__),
    .I0(__227__),
    .O(__2434__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6118__ (
    .I2(__1479__),
    .I1(__1418__),
    .I0(__1477__),
    .O(__2435__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6119__ (
    .I2(__1479__),
    .I1(__1474__),
    .I0(__1456__),
    .O(__2436__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __6120__ (
    .I2(__663__),
    .I1(__1606__),
    .I0(__203__),
    .O(__2437__)
  );
  LUT4 #(
    .INIT(16'hf8ff)
  ) __6121__ (
    .I3(__603__),
    .I2(__1570__),
    .I1(__1585__),
    .I0(__1580__),
    .O(__2438__)
  );
  LUT5 #(
    .INIT(32'h80000000)
  ) __6122__ (
    .I4(__1574__),
    .I3(__1569__),
    .I2(__1564__),
    .I1(__1561__),
    .I0(__2438__),
    .O(__2439__)
  );
  LUT6 #(
    .INIT(64'h4000000000000000)
  ) __6123__ (
    .I5(__1574__),
    .I4(__1569__),
    .I3(__1564__),
    .I2(__1561__),
    .I1(__1544__),
    .I0(__1542__),
    .O(__2440__)
  );
  LUT4 #(
    .INIT(16'h1428)
  ) __6124__ (
    .I3(__1422__),
    .I2(__1417__),
    .I1(__1546__),
    .I0(__1539__),
    .O(__2441__)
  );
  LUT4 #(
    .INIT(16'h0990)
  ) __6125__ (
    .I3(__1432__),
    .I2(__1550__),
    .I1(__1572__),
    .I0(__1540__),
    .O(__2442__)
  );
  LUT4 #(
    .INIT(16'h1428)
  ) __6126__ (
    .I3(__1419__),
    .I2(__1424__),
    .I1(__1537__),
    .I0(__1538__),
    .O(__2443__)
  );
  LUT4 #(
    .INIT(16'h0990)
  ) __6127__ (
    .I3(__1430__),
    .I2(__1548__),
    .I1(__1565__),
    .I0(__1536__),
    .O(__2444__)
  );
  LUT6 #(
    .INIT(64'h8000000000000000)
  ) __6128__ (
    .I5(__1581__),
    .I4(__1577__),
    .I3(__2444__),
    .I2(__2443__),
    .I1(__2442__),
    .I0(__2441__),
    .O(__2445__)
  );
  LUT3 #(
    .INIT(8'h10)
  ) __6129__ (
    .I2(__1544__),
    .I1(__1543__),
    .I0(__1542__),
    .O(__2446__)
  );
  LUT5 #(
    .INIT(32'hcd000000)
  ) __6130__ (
    .I4(__589__),
    .I3(__603__),
    .I2(__1570__),
    .I1(__2446__),
    .I0(__2445__),
    .O(__2447__)
  );
  LUT6 #(
    .INIT(64'hffff0707ff00ff00)
  ) __6131__ (
    .I5(__2447__),
    .I4(__1543__),
    .I3(__1155__),
    .I2(__2440__),
    .I1(__1542__),
    .I0(__2439__),
    .O(__2448__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __6132__ (
    .I3(__663__),
    .I2(__2282__),
    .I1(__2140__),
    .I0(__756__),
    .O(__2449__)
  );
  LUT5 #(
    .INIT(32'ha000cccc)
  ) __6133__ (
    .I4(__589__),
    .I3(__1682__),
    .I2(__1681__),
    .I1(__389__),
    .I0(__1680__),
    .O(__2450__)
  );
  LUT5 #(
    .INIT(32'ha000cccc)
  ) __6134__ (
    .I4(__663__),
    .I3(__1597__),
    .I2(__1596__),
    .I1(__782__),
    .I0(__1595__),
    .O(__2451__)
  );
  LUT4 #(
    .INIT(16'haccc)
  ) __6135__ (
    .I3(__589__),
    .I2(__603__),
    .I1(__815__),
    .I0(__1751__),
    .O(__2452__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6136__ (
    .I2(__662__),
    .I1(__1644__),
    .I0(__1181__),
    .O(__2453__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __6137__ (
    .I5(__764__),
    .I4(__573__),
    .I3(__858__),
    .I2(__745__),
    .I1(__688__),
    .I0(__741__),
    .O(__2454__)
  );
  LUT4 #(
    .INIT(16'h0008)
  ) __6138__ (
    .I3(__1448__),
    .I2(__1446__),
    .I1(__1444__),
    .I0(__1450__),
    .O(__2455__)
  );
  LUT5 #(
    .INIT(32'hb8f0f0f0)
  ) __6139__ (
    .I4(__663__),
    .I3(__1598__),
    .I2(__790__),
    .I1(__1635__),
    .I0(__2455__),
    .O(__2456__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __6140__ (
    .I3(__663__),
    .I2(__603__),
    .I1(__1442__),
    .I0(__839__),
    .O(__2457__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __6141__ (
    .I5(__944__),
    .I4(__93__),
    .I3(__73__),
    .I2(__748__),
    .I1(__1042__),
    .I0(__1047__),
    .O(__2458__)
  );
  LUT5 #(
    .INIT(32'h21a522aa)
  ) __6142__ (
    .I4(__944__),
    .I3(__954__),
    .I2(__229__),
    .I1(__231__),
    .I0(__367__),
    .O(__2459__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __6143__ (
    .I3(__663__),
    .I2(__603__),
    .I1(__1456__),
    .I0(__1324__),
    .O(__2460__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6144__ (
    .I2(__954__),
    .I1(__986__),
    .I0(__1396__),
    .O(__2461__)
  );
  LUT6 #(
    .INIT(64'haaaaa2a6aaaaa6a6)
  ) __6145__ (
    .I5(__603__),
    .I4(__1712__),
    .I3(__1710__),
    .I2(__1705__),
    .I1(__2089__),
    .I0(__2211__),
    .O(__2462__)
  );
  LUT6 #(
    .INIT(64'hfa000f0fcccccccc)
  ) __6146__ (
    .I5(__662__),
    .I4(__603__),
    .I3(__2462__),
    .I2(__2209__),
    .I1(__555__),
    .I0(__2210__),
    .O(__2463__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __6147__ (
    .I3(__589__),
    .I2(__603__),
    .I1(__1426__),
    .I0(__1313__),
    .O(__2464__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __6148__ (
    .I3(__589__),
    .I2(__603__),
    .I1(__1440__),
    .I0(__840__),
    .O(__2465__)
  );
  LUT5 #(
    .INIT(32'h21a522aa)
  ) __6149__ (
    .I4(__944__),
    .I3(__954__),
    .I2(__745__),
    .I1(__752__),
    .I0(__760__),
    .O(__2466__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __6150__ (
    .I2(__589__),
    .I1(__2212__),
    .I0(__553__),
    .O(__2467__)
  );
  LUT6 #(
    .INIT(64'h0f005555cccccccc)
  ) __6151__ (
    .I5(__662__),
    .I4(__603__),
    .I3(__1617__),
    .I2(__1614__),
    .I1(__1106__),
    .I0(__1613__),
    .O(__2468__)
  );
  LUT4 #(
    .INIT(16'h8000)
  ) __6152__ (
    .I3(__1499__),
    .I2(__1500__),
    .I1(__1498__),
    .I0(__215__),
    .O(__2469__)
  );
  LUT5 #(
    .INIT(32'h0000125a)
  ) __6153__ (
    .I4(g3234),
    .I3(__1623__),
    .I2(__1501__),
    .I1(__215__),
    .I0(__2469__),
    .O(__2470__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __6154__ (
    .I2(__663__),
    .I1(__2327__),
    .I0(__71__),
    .O(__2471__)
  );
  LUT5 #(
    .INIT(32'h0c66cccc)
  ) __6155__ (
    .I4(__589__),
    .I3(__1598__),
    .I2(__603__),
    .I1(__1236__),
    .I0(__1237__),
    .O(__2472__)
  );
  LUT5 #(
    .INIT(32'ha000cccc)
  ) __6156__ (
    .I4(__954__),
    .I3(__1951__),
    .I2(__2094__),
    .I1(__104__),
    .I0(__266__),
    .O(__2473__)
  );
  LUT5 #(
    .INIT(32'h6c9ccccc)
  ) __6157__ (
    .I4(__1597__),
    .I3(__1596__),
    .I2(__1595__),
    .I1(__1897__),
    .I0(__1877__),
    .O(__2474__)
  );
  LUT6 #(
    .INIT(64'hf0f03355f0f0f0f0)
  ) __6158__ (
    .I5(__2015__),
    .I4(__2012__),
    .I3(__2008__),
    .I2(__1454__),
    .I1(__2002__),
    .I0(__2474__),
    .O(__2475__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6159__ (
    .I2(__589__),
    .I1(__2475__),
    .I0(__534__),
    .O(__2476__)
  );
  LUT5 #(
    .INIT(32'hcd000000)
  ) __6160__ (
    .I4(__662__),
    .I3(__603__),
    .I2(__1899__),
    .I1(__1922__),
    .I0(__1921__),
    .O(__2477__)
  );
  LUT6 #(
    .INIT(64'hffff0707ff00ff00)
  ) __6161__ (
    .I5(__2477__),
    .I4(__1597__),
    .I3(__1078__),
    .I2(__1916__),
    .I1(__1595__),
    .I0(__1915__),
    .O(__2478__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __6162__ (
    .I5(__944__),
    .I4(__93__),
    .I3(__73__),
    .I2(__748__),
    .I1(__1046__),
    .I0(__797__),
    .O(__2479__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __6163__ (
    .I2(__662__),
    .I1(__2249__),
    .I0(__436__),
    .O(__2480__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __6164__ (
    .I5(__944__),
    .I4(__242__),
    .I3(__370__),
    .I2(__229__),
    .I1(__206__),
    .I0(__366__),
    .O(__2481__)
  );
  LUT6 #(
    .INIT(64'h8000010000000000)
  ) __6165__ (
    .I5(__1761__),
    .I4(__1760__),
    .I3(__1759__),
    .I2(__1755__),
    .I1(__1744__),
    .I0(__1735__),
    .O(__2482__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __6166__ (
    .I1(__1753__),
    .I0(__2482__),
    .O(__2483__)
  );
  LUT6 #(
    .INIT(64'hf0f03355f0f0f0f0)
  ) __6167__ (
    .I5(__1864__),
    .I4(__1861__),
    .I3(__1857__),
    .I2(__1442__),
    .I1(__1851__),
    .I0(__2483__),
    .O(__2484__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6168__ (
    .I2(__662__),
    .I1(__2484__),
    .I0(__718__),
    .O(__2485__)
  );
  LUT5 #(
    .INIT(32'h44ff00f0)
  ) __6169__ (
    .I4(__2094__),
    .I3(__1647__),
    .I2(__2056__),
    .I1(__266__),
    .I0(__1951__),
    .O(__2486__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6170__ (
    .I2(__663__),
    .I1(__2412__),
    .I0(__1109__),
    .O(__2487__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __6171__ (
    .I3(__663__),
    .I2(__603__),
    .I1(__1430__),
    .I0(__1300__),
    .O(__2488__)
  );
  LUT6 #(
    .INIT(64'h4f0f4f0000000000)
  ) __6172__ (
    .I5(__858__),
    .I4(__1674__),
    .I3(__1806__),
    .I2(__1647__),
    .I1(__1036__),
    .I0(__1805__),
    .O(__2489__)
  );
  LUT6 #(
    .INIT(64'h3fffff3faaaaaaaa)
  ) __6173__ (
    .I5(__2489__),
    .I4(g3229),
    .I3(__1810__),
    .I2(__1809__),
    .I1(__1808__),
    .I0(__976__),
    .O(__2490__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __6174__ (
    .I5(__764__),
    .I4(__573__),
    .I3(__858__),
    .I2(__745__),
    .I1(__651__),
    .I0(__768__),
    .O(__2491__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __6175__ (
    .I5(__944__),
    .I4(__936__),
    .I3(__927__),
    .I2(__924__),
    .I1(__887__),
    .I0(__913__),
    .O(__2492__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __6176__ (
    .I2(__663__),
    .I1(__2250__),
    .I0(__1125__),
    .O(__2493__)
  );
  LUT5 #(
    .INIT(32'ha000cccc)
  ) __6177__ (
    .I4(__858__),
    .I3(__1981__),
    .I2(__354__),
    .I1(__270__),
    .I0(__1800__),
    .O(__2494__)
  );
  LUT4 #(
    .INIT(16'haccc)
  ) __6178__ (
    .I3(__858__),
    .I2(__752__),
    .I1(__678__),
    .I0(__1646__),
    .O(__2495__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __6179__ (
    .I3(__662__),
    .I2(__603__),
    .I1(__1460__),
    .I0(__795__),
    .O(__2496__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __6180__ (
    .I2(__663__),
    .I1(__2211__),
    .I0(__150__),
    .O(__2497__)
  );
  LUT4 #(
    .INIT(16'h8000)
  ) __6181__ (
    .I3(__1491__),
    .I2(__1493__),
    .I1(__1492__),
    .I0(__1494__),
    .O(__2498__)
  );
  LUT4 #(
    .INIT(16'h0006)
  ) __6182__ (
    .I3(__1497__),
    .I2(__1611__),
    .I1(__1490__),
    .I0(__2498__),
    .O(__2499__)
  );
  LUT6 #(
    .INIT(64'hf0f0ff00aaaaaaaa)
  ) __6183__ (
    .I5(__858__),
    .I4(__142__),
    .I3(__1781__),
    .I2(__158__),
    .I1(__144__),
    .I0(__1378__),
    .O(__2500__)
  );
  LUT3 #(
    .INIT(8'h70)
  ) __6184__ (
    .I2(__2117__),
    .I1(__858__),
    .I0(__282__),
    .O(__2501__)
  );
  LUT6 #(
    .INIT(64'h5455555555555555)
  ) __6185__ (
    .I5(__1623__),
    .I4(__1506__),
    .I3(__1505__),
    .I2(__1508__),
    .I1(__1507__),
    .I0(__1982__),
    .O(__2502__)
  );
  LUT6 #(
    .INIT(64'h0f080f0f0f0f0f0f)
  ) __6186__ (
    .I5(__2118__),
    .I4(__2109__),
    .I3(__2104__),
    .I2(__2502__),
    .I1(__2501__),
    .I0(__2115__),
    .O(__2503__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __6187__ (
    .I2(__858__),
    .I1(__2503__),
    .I0(__272__),
    .O(__2504__)
  );
  LUT6 #(
    .INIT(64'hd8fad850d850d8fa)
  ) __6188__ (
    .I5(g3229),
    .I4(__1930__),
    .I3(__1928__),
    .I2(__135__),
    .I1(__1932__),
    .I0(__2173__),
    .O(__2505__)
  );
  LUT5 #(
    .INIT(32'h0030aaaa)
  ) __6189__ (
    .I4(__589__),
    .I3(__1544__),
    .I2(__1543__),
    .I1(__1542__),
    .I0(__1005__),
    .O(__2506__)
  );
  LUT3 #(
    .INIT(8'h10)
  ) __6190__ (
    .I2(__1643__),
    .I1(__1572__),
    .I0(__1565__),
    .O(__2507__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __6191__ (
    .I5(__589__),
    .I4(__1193__),
    .I3(__663__),
    .I2(__1195__),
    .I1(__662__),
    .I0(__1194__),
    .O(__2508__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __6192__ (
    .I5(__589__),
    .I4(__1187__),
    .I3(__663__),
    .I2(__1189__),
    .I1(__662__),
    .I0(__1188__),
    .O(__2509__)
  );
  LUT6 #(
    .INIT(64'h000300007773ffff)
  ) __6193__ (
    .I5(__1672__),
    .I4(__603__),
    .I3(__2509__),
    .I2(__2508__),
    .I1(__2507__),
    .I0(__1570__),
    .O(__2510__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __6194__ (
    .I2(__662__),
    .I1(__2510__),
    .I0(__1191__),
    .O(__2511__)
  );
  LUT6 #(
    .INIT(64'haaaaa2a6aaaaa6a6)
  ) __6195__ (
    .I5(__603__),
    .I4(__1751__),
    .I3(__1757__),
    .I2(__1742__),
    .I1(__2140__),
    .I0(__2279__),
    .O(__2512__)
  );
  LUT6 #(
    .INIT(64'hfa000f0fcccccccc)
  ) __6196__ (
    .I5(__662__),
    .I4(__603__),
    .I3(__2512__),
    .I2(__2277__),
    .I1(__621__),
    .I0(__2278__),
    .O(__2513__)
  );
  LUT5 #(
    .INIT(32'he0000000)
  ) __6197__ (
    .I4(__1597__),
    .I3(__1595__),
    .I2(__2015__),
    .I1(__2007__),
    .I0(__2005__),
    .O(__2514__)
  );
  LUT6 #(
    .INIT(64'hdffffff720000008)
  ) __6198__ (
    .I5(__1888__),
    .I4(__1895__),
    .I3(__1886__),
    .I2(__1879__),
    .I1(__2002__),
    .I0(__2361__),
    .O(__2515__)
  );
  LUT6 #(
    .INIT(64'h01000f000f000f00)
  ) __6199__ (
    .I5(__1597__),
    .I4(__1595__),
    .I3(__2015__),
    .I2(__2012__),
    .I1(__2007__),
    .I0(__2005__),
    .O(__2516__)
  );
  LUT6 #(
    .INIT(64'h0f0f4444ff00ff00)
  ) __6200__ (
    .I5(__589__),
    .I4(__2516__),
    .I3(__1207__),
    .I2(__2515__),
    .I1(__1458__),
    .I0(__2514__),
    .O(__2517__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6201__ (
    .I1(__568__),
    .I0(__2149__),
    .O(__2518__)
  );
  LUT6 #(
    .INIT(64'h00007fff00008000)
  ) __6202__ (
    .I5(__512__),
    .I4(__2151__),
    .I3(__567__),
    .I2(__605__),
    .I1(__604__),
    .I0(__2518__),
    .O(__2519__)
  );
  LUT4 #(
    .INIT(16'h0080)
  ) __6203__ (
    .I3(__745__),
    .I2(__944__),
    .I1(__764__),
    .I0(__573__),
    .O(__2520__)
  );
  LUT5 #(
    .INIT(32'h3f00aaaa)
  ) __6204__ (
    .I4(__2520__),
    .I3(__1838__),
    .I2(__1835__),
    .I1(__1822__),
    .I0(__670__),
    .O(__2521__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6205__ (
    .I2(__944__),
    .I1(__142__),
    .I0(__1363__),
    .O(__2522__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __6206__ (
    .I3(__662__),
    .I2(__603__),
    .I1(__1424__),
    .I0(__1317__),
    .O(__2523__)
  );
  LUT5 #(
    .INIT(32'he0000000)
  ) __6207__ (
    .I4(__1761__),
    .I3(__1759__),
    .I2(__1864__),
    .I1(__1856__),
    .I0(__1854__),
    .O(__2524__)
  );
  LUT5 #(
    .INIT(32'hdff72008)
  ) __6208__ (
    .I4(__1746__),
    .I3(__1753__),
    .I2(__1737__),
    .I1(__1851__),
    .I0(__2482__),
    .O(__2525__)
  );
  LUT6 #(
    .INIT(64'h01000f000f000f00)
  ) __6209__ (
    .I5(__1761__),
    .I4(__1759__),
    .I3(__1864__),
    .I2(__1861__),
    .I1(__1856__),
    .I0(__1854__),
    .O(__2526__)
  );
  LUT6 #(
    .INIT(64'h0f0f4444ff00ff00)
  ) __6210__ (
    .I5(__662__),
    .I4(__2526__),
    .I3(__712__),
    .I2(__2525__),
    .I1(__1446__),
    .I0(__2524__),
    .O(__2527__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __6211__ (
    .I2(__589__),
    .I1(__1593__),
    .I0(__1254__),
    .O(__2528__)
  );
  LUT5 #(
    .INIT(32'h0030aaaa)
  ) __6212__ (
    .I4(__662__),
    .I3(__1543__),
    .I2(__1544__),
    .I1(__1542__),
    .I0(__1003__),
    .O(__2529__)
  );
  LUT4 #(
    .INIT(16'h0baa)
  ) __6213__ (
    .I3(__858__),
    .I2(__1624__),
    .I1(__2048__),
    .I0(__973__),
    .O(__2530__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __6214__ (
    .I5(__944__),
    .I4(__764__),
    .I3(__573__),
    .I2(__745__),
    .I1(__689__),
    .I0(__772__),
    .O(__2531__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __6215__ (
    .I2(__944__),
    .I1(__2503__),
    .I0(__271__),
    .O(__2532__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __6216__ (
    .I5(__858__),
    .I4(__936__),
    .I3(__927__),
    .I2(__924__),
    .I1(__895__),
    .I0(__915__),
    .O(__2533__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __6217__ (
    .I3(__663__),
    .I2(__2282__),
    .I1(__1417__),
    .I0(__1282__),
    .O(__2534__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __6218__ (
    .I5(__944__),
    .I4(__936__),
    .I3(__927__),
    .I2(__924__),
    .I1(__884__),
    .I0(__912__),
    .O(__2535__)
  );
  LUT5 #(
    .INIT(32'h6c9ccccc)
  ) __6219__ (
    .I4(__1682__),
    .I3(__1681__),
    .I2(__1680__),
    .I1(__1679__),
    .I0(__1677__),
    .O(__2536__)
  );
  LUT6 #(
    .INIT(64'hf0f03355f0f0f0f0)
  ) __6220__ (
    .I5(__1732__),
    .I4(__1728__),
    .I3(__1697__),
    .I2(__1408__),
    .I1(__1684__),
    .I0(__2536__),
    .O(__2537__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6221__ (
    .I2(__662__),
    .I1(__2537__),
    .I0(__520__),
    .O(__2538__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6222__ (
    .I2(__663__),
    .I1(__1968__),
    .I0(__1244__),
    .O(__2539__)
  );
  LUT3 #(
    .INIT(8'he2)
  ) __6223__ (
    .I2(__988__),
    .I1(__954__),
    .I0(__1368__),
    .O(__2540__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __6224__ (
    .I5(__764__),
    .I4(__573__),
    .I3(__858__),
    .I2(__745__),
    .I1(__684__),
    .I0(__770__),
    .O(__2541__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6225__ (
    .I2(__589__),
    .I1(__1644__),
    .I0(__1179__),
    .O(__2542__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6226__ (
    .I2(__1479__),
    .I1(__1437__),
    .I0(__1468__),
    .O(__2543__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6227__ (
    .I2(__589__),
    .I1(__1962__),
    .I0(__439__),
    .O(__2544__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __6228__ (
    .I5(__944__),
    .I4(__764__),
    .I3(__573__),
    .I2(__745__),
    .I1(__692__),
    .I0(__765__),
    .O(__2545__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __6229__ (
    .I5(__858__),
    .I4(__936__),
    .I3(__927__),
    .I2(__924__),
    .I1(__886__),
    .I0(__912__),
    .O(__2546__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __6230__ (
    .I2(__589__),
    .I1(__1957__),
    .I0(__361__),
    .O(__2547__)
  );
  LUT4 #(
    .INIT(16'h125a)
  ) __6231__ (
    .I3(__954__),
    .I2(__796__),
    .I1(__875__),
    .I0(__1667__),
    .O(__2548__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __6232__ (
    .I2(__662__),
    .I1(__2411__),
    .I0(__447__),
    .O(__2549__)
  );
  LUT6 #(
    .INIT(64'h0100000100000000)
  ) __6233__ (
    .I5(__868__),
    .I4(__1817__),
    .I3(__1646__),
    .I2(__1966__),
    .I1(g1943),
    .I0(__867__),
    .O(__2550__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __6234__ (
    .I5(__944__),
    .I4(__670__),
    .I3(__858__),
    .I2(__672__),
    .I1(__954__),
    .I0(__671__),
    .O(__2551__)
  );
  LUT3 #(
    .INIT(8'h08)
  ) __6235__ (
    .I2(__1818__),
    .I1(__2343__),
    .I0(__2342__),
    .O(__2552__)
  );
  LUT6 #(
    .INIT(64'h0000df0f00000000)
  ) __6236__ (
    .I5(__969__),
    .I4(__968__),
    .I3(__868__),
    .I2(__2346__),
    .I1(__2552__),
    .I0(__2551__),
    .O(__2553__)
  );
  LUT6 #(
    .INIT(64'hffffffff000f00bb)
  ) __6237__ (
    .I5(__2553__),
    .I4(__2348__),
    .I3(__2347__),
    .I2(__2550__),
    .I1(__2346__),
    .I0(__762__),
    .O(__2554__)
  );
  LUT2 #(
    .INIT(4'h7)
  ) __6238__ (
    .I1(__1682__),
    .I0(__1680__),
    .O(__2555__)
  );
  LUT6 #(
    .INIT(64'h5555fccf55555555)
  ) __6239__ (
    .I5(__1732__),
    .I4(__1728__),
    .I3(__1677__),
    .I2(__2555__),
    .I1(__1697__),
    .I0(__1407__),
    .O(__2556__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __6240__ (
    .I2(__589__),
    .I1(__2556__),
    .I0(__617__),
    .O(__2557__)
  );
  LUT4 #(
    .INIT(16'hf0ee)
  ) __6241__ (
    .I3(__939__),
    .I2(__938__),
    .I1(__954__),
    .I0(__937__),
    .O(__2558__)
  );
  LUT5 #(
    .INIT(32'hf0f0ccaa)
  ) __6242__ (
    .I4(__98__),
    .I3(__954__),
    .I2(__97__),
    .I1(__2558__),
    .I0(__94__),
    .O(__2559__)
  );
  LUT5 #(
    .INIT(32'hf0f0ccaa)
  ) __6243__ (
    .I4(__848__),
    .I3(__954__),
    .I2(__744__),
    .I1(__2559__),
    .I0(__771__),
    .O(__2560__)
  );
  LUT5 #(
    .INIT(32'ha000cccc)
  ) __6244__ (
    .I4(__954__),
    .I3(__968__),
    .I2(__1646__),
    .I1(__803__),
    .I0(__1648__),
    .O(__2561__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __6245__ (
    .I3(__663__),
    .I2(__603__),
    .I1(__1446__),
    .I0(__833__),
    .O(__2562__)
  );
  LUT6 #(
    .INIT(64'hd8fad850d850d8fa)
  ) __6246__ (
    .I5(g3229),
    .I4(__2287__),
    .I3(__2286__),
    .I2(__560__),
    .I1(__2285__),
    .I0(__2427__),
    .O(__2563__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6247__ (
    .I2(__944__),
    .I1(__356__),
    .I0(__354__),
    .O(__2564__)
  );
  LUT6 #(
    .INIT(64'haa3aaaaaaaaaaaaa)
  ) __6248__ (
    .I5(__858__),
    .I4(__93__),
    .I3(__748__),
    .I2(__73__),
    .I1(__1055__),
    .I0(__732__),
    .O(__2565__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __6249__ (
    .I5(__944__),
    .I4(__474__),
    .I3(__858__),
    .I2(__361__),
    .I1(__954__),
    .I0(__477__),
    .O(__2566__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6250__ (
    .I2(__944__),
    .I1(__269__),
    .I0(__266__),
    .O(__2567__)
  );
  LUT5 #(
    .INIT(32'h80ef0000)
  ) __6251__ (
    .I4(__662__),
    .I3(__1598__),
    .I2(__1543__),
    .I1(__1544__),
    .I0(__1542__),
    .O(__2568__)
  );
  LUT6 #(
    .INIT(64'hd8fad850d850d8fa)
  ) __6252__ (
    .I5(g3229),
    .I4(__2065__),
    .I3(__2064__),
    .I2(__1211__),
    .I1(__2063__),
    .I0(__2568__),
    .O(__2569__)
  );
  LUT5 #(
    .INIT(32'hdff72008)
  ) __6253__ (
    .I4(__1883__),
    .I3(__1890__),
    .I2(__1881__),
    .I1(__2002__),
    .I0(__2362__),
    .O(__2570__)
  );
  LUT6 #(
    .INIT(64'h0f0f33550f0f0f0f)
  ) __6254__ (
    .I5(__2015__),
    .I4(__2012__),
    .I3(__2008__),
    .I2(__1884__),
    .I1(__2002__),
    .I0(__2570__),
    .O(__2571__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6255__ (
    .I2(__662__),
    .I1(__2571__),
    .I0(__649__),
    .O(__2572__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6256__ (
    .I2(__944__),
    .I1(__868__),
    .I0(__1360__),
    .O(__2573__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6257__ (
    .I2(__663__),
    .I1(__2537__),
    .I0(__616__),
    .O(__2574__)
  );
  LUT4 #(
    .INIT(16'haccc)
  ) __6258__ (
    .I3(__944__),
    .I2(__752__),
    .I1(__673__),
    .I0(__1649__),
    .O(__2575__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __6259__ (
    .I3(__662__),
    .I2(__2282__),
    .I1(__1454__),
    .I0(__1260__),
    .O(__2576__)
  );
  LUT6 #(
    .INIT(64'h4545ff000505ff00)
  ) __6260__ (
    .I5(__858__),
    .I4(__944__),
    .I3(__971__),
    .I2(__2048__),
    .I1(__973__),
    .I0(__1624__),
    .O(__2577__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6261__ (
    .I2(__944__),
    .I1(__1953__),
    .I0(__110__),
    .O(__2578__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __6262__ (
    .I3(__663__),
    .I2(__603__),
    .I1(__1408__),
    .I0(__430__),
    .O(__2579__)
  );
  LUT5 #(
    .INIT(32'hf0f0ccaa)
  ) __6263__ (
    .I4(__267__),
    .I3(__954__),
    .I2(__264__),
    .I1(__2560__),
    .I0(__244__),
    .O(__2580__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __6264__ (
    .I5(__589__),
    .I4(__625__),
    .I3(__663__),
    .I2(__628__),
    .I1(__662__),
    .I0(__627__),
    .O(__2581__)
  );
  LUT5 #(
    .INIT(32'h80ef0000)
  ) __6265__ (
    .I4(__663__),
    .I3(__1598__),
    .I2(__1761__),
    .I1(__1760__),
    .I0(__1759__),
    .O(__2582__)
  );
  LUT6 #(
    .INIT(64'hcc77f0f077ccf0f0)
  ) __6266__ (
    .I5(g3229),
    .I4(__2582__),
    .I3(__2070__),
    .I2(__631__),
    .I1(__2069__),
    .I0(__2581__),
    .O(__2583__)
  );
  LUT3 #(
    .INIT(8'h4f)
  ) __6267__ (
    .I2(__1511__),
    .I1(__1509__),
    .I0(__1510__),
    .O(__2584__)
  );
  LUT6 #(
    .INIT(64'haaaaa2a6aaaaa6a6)
  ) __6268__ (
    .I5(__603__),
    .I4(__1572__),
    .I3(__1570__),
    .I2(__1565__),
    .I1(__1643__),
    .I0(__1672__),
    .O(__2585__)
  );
  LUT6 #(
    .INIT(64'hfa000f0fcccccccc)
  ) __6269__ (
    .I5(__662__),
    .I4(__603__),
    .I3(__2585__),
    .I2(__2508__),
    .I1(__1194__),
    .I0(__2509__),
    .O(__2586__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __6270__ (
    .I3(__663__),
    .I2(__2282__),
    .I1(__1643__),
    .I0(__1279__),
    .O(__2587__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6271__ (
    .I2(__589__),
    .I1(__1865__),
    .I0(__723__),
    .O(__2588__)
  );
  LUT5 #(
    .INIT(32'ha000cccc)
  ) __6272__ (
    .I4(__662__),
    .I3(__1597__),
    .I2(__1596__),
    .I1(__784__),
    .I0(__1595__),
    .O(__2589__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6273__ (
    .I2(__589__),
    .I1(__2537__),
    .I0(__452__),
    .O(__2590__)
  );
  LUT6 #(
    .INIT(64'h8000000000000000)
  ) __6274__ (
    .I5(__646__),
    .I4(__656__),
    .I3(__657__),
    .I2(__658__),
    .I1(__2148__),
    .I0(__645__),
    .O(__2591__)
  );
  LUT6 #(
    .INIT(64'h0078787878787878)
  ) __6275__ (
    .I5(__589__),
    .I4(__1598__),
    .I3(__603__),
    .I2(__643__),
    .I1(__644__),
    .I0(__2591__),
    .O(__2592__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6276__ (
    .I2(__1511__),
    .I1(__127__),
    .I0(__105__),
    .O(__2593__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __6277__ (
    .I3(__662__),
    .I2(__603__),
    .I1(__1426__),
    .I0(__1314__),
    .O(__2594__)
  );
  LUT6 #(
    .INIT(64'h8000010000000000)
  ) __6278__ (
    .I5(__1682__),
    .I4(__1681__),
    .I3(__1680__),
    .I2(__1679__),
    .I1(__1678__),
    .I0(__1677__),
    .O(__2595__)
  );
  LUT6 #(
    .INIT(64'h9393399393939393)
  ) __6279__ (
    .I5(__1682__),
    .I4(__1681__),
    .I3(__1680__),
    .I2(__1686__),
    .I1(__1689__),
    .I0(__2595__),
    .O(__2596__)
  );
  LUT5 #(
    .INIT(32'h0fbb0f0f)
  ) __6280__ (
    .I4(__1732__),
    .I3(__1728__),
    .I2(__1411__),
    .I1(__2596__),
    .I0(__1697__),
    .O(__2597__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __6281__ (
    .I2(__663__),
    .I1(__2597__),
    .I0(__579__),
    .O(__2598__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __6282__ (
    .I3(__663__),
    .I2(__603__),
    .I1(__1438__),
    .I0(__845__),
    .O(__2599__)
  );
  LUT5 #(
    .INIT(32'h06666666)
  ) __6283__ (
    .I4(__589__),
    .I3(__1598__),
    .I2(__603__),
    .I1(__568__),
    .I0(__2149__),
    .O(__2600__)
  );
  LUT5 #(
    .INIT(32'hcd000000)
  ) __6284__ (
    .I4(__662__),
    .I3(__603__),
    .I2(__1570__),
    .I1(__2446__),
    .I0(__2445__),
    .O(__2601__)
  );
  LUT6 #(
    .INIT(64'hffff0707ff00ff00)
  ) __6285__ (
    .I5(__2601__),
    .I4(__1543__),
    .I3(__1156__),
    .I2(__2440__),
    .I1(__1542__),
    .I0(__2439__),
    .O(__2602__)
  );
  LUT5 #(
    .INIT(32'h21a522aa)
  ) __6286__ (
    .I4(__944__),
    .I3(__954__),
    .I2(__924__),
    .I1(__925__),
    .I0(__921__),
    .O(__2603__)
  );
  LUT6 #(
    .INIT(64'he4ee4e4e4eeee4e4)
  ) __6287__ (
    .I5(g3229),
    .I4(__1932__),
    .I3(__1929__),
    .I2(__1930__),
    .I1(__131__),
    .I0(__2173__),
    .O(__2604__)
  );
  LUT6 #(
    .INIT(64'h0000baaaaaaaaaaa)
  ) __6288__ (
    .I5(__944__),
    .I4(__875__),
    .I3(__93__),
    .I2(__73__),
    .I1(__748__),
    .I0(__757__),
    .O(__2605__)
  );
  LUT5 #(
    .INIT(32'ha000cccc)
  ) __6289__ (
    .I4(__954__),
    .I3(__1981__),
    .I2(__354__),
    .I1(__268__),
    .I0(__1800__),
    .O(__2606__)
  );
  LUT5 #(
    .INIT(32'h6c9ccccc)
  ) __6290__ (
    .I4(__1543__),
    .I3(__1544__),
    .I2(__1542__),
    .I1(__1538__),
    .I0(__1546__),
    .O(__2607__)
  );
  LUT6 #(
    .INIT(64'hf0f03355f0f0f0f0)
  ) __6291__ (
    .I5(__1592__),
    .I4(__1588__),
    .I3(__1555__),
    .I2(__1419__),
    .I1(__1545__),
    .I0(__2607__),
    .O(__2608__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6292__ (
    .I2(__663__),
    .I1(__2608__),
    .I0(__1273__),
    .O(__2609__)
  );
  LUT5 #(
    .INIT(32'hfcccaaaa)
  ) __6293__ (
    .I4(__944__),
    .I3(__862__),
    .I2(__868__),
    .I1(__1782__),
    .I0(__1373__),
    .O(__2610__)
  );
  LUT5 #(
    .INIT(32'h4ecccccc)
  ) __6294__ (
    .I4(__589__),
    .I3(__1598__),
    .I2(__1436__),
    .I1(__775__),
    .I0(__1635__),
    .O(__2611__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6295__ (
    .I2(__1511__),
    .I1(__117__),
    .I0(__193__),
    .O(__2612__)
  );
  LUT4 #(
    .INIT(16'h0080)
  ) __6296__ (
    .I3(__745__),
    .I2(__944__),
    .I1(__768__),
    .I0(__760__),
    .O(__2613__)
  );
  LUT4 #(
    .INIT(16'h125a)
  ) __6297__ (
    .I3(__954__),
    .I2(__767__),
    .I1(__752__),
    .I0(__2613__),
    .O(__2614__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __6298__ (
    .I5(__764__),
    .I4(__573__),
    .I3(__858__),
    .I2(__745__),
    .I1(__691__),
    .I0(__772__),
    .O(__2615__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6299__ (
    .I2(__589__),
    .I1(__2355__),
    .I0(__702__),
    .O(__2616__)
  );
  LUT5 #(
    .INIT(32'haa20cf45)
  ) __6300__ (
    .I4(g3229),
    .I3(__1602__),
    .I2(__1601__),
    .I1(__1600__),
    .I0(__1632__),
    .O(__2617__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6301__ (
    .I2(__1633__),
    .I1(__2617__),
    .I0(__1114__),
    .O(__2618__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __6302__ (
    .I1(__603__),
    .I0(__1570__),
    .O(__2619__)
  );
  LUT6 #(
    .INIT(64'hffff00ffd5ffd5d5)
  ) __6303__ (
    .I5(__1543__),
    .I4(__1544__),
    .I3(__1542__),
    .I2(__1585__),
    .I1(__1580__),
    .I0(__2619__),
    .O(__2620__)
  );
  LUT5 #(
    .INIT(32'h00008000)
  ) __6304__ (
    .I4(__1591__),
    .I3(__1574__),
    .I2(__1569__),
    .I1(__1564__),
    .I0(__1561__),
    .O(__2621__)
  );
  LUT4 #(
    .INIT(16'h11f0)
  ) __6305__ (
    .I3(__589__),
    .I2(__1168__),
    .I1(__2621__),
    .I0(__2620__),
    .O(__2622__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __6306__ (
    .I3(__589__),
    .I2(__603__),
    .I1(__1454__),
    .I0(__1328__),
    .O(__2623__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6307__ (
    .I2(__944__),
    .I1(__1647__),
    .I0(__748__),
    .O(__2624__)
  );
  LUT6 #(
    .INIT(64'h4545ff000505ff00)
  ) __6308__ (
    .I5(__858__),
    .I4(__954__),
    .I3(__120__),
    .I2(__1949__),
    .I1(__121__),
    .I0(__1624__),
    .O(__2625__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6309__ (
    .I2(__1511__),
    .I1(__123__),
    .I0(__83__),
    .O(__2626__)
  );
  LUT6 #(
    .INIT(64'h0000000f00000011)
  ) __6310__ (
    .I5(__988__),
    .I4(g563),
    .I3(__986__),
    .I2(__991__),
    .I1(__858__),
    .I0(__990__),
    .O(__2627__)
  );
  LUT4 #(
    .INIT(16'h8040)
  ) __6311__ (
    .I3(__2219__),
    .I2(__988__),
    .I1(__2627__),
    .I0(__1805__),
    .O(__2628__)
  );
  LUT3 #(
    .INIT(8'hf1)
  ) __6312__ (
    .I2(__1037__),
    .I1(__936__),
    .I0(__1036__),
    .O(__2629__)
  );
  LUT3 #(
    .INIT(8'hf1)
  ) __6313__ (
    .I2(__1036__),
    .I1(__936__),
    .I0(__1037__),
    .O(__2630__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __6314__ (
    .I5(__944__),
    .I4(__856__),
    .I3(__858__),
    .I2(__871__),
    .I1(__954__),
    .I0(__861__),
    .O(__2631__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6315__ (
    .I1(__2226__),
    .I0(__2222__),
    .O(__2632__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __6316__ (
    .I1(__2239__),
    .I0(__2234__),
    .O(__2633__)
  );
  LUT6 #(
    .INIT(64'h0000000000008000)
  ) __6317__ (
    .I5(__2225__),
    .I4(__2228__),
    .I3(__2219__),
    .I2(__2232__),
    .I1(__2633__),
    .I0(__2632__),
    .O(__2634__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __6318__ (
    .I5(__944__),
    .I4(__851__),
    .I3(__858__),
    .I2(__854__),
    .I1(__954__),
    .I0(__852__),
    .O(__2635__)
  );
  LUT5 #(
    .INIT(32'h00000008)
  ) __6319__ (
    .I4(__2635__),
    .I3(__2218__),
    .I2(__2220__),
    .I1(__2634__),
    .I0(__2230__),
    .O(__2636__)
  );
  LUT6 #(
    .INIT(64'h0000df0f00000000)
  ) __6320__ (
    .I5(__1037__),
    .I4(__1036__),
    .I3(__988__),
    .I2(__2627__),
    .I1(__2636__),
    .I0(__2631__),
    .O(__2637__)
  );
  LUT6 #(
    .INIT(64'hffffffff000f00bb)
  ) __6321__ (
    .I5(__2637__),
    .I4(__2630__),
    .I3(__2629__),
    .I2(__2628__),
    .I1(__2627__),
    .I0(__934__),
    .O(__2638__)
  );
  LUT6 #(
    .INIT(64'h0f007f00ff00ff00)
  ) __6322__ (
    .I5(__603__),
    .I4(__1570__),
    .I3(__1544__),
    .I2(__1542__),
    .I1(__1585__),
    .I0(__1580__),
    .O(__2639__)
  );
  LUT5 #(
    .INIT(32'hfcf9f0f0)
  ) __6323__ (
    .I4(__603__),
    .I3(__1570__),
    .I2(__1544__),
    .I1(__1542__),
    .I0(__2445__),
    .O(__2640__)
  );
  LUT5 #(
    .INIT(32'h000b0004)
  ) __6324__ (
    .I4(__1542__),
    .I3(__1543__),
    .I2(__2621__),
    .I1(__2640__),
    .I0(__2639__),
    .O(__2641__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6325__ (
    .I2(__589__),
    .I1(__2641__),
    .I0(__1158__),
    .O(__2642__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __6326__ (
    .I5(__954__),
    .I4(__242__),
    .I3(__370__),
    .I2(__229__),
    .I1(__255__),
    .I0(__366__),
    .O(__2643__)
  );
  LUT6 #(
    .INIT(64'h0100000100000000)
  ) __6327__ (
    .I5(__300__),
    .I4(__1982__),
    .I3(__1785__),
    .I2(__297__),
    .I1(g2637),
    .I0(__1784__),
    .O(__2644__)
  );
  LUT3 #(
    .INIT(8'hf1)
  ) __6328__ (
    .I2(__356__),
    .I1(__242__),
    .I0(__354__),
    .O(__2645__)
  );
  LUT3 #(
    .INIT(8'hf1)
  ) __6329__ (
    .I2(__354__),
    .I1(__242__),
    .I0(__356__),
    .O(__2646__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __6330__ (
    .I5(__944__),
    .I4(__147__),
    .I3(__858__),
    .I2(__146__),
    .I1(__954__),
    .I0(__248__),
    .O(__2647__)
  );
  LUT3 #(
    .INIT(8'h08)
  ) __6331__ (
    .I2(__1788__),
    .I1(__1798__),
    .I0(__1791__),
    .O(__2648__)
  );
  LUT6 #(
    .INIT(64'h0000df0f00000000)
  ) __6332__ (
    .I5(__356__),
    .I4(__354__),
    .I3(__300__),
    .I2(__1802__),
    .I1(__2648__),
    .I0(__2647__),
    .O(__2649__)
  );
  LUT6 #(
    .INIT(64'hffffffff000f00bb)
  ) __6333__ (
    .I5(__2649__),
    .I4(__2646__),
    .I3(__2645__),
    .I2(__2644__),
    .I1(__1802__),
    .I0(__239__),
    .O(__2650__)
  );
  LUT5 #(
    .INIT(32'he0000000)
  ) __6334__ (
    .I4(__1543__),
    .I3(__1542__),
    .I2(__1592__),
    .I1(__1554__),
    .I0(__1552__),
    .O(__2651__)
  );
  LUT5 #(
    .INIT(32'hdff72008)
  ) __6335__ (
    .I4(__1549__),
    .I3(__1537__),
    .I2(__1547__),
    .I1(__1545__),
    .I0(__1556__),
    .O(__2652__)
  );
  LUT6 #(
    .INIT(64'h01000f000f000f00)
  ) __6336__ (
    .I5(__1543__),
    .I4(__1542__),
    .I3(__1592__),
    .I2(__1588__),
    .I1(__1554__),
    .I0(__1552__),
    .O(__2653__)
  );
  LUT6 #(
    .INIT(64'h0f0f4444ff00ff00)
  ) __6337__ (
    .I5(__663__),
    .I4(__2653__),
    .I3(__1253__),
    .I2(__2652__),
    .I1(__1428__),
    .I0(__2651__),
    .O(__2654__)
  );
  LUT4 #(
    .INIT(16'haccc)
  ) __6338__ (
    .I3(__589__),
    .I2(__603__),
    .I1(__1292__),
    .I0(__1565__),
    .O(__2655__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __6339__ (
    .I5(__858__),
    .I4(__936__),
    .I3(__927__),
    .I2(__924__),
    .I1(__883__),
    .I0(__911__),
    .O(__2656__)
  );
  LUT6 #(
    .INIT(64'h8000000000000000)
  ) __6340__ (
    .I5(__1501__),
    .I4(__1502__),
    .I3(__1499__),
    .I2(__1500__),
    .I1(__1498__),
    .I0(__215__),
    .O(__2657__)
  );
  LUT6 #(
    .INIT(64'h0000000012305af0)
  ) __6341__ (
    .I5(g3234),
    .I4(__1623__),
    .I3(__1503__),
    .I2(__1504__),
    .I1(__215__),
    .I0(__2657__),
    .O(__2658__)
  );
  LUT5 #(
    .INIT(32'h77f0f0f0)
  ) __6342__ (
    .I4(__662__),
    .I3(__603__),
    .I2(__1153__),
    .I1(__1591__),
    .I0(__1575__),
    .O(__2659__)
  );
  LUT4 #(
    .INIT(16'he7ee)
  ) __6343__ (
    .I3(__1617__),
    .I2(__1614__),
    .I1(__2411__),
    .I0(__1613__),
    .O(__2660__)
  );
  LUT6 #(
    .INIT(64'h108000c000000000)
  ) __6344__ (
    .I5(__603__),
    .I4(__1617__),
    .I3(__2411__),
    .I2(__2410__),
    .I1(__1613__),
    .I0(__1614__),
    .O(__2661__)
  );
  LUT5 #(
    .INIT(32'h00f4f0f0)
  ) __6345__ (
    .I4(__589__),
    .I3(__2661__),
    .I2(__1119__),
    .I1(__603__),
    .I0(__2660__),
    .O(__2662__)
  );
  LUT6 #(
    .INIT(64'hfa000f0fcccccccc)
  ) __6346__ (
    .I5(__589__),
    .I4(__603__),
    .I3(__2585__),
    .I2(__2508__),
    .I1(__1193__),
    .I0(__2509__),
    .O(__2663__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __6347__ (
    .I5(__944__),
    .I4(__242__),
    .I3(__370__),
    .I2(__229__),
    .I1(__156__),
    .I0(__365__),
    .O(__2664__)
  );
  LUT4 #(
    .INIT(16'h0001)
  ) __6348__ (
    .I3(__2178__),
    .I2(__140__),
    .I1(g1249),
    .I0(__74__),
    .O(__2665__)
  );
  LUT6 #(
    .INIT(64'h0100000100000000)
  ) __6349__ (
    .I5(__142__),
    .I4(__2190__),
    .I3(__1951__),
    .I2(__2178__),
    .I1(__140__),
    .I0(g1249),
    .O(__2666__)
  );
  LUT6 #(
    .INIT(64'h0100000000000000)
  ) __6350__ (
    .I5(__2180__),
    .I4(__2190__),
    .I3(__2191__),
    .I2(__2193__),
    .I1(__2192__),
    .I0(__2195__),
    .O(__2667__)
  );
  LUT6 #(
    .INIT(64'h0000000000000008)
  ) __6351__ (
    .I5(__2188__),
    .I4(__2196__),
    .I3(__2197__),
    .I2(__2187__),
    .I1(__2185__),
    .I0(__2184__),
    .O(__2668__)
  );
  LUT4 #(
    .INIT(16'h0010)
  ) __6352__ (
    .I3(__2178__),
    .I2(__142__),
    .I1(__140__),
    .I0(g1249),
    .O(__2669__)
  );
  LUT5 #(
    .INIT(32'hf8070000)
  ) __6353__ (
    .I4(__2669__),
    .I3(__1951__),
    .I2(__2196__),
    .I1(__2668__),
    .I0(__2667__),
    .O(__2670__)
  );
  LUT5 #(
    .INIT(32'h00330f55)
  ) __6354__ (
    .I4(__2183__),
    .I3(__2182__),
    .I2(__2670__),
    .I1(__2666__),
    .I0(__2665__),
    .O(__2671__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __6355__ (
    .I2(__662__),
    .I1(__2556__),
    .I0(__441__),
    .O(__2672__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6356__ (
    .I2(__663__),
    .I1(__1733__),
    .I0(__455__),
    .O(__2673__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __6357__ (
    .I2(__663__),
    .I1(__2212__),
    .I0(__554__),
    .O(__2674__)
  );
  LUT6 #(
    .INIT(64'h0000baaaaaaaaaaa)
  ) __6358__ (
    .I5(__954__),
    .I4(__752__),
    .I3(__764__),
    .I2(__573__),
    .I1(__745__),
    .I0(__668__),
    .O(__2675__)
  );
  LUT5 #(
    .INIT(32'haa20cf45)
  ) __6359__ (
    .I4(g3229),
    .I3(__1930__),
    .I2(__1928__),
    .I1(__1932__),
    .I0(__1929__),
    .O(__2676__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6360__ (
    .I2(__2095__),
    .I1(__2676__),
    .I0(__136__),
    .O(__2677__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __6361__ (
    .I5(__944__),
    .I4(__1009__),
    .I3(__858__),
    .I2(__1008__),
    .I1(__954__),
    .I0(__1010__),
    .O(__2678__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __6362__ (
    .I5(__589__),
    .I4(__1196__),
    .I3(__663__),
    .I2(__1199__),
    .I1(__662__),
    .I0(__1197__),
    .O(__2679__)
  );
  LUT6 #(
    .INIT(64'hcc77f0f077ccf0f0)
  ) __6363__ (
    .I5(g3229),
    .I4(__2568__),
    .I3(__2065__),
    .I2(__1208__),
    .I1(__2063__),
    .I0(__2679__),
    .O(__2680__)
  );
  LUT4 #(
    .INIT(16'h11f0)
  ) __6364__ (
    .I3(__589__),
    .I2(__473__),
    .I1(__1778__),
    .I0(__1762__),
    .O(__2681__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __6365__ (
    .I1(__1494__),
    .I0(g51),
    .O(__2682__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __6366__ (
    .I2(g3229),
    .I1(__1058__),
    .I0(__1056__),
    .O(__2683__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6367__ (
    .I2(__1479__),
    .I1(__1477__),
    .I0(__1453__),
    .O(__2684__)
  );
  LUT6 #(
    .INIT(64'h9333363333333333)
  ) __6368__ (
    .I5(__1543__),
    .I4(__1544__),
    .I3(__1542__),
    .I2(__1538__),
    .I1(__1539__),
    .I0(__1546__),
    .O(__2685__)
  );
  LUT6 #(
    .INIT(64'hf0f033aaf0f0f0f0)
  ) __6369__ (
    .I5(__1592__),
    .I4(__1588__),
    .I3(__1555__),
    .I2(__1422__),
    .I1(__1545__),
    .I0(__2685__),
    .O(__2686__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6370__ (
    .I2(__663__),
    .I1(__2686__),
    .I0(__1270__),
    .O(__2687__)
  );
  LUT5 #(
    .INIT(32'h0030aaaa)
  ) __6371__ (
    .I4(__663__),
    .I3(__1760__),
    .I2(__1761__),
    .I1(__1759__),
    .I0(__196__),
    .O(__2688__)
  );
  LUT6 #(
    .INIT(64'hdffffff720000008)
  ) __6372__ (
    .I5(__1540__),
    .I4(__1550__),
    .I3(__1536__),
    .I2(__1548__),
    .I1(__1545__),
    .I0(__1656__),
    .O(__2689__)
  );
  LUT6 #(
    .INIT(64'h0f0f33550f0f0f0f)
  ) __6373__ (
    .I5(__1592__),
    .I4(__1588__),
    .I3(__1555__),
    .I2(__1572__),
    .I1(__1545__),
    .I0(__2689__),
    .O(__2690__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6374__ (
    .I2(__663__),
    .I1(__2690__),
    .I0(__1240__),
    .O(__2691__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __6375__ (
    .I3(__663__),
    .I2(__603__),
    .I1(__1454__),
    .I0(__1331__),
    .O(__2692__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __6376__ (
    .I5(__764__),
    .I4(__573__),
    .I3(__954__),
    .I2(__745__),
    .I1(__693__),
    .I0(__765__),
    .O(__2693__)
  );
  LUT6 #(
    .INIT(64'h3fffff3faaaaaaaa)
  ) __6377__ (
    .I5(__1807__),
    .I4(g3229),
    .I3(__1810__),
    .I2(__1809__),
    .I1(__1808__),
    .I0(__975__),
    .O(__2694__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6378__ (
    .I2(__944__),
    .I1(__2051__),
    .I0(__947__),
    .O(__2695__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __6379__ (
    .I5(__858__),
    .I4(__242__),
    .I3(__370__),
    .I2(__229__),
    .I1(__199__),
    .I0(__225__),
    .O(__2696__)
  );
  LUT5 #(
    .INIT(32'hcd000000)
  ) __6380__ (
    .I4(__663__),
    .I3(__603__),
    .I2(__1570__),
    .I1(__2446__),
    .I0(__2445__),
    .O(__2697__)
  );
  LUT6 #(
    .INIT(64'hffff0707ff00ff00)
  ) __6381__ (
    .I5(__2697__),
    .I4(__1543__),
    .I3(__1157__),
    .I2(__2440__),
    .I1(__1542__),
    .I0(__2439__),
    .O(__2698__)
  );
  LUT4 #(
    .INIT(16'h0666)
  ) __6382__ (
    .I3(__954__),
    .I2(__925__),
    .I1(__916__),
    .I0(__1868__),
    .O(__2699__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __6383__ (
    .I3(__589__),
    .I2(__603__),
    .I1(__1444__),
    .I0(__834__),
    .O(__2700__)
  );
  LUT5 #(
    .INIT(32'h80ef0000)
  ) __6384__ (
    .I4(__663__),
    .I3(__1598__),
    .I2(__1543__),
    .I1(__1544__),
    .I0(__1542__),
    .O(__2701__)
  );
  LUT6 #(
    .INIT(64'hcc77f0f077ccf0f0)
  ) __6385__ (
    .I5(g3229),
    .I4(__2701__),
    .I3(__2065__),
    .I2(__1209__),
    .I1(__2063__),
    .I0(__2679__),
    .O(__2702__)
  );
  LUT5 #(
    .INIT(32'ha000cccc)
  ) __6386__ (
    .I4(__858__),
    .I3(__1036__),
    .I2(__1806__),
    .I1(__942__),
    .I0(__1805__),
    .O(__2703__)
  );
  LUT5 #(
    .INIT(32'ha000cccc)
  ) __6387__ (
    .I4(__944__),
    .I3(__1951__),
    .I2(__2094__),
    .I1(__100__),
    .I0(__266__),
    .O(__2704__)
  );
  LUT5 #(
    .INIT(32'h0c66cccc)
  ) __6388__ (
    .I4(__589__),
    .I3(__1598__),
    .I2(__603__),
    .I1(__1178__),
    .I0(__1180__),
    .O(__2705__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6389__ (
    .I2(__954__),
    .I1(__300__),
    .I0(__1358__),
    .O(__2706__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __6390__ (
    .I5(__944__),
    .I4(__764__),
    .I3(__573__),
    .I2(__745__),
    .I1(__506__),
    .I0(__768__),
    .O(__2707__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __6391__ (
    .I1(__1537__),
    .I0(__1556__),
    .O(__2708__)
  );
  LUT6 #(
    .INIT(64'hf0f03355f0f0f0f0)
  ) __6392__ (
    .I5(__1592__),
    .I4(__1588__),
    .I3(__1555__),
    .I2(__1424__),
    .I1(__1545__),
    .I0(__2708__),
    .O(__2709__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6393__ (
    .I2(__663__),
    .I1(__2709__),
    .I0(__1267__),
    .O(__2710__)
  );
  LUT5 #(
    .INIT(32'hf8070000)
  ) __6394__ (
    .I4(__2669__),
    .I3(__1951__),
    .I2(__2192__),
    .I1(__2668__),
    .I0(__2667__),
    .O(__2711__)
  );
  LUT6 #(
    .INIT(64'h000033330f0faf00)
  ) __6395__ (
    .I5(__266__),
    .I4(__269__),
    .I3(__93__),
    .I2(__2179__),
    .I1(__2711__),
    .I0(__76__),
    .O(__2712__)
  );
  LUT6 #(
    .INIT(64'h8000000000000000)
  ) __6396__ (
    .I5(__2148__),
    .I4(__1232__),
    .I3(__1236__),
    .I2(__1235__),
    .I1(__1237__),
    .I0(__1234__),
    .O(__2713__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6397__ (
    .I1(__1228__),
    .I0(__2713__),
    .O(__2714__)
  );
  LUT6 #(
    .INIT(64'h00007fff00008000)
  ) __6398__ (
    .I5(__1220__),
    .I4(__2151__),
    .I3(__1222__),
    .I2(__1224__),
    .I1(__1223__),
    .I0(__2714__),
    .O(__2715__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6399__ (
    .I2(__589__),
    .I1(__1968__),
    .I0(__1241__),
    .O(__2716__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __6400__ (
    .I2(__662__),
    .I1(__1872__),
    .I0(__1275__),
    .O(__2717__)
  );
  LUT4 #(
    .INIT(16'haccc)
  ) __6401__ (
    .I3(__663__),
    .I2(__603__),
    .I1(__1294__),
    .I0(__1565__),
    .O(__2718__)
  );
  LUT6 #(
    .INIT(64'hf000b00000000000)
  ) __6402__ (
    .I5(__603__),
    .I4(__1570__),
    .I3(__1544__),
    .I2(__1542__),
    .I1(__1585__),
    .I0(__2445__),
    .O(__2719__)
  );
  LUT6 #(
    .INIT(64'hff5fffff2222ffff)
  ) __6403__ (
    .I5(__1544__),
    .I4(__1542__),
    .I3(__1587__),
    .I2(__1575__),
    .I1(__1585__),
    .I0(__1580__),
    .O(__2720__)
  );
  LUT6 #(
    .INIT(64'h00000000bfffffff)
  ) __6404__ (
    .I5(__1590__),
    .I4(__1574__),
    .I3(__1569__),
    .I2(__1564__),
    .I1(__1561__),
    .I0(__1587__),
    .O(__2721__)
  );
  LUT6 #(
    .INIT(64'hfafffaccfafffaff)
  ) __6405__ (
    .I5(__603__),
    .I4(__1570__),
    .I3(__1544__),
    .I2(__1542__),
    .I1(__1580__),
    .I0(__2721__),
    .O(__2722__)
  );
  LUT6 #(
    .INIT(64'h00ff000040400000)
  ) __6406__ (
    .I5(__1543__),
    .I4(__1544__),
    .I3(__1542__),
    .I2(__2722__),
    .I1(__2720__),
    .I0(__2719__),
    .O(__2723__)
  );
  LUT3 #(
    .INIT(8'h10)
  ) __6407__ (
    .I2(__603__),
    .I1(__1570__),
    .I0(__2445__),
    .O(__2724__)
  );
  LUT5 #(
    .INIT(32'h0000004f)
  ) __6408__ (
    .I4(__1543__),
    .I3(__1544__),
    .I2(__2722__),
    .I1(__2724__),
    .I0(__2720__),
    .O(__2725__)
  );
  LUT5 #(
    .INIT(32'h00eef0f0)
  ) __6409__ (
    .I4(__663__),
    .I3(__2621__),
    .I2(__1167__),
    .I1(__2725__),
    .I0(__2723__),
    .O(__2726__)
  );
  LUT6 #(
    .INIT(64'hf000b00000000000)
  ) __6410__ (
    .I5(__603__),
    .I4(__1757__),
    .I3(__1760__),
    .I2(__1759__),
    .I1(__1756__),
    .I0(__1997__),
    .O(__2727__)
  );
  LUT6 #(
    .INIT(64'hff5fffff2222ffff)
  ) __6411__ (
    .I5(__1760__),
    .I4(__1759__),
    .I3(__1860__),
    .I2(__1858__),
    .I1(__1756__),
    .I0(__1745__),
    .O(__2728__)
  );
  LUT6 #(
    .INIT(64'h00000000bfffffff)
  ) __6412__ (
    .I5(__1863__),
    .I4(__1776__),
    .I3(__1773__),
    .I2(__1769__),
    .I1(__1766__),
    .I0(__1860__),
    .O(__2729__)
  );
  LUT6 #(
    .INIT(64'hfafffaccfafffaff)
  ) __6413__ (
    .I5(__603__),
    .I4(__1757__),
    .I3(__1760__),
    .I2(__1759__),
    .I1(__1745__),
    .I0(__2729__),
    .O(__2730__)
  );
  LUT6 #(
    .INIT(64'h00ff000040400000)
  ) __6414__ (
    .I5(__1761__),
    .I4(__1760__),
    .I3(__1759__),
    .I2(__2730__),
    .I1(__2728__),
    .I0(__2727__),
    .O(__2731__)
  );
  LUT3 #(
    .INIT(8'h10)
  ) __6415__ (
    .I2(__603__),
    .I1(__1757__),
    .I0(__1997__),
    .O(__2732__)
  );
  LUT5 #(
    .INIT(32'h0000004f)
  ) __6416__ (
    .I4(__1761__),
    .I3(__1760__),
    .I2(__2730__),
    .I1(__2732__),
    .I0(__2728__),
    .O(__2733__)
  );
  LUT5 #(
    .INIT(32'h00eef0f0)
  ) __6417__ (
    .I4(__589__),
    .I3(__1778__),
    .I2(__418__),
    .I1(__2733__),
    .I0(__2731__),
    .O(__2734__)
  );
  LUT6 #(
    .INIT(64'h0000baaaaaaaaaaa)
  ) __6418__ (
    .I5(__944__),
    .I4(__231__),
    .I3(__242__),
    .I2(__370__),
    .I1(__229__),
    .I0(__245__),
    .O(__2735__)
  );
  LUT4 #(
    .INIT(16'h0006)
  ) __6419__ (
    .I3(__1497__),
    .I2(__1611__),
    .I1(__1489__),
    .I0(__1608__),
    .O(__2736__)
  );
  LUT5 #(
    .INIT(32'h00000708)
  ) __6420__ (
    .I4(__1497__),
    .I3(__1492__),
    .I2(__1611__),
    .I1(__1493__),
    .I0(__1494__),
    .O(__2737__)
  );
  LUT4 #(
    .INIT(16'haccc)
  ) __6421__ (
    .I3(__858__),
    .I2(__875__),
    .I1(__1364__),
    .I0(__2056__),
    .O(__2738__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6422__ (
    .I2(__663__),
    .I1(__2155__),
    .I0(__525__),
    .O(__2739__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __6423__ (
    .I2(g3229),
    .I1(__502__),
    .I0(__500__),
    .O(__2740__)
  );
  LUT5 #(
    .INIT(32'h4ecccccc)
  ) __6424__ (
    .I4(__663__),
    .I3(__1598__),
    .I2(__1407__),
    .I1(__623__),
    .I0(__1635__),
    .O(__2741__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __6425__ (
    .I1(__1686__),
    .I0(__2595__),
    .O(__2742__)
  );
  LUT6 #(
    .INIT(64'hf0f03355f0f0f0f0)
  ) __6426__ (
    .I5(__1732__),
    .I4(__1728__),
    .I3(__1697__),
    .I2(__1410__),
    .I1(__1684__),
    .I0(__2742__),
    .O(__2743__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6427__ (
    .I2(__662__),
    .I1(__2743__),
    .I0(__587__),
    .O(__2744__)
  );
  LUT6 #(
    .INIT(64'h0f0f4444ff00ff00)
  ) __6428__ (
    .I5(__663__),
    .I4(__2526__),
    .I3(__713__),
    .I2(__2525__),
    .I1(__1446__),
    .I0(__2524__),
    .O(__2745__)
  );
  LUT4 #(
    .INIT(16'h0080)
  ) __6429__ (
    .I3(__924__),
    .I2(__944__),
    .I1(__920__),
    .I0(__921__),
    .O(__2746__)
  );
  LUT5 #(
    .INIT(32'h12305af0)
  ) __6430__ (
    .I4(__954__),
    .I3(__918__),
    .I2(__917__),
    .I1(__925__),
    .I0(__2746__),
    .O(__2747__)
  );
  LUT6 #(
    .INIT(64'h4545ff000505ff00)
  ) __6431__ (
    .I5(__858__),
    .I4(__944__),
    .I3(__280__),
    .I2(__2117__),
    .I1(__282__),
    .I0(__1624__),
    .O(__2748__)
  );
  LUT4 #(
    .INIT(16'h0080)
  ) __6432__ (
    .I3(__924__),
    .I2(__954__),
    .I1(__936__),
    .I0(__927__),
    .O(__2749__)
  );
  LUT5 #(
    .INIT(32'h3f00aaaa)
  ) __6433__ (
    .I4(__2749__),
    .I3(__2240__),
    .I2(__2237__),
    .I1(__2224__),
    .I0(__861__),
    .O(__2750__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __6434__ (
    .I3(__589__),
    .I2(__2282__),
    .I1(__2140__),
    .I0(__751__),
    .O(__2751__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __6435__ (
    .I2(__662__),
    .I1(__2597__),
    .I0(__612__),
    .O(__2752__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __6436__ (
    .I3(__662__),
    .I2(__603__),
    .I1(__1457__),
    .I0(__1310__),
    .O(__2753__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __6437__ (
    .I5(__954__),
    .I4(__936__),
    .I3(__927__),
    .I2(__924__),
    .I1(__882__),
    .I0(__911__),
    .O(__2754__)
  );
  LUT6 #(
    .INIT(64'hfa000f0fcccccccc)
  ) __6438__ (
    .I5(__663__),
    .I4(__603__),
    .I3(__2512__),
    .I2(__2277__),
    .I1(__624__),
    .I0(__2278__),
    .O(__2755__)
  );
  LUT4 #(
    .INIT(16'h0080)
  ) __6439__ (
    .I3(__745__),
    .I2(__764__),
    .I1(__573__),
    .I0(__858__),
    .O(__2756__)
  );
  LUT5 #(
    .INIT(32'h3f00aaaa)
  ) __6440__ (
    .I4(__2756__),
    .I3(__1838__),
    .I2(__1835__),
    .I1(__1822__),
    .I0(__672__),
    .O(__2757__)
  );
  LUT5 #(
    .INIT(32'ha000cccc)
  ) __6441__ (
    .I4(__662__),
    .I3(__1761__),
    .I2(__1760__),
    .I1(__179__),
    .I0(__1759__),
    .O(__2758__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __6442__ (
    .I3(__662__),
    .I2(__603__),
    .I1(__1454__),
    .I0(__1330__),
    .O(__2759__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __6443__ (
    .I5(__764__),
    .I4(__573__),
    .I3(__858__),
    .I2(__745__),
    .I1(__740__),
    .I0(__760__),
    .O(__2760__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __6444__ (
    .I2(__589__),
    .I1(__2280__),
    .I0(__540__),
    .O(__2761__)
  );
  LUT6 #(
    .INIT(64'h0f007f00ff00ff00)
  ) __6445__ (
    .I5(__1595__),
    .I4(__1899__),
    .I3(__1596__),
    .I2(__603__),
    .I1(__1898__),
    .I0(__1887__),
    .O(__2762__)
  );
  LUT5 #(
    .INIT(32'hfcf9f0f0)
  ) __6446__ (
    .I4(__603__),
    .I3(__1899__),
    .I2(__1596__),
    .I1(__1595__),
    .I0(__1921__),
    .O(__2763__)
  );
  LUT5 #(
    .INIT(32'h00008000)
  ) __6447__ (
    .I4(__1972__),
    .I3(__1914__),
    .I2(__1910__),
    .I1(__1907__),
    .I0(__1903__),
    .O(__2764__)
  );
  LUT5 #(
    .INIT(32'h000b0004)
  ) __6448__ (
    .I4(__1595__),
    .I3(__1597__),
    .I2(__2764__),
    .I1(__2763__),
    .I0(__2762__),
    .O(__2765__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6449__ (
    .I2(__589__),
    .I1(__2765__),
    .I0(__1081__),
    .O(__2766__)
  );
  LUT5 #(
    .INIT(32'hf8070000)
  ) __6450__ (
    .I4(__2669__),
    .I3(__2056__),
    .I2(__2187__),
    .I1(__2668__),
    .I0(__2667__),
    .O(__2767__)
  );
  LUT6 #(
    .INIT(64'h000033330f0faf00)
  ) __6451__ (
    .I5(__266__),
    .I4(__269__),
    .I3(__93__),
    .I2(__2179__),
    .I1(__2767__),
    .I0(__84__),
    .O(__2768__)
  );
  LUT2 #(
    .INIT(4'hd)
  ) __6452__ (
    .I1(g3230),
    .I0(g3233),
    .O(__2769__)
  );
  LUT5 #(
    .INIT(32'ha000cccc)
  ) __6453__ (
    .I4(__858__),
    .I3(__968__),
    .I2(__1646__),
    .I1(__574__),
    .I0(__1648__),
    .O(__2770__)
  );
  LUT6 #(
    .INIT(64'hcc77f0f077ccf0f0)
  ) __6454__ (
    .I5(g3229),
    .I4(__2288__),
    .I3(__2287__),
    .I2(__559__),
    .I1(__2285__),
    .I0(__2369__),
    .O(__2771__)
  );
  LUT6 #(
    .INIT(64'hfa000f0fcccccccc)
  ) __6455__ (
    .I5(__662__),
    .I4(__603__),
    .I3(__2417__),
    .I2(__2248__),
    .I1(__1127__),
    .I0(__2247__),
    .O(__2772__)
  );
  LUT6 #(
    .INIT(64'haa3aaaaaaaaaaaaa)
  ) __6456__ (
    .I5(__858__),
    .I4(__93__),
    .I3(__748__),
    .I2(__73__),
    .I1(__747__),
    .I0(__734__),
    .O(__2773__)
  );
  LUT5 #(
    .INIT(32'h80ef0000)
  ) __6457__ (
    .I4(__589__),
    .I3(__1598__),
    .I2(__1761__),
    .I1(__1760__),
    .I0(__1759__),
    .O(__2774__)
  );
  LUT6 #(
    .INIT(64'h3fffff3faaaaaaaa)
  ) __6458__ (
    .I5(__2774__),
    .I4(g3229),
    .I3(__2070__),
    .I2(__2069__),
    .I1(__2068__),
    .I0(__625__),
    .O(__2775__)
  );
  LUT6 #(
    .INIT(64'haa3aaaaaaaaaaaaa)
  ) __6459__ (
    .I5(__944__),
    .I4(__93__),
    .I3(__748__),
    .I2(__73__),
    .I1(__788__),
    .I0(__1054__),
    .O(__2776__)
  );
  LUT5 #(
    .INIT(32'h12305af0)
  ) __6460__ (
    .I4(__954__),
    .I3(__916__),
    .I2(__915__),
    .I1(__925__),
    .I0(__1868__),
    .O(__2777__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __6461__ (
    .I5(__858__),
    .I4(__936__),
    .I3(__927__),
    .I2(__924__),
    .I1(__904__),
    .I0(__918__),
    .O(__2778__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6462__ (
    .I2(__1511__),
    .I1(__125__),
    .I0(__81__),
    .O(__2779__)
  );
  LUT5 #(
    .INIT(32'h12305af0)
  ) __6463__ (
    .I4(__954__),
    .I3(__796__),
    .I2(__788__),
    .I1(__875__),
    .I0(__1667__),
    .O(__2780__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __6464__ (
    .I2(__954__),
    .I1(__2503__),
    .I0(__205__),
    .O(__2781__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6465__ (
    .I2(__663__),
    .I1(__2176__),
    .I0(__444__),
    .O(__2782__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __6466__ (
    .I1(__1895__),
    .I0(__2325__),
    .O(__2783__)
  );
  LUT6 #(
    .INIT(64'hf0f03355f0f0f0f0)
  ) __6467__ (
    .I5(__2015__),
    .I4(__2012__),
    .I3(__2008__),
    .I2(__1456__),
    .I1(__2002__),
    .I0(__2783__),
    .O(__2784__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6468__ (
    .I2(__663__),
    .I1(__2784__),
    .I0(__728__),
    .O(__2785__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __6469__ (
    .I5(__764__),
    .I4(__573__),
    .I3(__954__),
    .I2(__745__),
    .I1(__697__),
    .I0(__750__),
    .O(__2786__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6470__ (
    .I2(__662__),
    .I1(__2765__),
    .I0(__1083__),
    .O(__2787__)
  );
  LUT5 #(
    .INIT(32'haa20cf45)
  ) __6471__ (
    .I4(g3229),
    .I3(__2070__),
    .I2(__2068__),
    .I1(__2069__),
    .I0(__2581__),
    .O(__2788__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6472__ (
    .I2(__2071__),
    .I1(__2788__),
    .I0(__636__),
    .O(__2789__)
  );
  LUT6 #(
    .INIT(64'h7878d27878787878)
  ) __6473__ (
    .I5(__1597__),
    .I4(__1596__),
    .I3(__1595__),
    .I2(__1890__),
    .I1(__1881__),
    .I0(__2362__),
    .O(__2790__)
  );
  LUT5 #(
    .INIT(32'hf011f0f0)
  ) __6474__ (
    .I4(__2015__),
    .I3(__2012__),
    .I2(__1460__),
    .I1(__2008__),
    .I0(__2790__),
    .O(__2791__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6475__ (
    .I2(__663__),
    .I1(__2791__),
    .I0(__1201__),
    .O(__2792__)
  );
  LUT4 #(
    .INIT(16'h11f0)
  ) __6476__ (
    .I3(__662__),
    .I2(__475__),
    .I1(__1778__),
    .I0(__1762__),
    .O(__2793__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __6477__ (
    .I3(__589__),
    .I2(__603__),
    .I1(__1459__),
    .I0(__652__),
    .O(__2794__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6478__ (
    .I2(__858__),
    .I1(__297__),
    .I0(__1384__),
    .O(__2795__)
  );
  LUT4 #(
    .INIT(16'h0baa)
  ) __6479__ (
    .I3(__858__),
    .I2(__1624__),
    .I1(__2023__),
    .I0(__955__),
    .O(__2796__)
  );
  LUT4 #(
    .INIT(16'h0080)
  ) __6480__ (
    .I3(__748__),
    .I2(__944__),
    .I1(__747__),
    .I0(__802__),
    .O(__2797__)
  );
  LUT4 #(
    .INIT(16'h125a)
  ) __6481__ (
    .I3(__954__),
    .I2(__799__),
    .I1(__875__),
    .I0(__2797__),
    .O(__2798__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __6482__ (
    .I3(__589__),
    .I2(__603__),
    .I1(__1436__),
    .I0(__846__),
    .O(__2799__)
  );
  LUT6 #(
    .INIT(64'h00007fff00008000)
  ) __6483__ (
    .I5(__1175__),
    .I4(__2151__),
    .I3(__2148__),
    .I2(__1178__),
    .I1(__1176__),
    .I0(__1180__),
    .O(__2800__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6484__ (
    .I2(__954__),
    .I1(__297__),
    .I0(__1383__),
    .O(__2801__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6485__ (
    .I2(__589__),
    .I1(__2484__),
    .I0(__717__),
    .O(__2802__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __6486__ (
    .I3(__663__),
    .I2(__603__),
    .I1(__1414__),
    .I0(__536__),
    .O(__2803__)
  );
  LUT5 #(
    .INIT(32'h4ecccccc)
  ) __6487__ (
    .I4(__663__),
    .I3(__1598__),
    .I2(__1453__),
    .I1(__1259__),
    .I0(__1635__),
    .O(__2804__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __6488__ (
    .I2(__944__),
    .I1(__1624__),
    .I0(__445__),
    .O(__2805__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __6489__ (
    .I3(__662__),
    .I2(__603__),
    .I1(__1409__),
    .I0(__485__),
    .O(__2806__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __6490__ (
    .I3(__589__),
    .I2(__603__),
    .I1(__1413__),
    .I0(__221__),
    .O(__2807__)
  );
  LUT6 #(
    .INIT(64'h000a000c00000000)
  ) __6491__ (
    .I5(__242__),
    .I4(g3229),
    .I3(__354__),
    .I2(__356__),
    .I1(__369__),
    .I0(__370__),
    .O(__2808__)
  );
  LUT3 #(
    .INIT(8'h07)
  ) __6492__ (
    .I2(__1789__),
    .I1(__1798__),
    .I0(__1791__),
    .O(__2809__)
  );
  LUT6 #(
    .INIT(64'h0001010000000000)
  ) __6493__ (
    .I5(__300__),
    .I4(__1800__),
    .I3(__2809__),
    .I2(__297__),
    .I1(g2637),
    .I0(__1784__),
    .O(__2810__)
  );
  LUT3 #(
    .INIT(8'h07)
  ) __6494__ (
    .I2(__1788__),
    .I1(__1798__),
    .I0(__1791__),
    .O(__2811__)
  );
  LUT6 #(
    .INIT(64'h0001010000000000)
  ) __6495__ (
    .I5(__300__),
    .I4(__1982__),
    .I3(__2811__),
    .I2(__297__),
    .I1(g2637),
    .I0(__1784__),
    .O(__2812__)
  );
  LUT5 #(
    .INIT(32'h70077777)
  ) __6496__ (
    .I4(__356__),
    .I3(__2812__),
    .I2(__2810__),
    .I1(__1802__),
    .I0(__2808__),
    .O(__2813__)
  );
  LUT3 #(
    .INIT(8'h07)
  ) __6497__ (
    .I2(__1787__),
    .I1(__1798__),
    .I0(__1791__),
    .O(__2814__)
  );
  LUT6 #(
    .INIT(64'h0001010000000000)
  ) __6498__ (
    .I5(__300__),
    .I4(__1982__),
    .I3(__2814__),
    .I2(__297__),
    .I1(g2637),
    .I0(__1784__),
    .O(__2815__)
  );
  LUT6 #(
    .INIT(64'h0100000100000000)
  ) __6499__ (
    .I5(__300__),
    .I4(__1800__),
    .I3(__1795__),
    .I2(__297__),
    .I1(g2637),
    .I0(__1784__),
    .O(__2816__)
  );
  LUT3 #(
    .INIT(8'h07)
  ) __6500__ (
    .I2(__1793__),
    .I1(__1798__),
    .I0(__1791__),
    .O(__2817__)
  );
  LUT6 #(
    .INIT(64'h0001010000000000)
  ) __6501__ (
    .I5(__300__),
    .I4(__1982__),
    .I3(__2817__),
    .I2(__297__),
    .I1(g2637),
    .I0(__1784__),
    .O(__2818__)
  );
  LUT4 #(
    .INIT(16'h6996)
  ) __6502__ (
    .I3(__2818__),
    .I2(__2816__),
    .I1(__2815__),
    .I0(__1801__),
    .O(__2819__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __6503__ (
    .I1(__1982__),
    .I0(__1785__),
    .O(__2820__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __6504__ (
    .I1(__1800__),
    .I0(__1786__),
    .O(__2821__)
  );
  LUT6 #(
    .INIT(64'h0001010000000000)
  ) __6505__ (
    .I5(__300__),
    .I4(__2821__),
    .I3(__2820__),
    .I2(__297__),
    .I1(g2637),
    .I0(__1784__),
    .O(__2822__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __6506__ (
    .I1(__1800__),
    .I0(__1796__),
    .O(__2823__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __6507__ (
    .I1(__1982__),
    .I0(__1797__),
    .O(__2824__)
  );
  LUT6 #(
    .INIT(64'hfffefeffffffffff)
  ) __6508__ (
    .I5(__300__),
    .I4(__2824__),
    .I3(__2823__),
    .I2(__297__),
    .I1(g2637),
    .I0(__1784__),
    .O(__2825__)
  );
  LUT5 #(
    .INIT(32'h7dd75555)
  ) __6509__ (
    .I4(__354__),
    .I3(__2825__),
    .I2(__2822__),
    .I1(__2819__),
    .I0(__2813__),
    .O(__2826__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6510__ (
    .I2(__1511__),
    .I1(__80__),
    .I0(__168__),
    .O(__2827__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __6511__ (
    .I1(__1461__),
    .I0(__1462__),
    .O(__2828__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __6512__ (
    .I1(__1463__),
    .I0(__1464__),
    .O(__2829__)
  );
  LUT6 #(
    .INIT(64'h6996966996696996)
  ) __6513__ (
    .I5(__1467__),
    .I4(__1465__),
    .I3(__1466__),
    .I2(__1468__),
    .I1(__2829__),
    .I0(__2828__),
    .O(__2830__)
  );
  LUT5 #(
    .INIT(32'hf0f06633)
  ) __6514__ (
    .I4(__1479__),
    .I3(__1349__),
    .I2(__1435__),
    .I1(__2830__),
    .I0(g3231),
    .O(__2831__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6515__ (
    .I2(__1479__),
    .I1(__1466__),
    .I0(__1409__),
    .O(__2832__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __6516__ (
    .I5(__944__),
    .I4(__936__),
    .I3(__927__),
    .I2(__924__),
    .I1(__890__),
    .I0(__914__),
    .O(__2833__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __6517__ (
    .I2(__662__),
    .I1(__1640__),
    .I0(__1009__),
    .O(__2834__)
  );
  LUT5 #(
    .INIT(32'h0030aaaa)
  ) __6518__ (
    .I4(__589__),
    .I3(__1596__),
    .I2(__1597__),
    .I1(__1595__),
    .I0(__433__),
    .O(__2835__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __6519__ (
    .I2(__663__),
    .I1(__2556__),
    .I0(__618__),
    .O(__2836__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __6520__ (
    .I3(__589__),
    .I2(__2282__),
    .I1(__1454__),
    .I0(__1229__),
    .O(__2837__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6521__ (
    .I2(__1479__),
    .I1(__1431__),
    .I0(__1471__),
    .O(__2838__)
  );
  LUT6 #(
    .INIT(64'h0078787878787878)
  ) __6522__ (
    .I5(__589__),
    .I4(__1598__),
    .I3(__603__),
    .I2(__1224__),
    .I1(__1228__),
    .I0(__2713__),
    .O(__2839__)
  );
  LUT6 #(
    .INIT(64'hbfffffffa0000000)
  ) __6523__ (
    .I5(__1188__),
    .I4(__662__),
    .I3(__603__),
    .I2(__2585__),
    .I1(__2509__),
    .I0(__2508__),
    .O(__2840__)
  );
  LUT5 #(
    .INIT(32'h77f0f0f0)
  ) __6524__ (
    .I4(__662__),
    .I3(__603__),
    .I2(__470__),
    .I1(__1731__),
    .I0(__1715__),
    .O(__2841__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __6525__ (
    .I3(__663__),
    .I2(__603__),
    .I1(__1426__),
    .I0(__1315__),
    .O(__2842__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __6526__ (
    .I3(__662__),
    .I2(__603__),
    .I1(__1458__),
    .I0(__1307__),
    .O(__2843__)
  );
  LUT6 #(
    .INIT(64'h0f0f4444ff00ff00)
  ) __6527__ (
    .I5(__589__),
    .I4(__2653__),
    .I3(__1251__),
    .I2(__2652__),
    .I1(__1428__),
    .I0(__2651__),
    .O(__2844__)
  );
  LUT6 #(
    .INIT(64'h0000077007700000)
  ) __6528__ (
    .I5(__1744__),
    .I4(__656__),
    .I3(__1741__),
    .I2(__641__),
    .I1(__1750__),
    .I0(__640__),
    .O(__2845__)
  );
  LUT6 #(
    .INIT(64'h00000eee0eee0000)
  ) __6529__ (
    .I5(__1748__),
    .I4(__642__),
    .I3(__1746__),
    .I2(__644__),
    .I1(__1750__),
    .I0(__640__),
    .O(__2846__)
  );
  LUT5 #(
    .INIT(32'heee0eeee)
  ) __6530__ (
    .I4(__1761__),
    .I3(__1760__),
    .I2(__1759__),
    .I1(__1737__),
    .I0(__645__),
    .O(__2847__)
  );
  LUT6 #(
    .INIT(64'h0000077707770000)
  ) __6531__ (
    .I5(__1753__),
    .I4(__646__),
    .I3(__1737__),
    .I2(__645__),
    .I1(__1735__),
    .I0(__658__),
    .O(__2848__)
  );
  LUT6 #(
    .INIT(64'h0e00000000000000)
  ) __6532__ (
    .I5(__2848__),
    .I4(__2847__),
    .I3(__2846__),
    .I2(__1598__),
    .I1(__1746__),
    .I0(__644__),
    .O(__2849__)
  );
  LUT4 #(
    .INIT(16'h0ee0)
  ) __6533__ (
    .I3(__1739__),
    .I2(__643__),
    .I1(__1735__),
    .I0(__658__),
    .O(__2850__)
  );
  LUT6 #(
    .INIT(64'h155555559fffffff)
  ) __6534__ (
    .I5(__1857__),
    .I4(__2850__),
    .I3(__2849__),
    .I2(__2845__),
    .I1(__657__),
    .I0(__1755__),
    .O(__2851__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __6535__ (
    .I5(__944__),
    .I4(__242__),
    .I3(__370__),
    .I2(__229__),
    .I1(__172__),
    .I0(__222__),
    .O(__2852__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6536__ (
    .I2(__662__),
    .I1(__2641__),
    .I0(__1159__),
    .O(__2853__)
  );
  LUT4 #(
    .INIT(16'h25aa)
  ) __6537__ (
    .I3(__589__),
    .I2(__1598__),
    .I1(__603__),
    .I0(__658__),
    .O(__2854__)
  );
  LUT5 #(
    .INIT(32'h0030aaaa)
  ) __6538__ (
    .I4(__662__),
    .I3(__1682__),
    .I2(__1681__),
    .I1(__1680__),
    .I0(__151__),
    .O(__2855__)
  );
  LUT5 #(
    .INIT(32'hcd000000)
  ) __6539__ (
    .I4(__589__),
    .I3(__603__),
    .I2(__1710__),
    .I1(__2263__),
    .I0(__2262__),
    .O(__2856__)
  );
  LUT6 #(
    .INIT(64'hffff0707ff00ff00)
  ) __6540__ (
    .I5(__2856__),
    .I4(__1682__),
    .I3(__421__),
    .I2(__2257__),
    .I1(__1680__),
    .I0(__2256__),
    .O(__2857__)
  );
  LUT5 #(
    .INIT(32'h4ecccccc)
  ) __6541__ (
    .I4(__662__),
    .I3(__1598__),
    .I2(__1417__),
    .I1(__1281__),
    .I0(__1635__),
    .O(__2858__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6542__ (
    .I2(__954__),
    .I1(__868__),
    .I0(__1361__),
    .O(__2859__)
  );
  LUT6 #(
    .INIT(64'haa3aaaaaaaaaaaaa)
  ) __6543__ (
    .I5(__954__),
    .I4(__93__),
    .I3(__748__),
    .I2(__73__),
    .I1(__802__),
    .I0(__1421__),
    .O(__2860__)
  );
  LUT6 #(
    .INIT(64'hbfffffffa0000000)
  ) __6544__ (
    .I5(__1189__),
    .I4(__663__),
    .I3(__603__),
    .I2(__2585__),
    .I1(__2509__),
    .I0(__2508__),
    .O(__2861__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __6545__ (
    .I5(__764__),
    .I4(__573__),
    .I3(__858__),
    .I2(__745__),
    .I1(__694__),
    .I0(__765__),
    .O(__2862__)
  );
  LUT5 #(
    .INIT(32'h12305af0)
  ) __6546__ (
    .I4(__954__),
    .I3(__750__),
    .I2(__765__),
    .I1(__752__),
    .I0(__1985__),
    .O(__2863__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6547__ (
    .I2(__662__),
    .I1(__2784__),
    .I0(__726__),
    .O(__2864__)
  );
  LUT5 #(
    .INIT(32'he0000000)
  ) __6548__ (
    .I4(__1682__),
    .I3(__1680__),
    .I2(__1732__),
    .I1(__1696__),
    .I0(__1694__),
    .O(__2865__)
  );
  LUT5 #(
    .INIT(32'hdff72008)
  ) __6549__ (
    .I4(__1691__),
    .I3(__1686__),
    .I2(__1689__),
    .I1(__1684__),
    .I0(__2595__),
    .O(__2866__)
  );
  LUT6 #(
    .INIT(64'h01000f000f000f00)
  ) __6550__ (
    .I5(__1682__),
    .I4(__1680__),
    .I3(__1732__),
    .I2(__1728__),
    .I1(__1696__),
    .I0(__1694__),
    .O(__2867__)
  );
  LUT6 #(
    .INIT(64'h0f0f4444ff00ff00)
  ) __6551__ (
    .I5(__663__),
    .I4(__2867__),
    .I3(__446__),
    .I2(__2866__),
    .I1(__1412__),
    .I0(__2865__),
    .O(__2868__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __6552__ (
    .I5(__944__),
    .I4(__435__),
    .I3(__858__),
    .I2(__416__),
    .I1(__954__),
    .I0(__423__),
    .O(__2869__)
  );
  LUT5 #(
    .INIT(32'h80ef0000)
  ) __6553__ (
    .I4(__663__),
    .I3(__1598__),
    .I2(__1597__),
    .I1(__1596__),
    .I0(__1595__),
    .O(__2870__)
  );
  LUT6 #(
    .INIT(64'hd8fad850d850d8fa)
  ) __6554__ (
    .I5(g3229),
    .I4(__1602__),
    .I3(__1601__),
    .I2(__1137__),
    .I1(__1600__),
    .I0(__2870__),
    .O(__2871__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __6555__ (
    .I5(__954__),
    .I4(__936__),
    .I3(__927__),
    .I2(__924__),
    .I1(__909__),
    .I0(__921__),
    .O(__2872__)
  );
  LUT6 #(
    .INIT(64'haa3aaaaaaaaaaaaa)
  ) __6556__ (
    .I5(__858__),
    .I4(__93__),
    .I3(__748__),
    .I2(__73__),
    .I1(__796__),
    .I0(__1398__),
    .O(__2873__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6557__ (
    .I2(__1511__),
    .I1(__82__),
    .I0(__155__),
    .O(__2874__)
  );
  LUT6 #(
    .INIT(64'h0100000000000000)
  ) __6558__ (
    .I5(__2219__),
    .I4(__2232__),
    .I3(__2230__),
    .I2(__2225__),
    .I1(__2228__),
    .I0(__2635__),
    .O(__2875__)
  );
  LUT6 #(
    .INIT(64'h0000000000000008)
  ) __6559__ (
    .I5(__2239__),
    .I4(__2218__),
    .I3(__2220__),
    .I2(__2234__),
    .I1(__2226__),
    .I0(__2222__),
    .O(__2876__)
  );
  LUT6 #(
    .INIT(64'hf087000000000000)
  ) __6560__ (
    .I5(__988__),
    .I4(__2627__),
    .I3(__2234__),
    .I2(__1674__),
    .I1(__2876__),
    .I0(__2875__),
    .O(__2877__)
  );
  LUT6 #(
    .INIT(64'h000033330f0faf00)
  ) __6561__ (
    .I5(__1036__),
    .I4(__1037__),
    .I3(__936__),
    .I2(__2627__),
    .I1(__2877__),
    .I0(__931__),
    .O(__2878__)
  );
  LUT5 #(
    .INIT(32'h12305af0)
  ) __6562__ (
    .I4(__954__),
    .I3(__741__),
    .I2(__770__),
    .I1(__752__),
    .I0(__1986__),
    .O(__2879__)
  );
  LUT4 #(
    .INIT(16'h25aa)
  ) __6563__ (
    .I3(__589__),
    .I2(__1598__),
    .I1(__603__),
    .I0(__1237__),
    .O(__2880__)
  );
  LUT5 #(
    .INIT(32'haa20cf45)
  ) __6564__ (
    .I4(g3229),
    .I3(__2065__),
    .I2(__2064__),
    .I1(__2063__),
    .I0(__2679__),
    .O(__2881__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6565__ (
    .I2(__2062__),
    .I1(__2881__),
    .I0(__1214__),
    .O(__2882__)
  );
  LUT6 #(
    .INIT(64'haa3aaaaaaaaaaaaa)
  ) __6566__ (
    .I5(__944__),
    .I4(__93__),
    .I3(__748__),
    .I2(__73__),
    .I1(__1051__),
    .I0(__1399__),
    .O(__2883__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __6567__ (
    .I3(__662__),
    .I2(__2282__),
    .I1(__1643__),
    .I0(__1278__),
    .O(__2884__)
  );
  LUT6 #(
    .INIT(64'h7878d27878787878)
  ) __6568__ (
    .I5(__1543__),
    .I4(__1544__),
    .I3(__1542__),
    .I2(__1550__),
    .I1(__1548__),
    .I0(__1656__),
    .O(__2885__)
  );
  LUT5 #(
    .INIT(32'hf011f0f0)
  ) __6569__ (
    .I4(__1592__),
    .I3(__1588__),
    .I2(__1432__),
    .I1(__1555__),
    .I0(__2885__),
    .O(__2886__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6570__ (
    .I2(__662__),
    .I1(__2886__),
    .I0(__1246__),
    .O(__2887__)
  );
  LUT6 #(
    .INIT(64'h9393399393939393)
  ) __6571__ (
    .I5(__1761__),
    .I4(__1760__),
    .I3(__1759__),
    .I2(__1753__),
    .I1(__1737__),
    .I0(__2482__),
    .O(__2888__)
  );
  LUT5 #(
    .INIT(32'h0fbb0f0f)
  ) __6572__ (
    .I4(__1864__),
    .I3(__1861__),
    .I2(__1444__),
    .I1(__2888__),
    .I0(__1857__),
    .O(__2889__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __6573__ (
    .I2(__663__),
    .I1(__2889__),
    .I0(__716__),
    .O(__2890__)
  );
  LUT5 #(
    .INIT(32'h4ecccccc)
  ) __6574__ (
    .I4(__589__),
    .I3(__1598__),
    .I2(__1408__),
    .I1(__461__),
    .I0(__1635__),
    .O(__2891__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __6575__ (
    .I3(__662__),
    .I2(__603__),
    .I1(__1412__),
    .I0(__344__),
    .O(__2892__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __6576__ (
    .I2(__944__),
    .I1(__1624__),
    .I0(__357__),
    .O(__2893__)
  );
  LUT6 #(
    .INIT(64'h0100000100000000)
  ) __6577__ (
    .I5(__300__),
    .I4(__1800__),
    .I3(__1796__),
    .I2(__297__),
    .I1(g2637),
    .I0(__1784__),
    .O(__2894__)
  );
  LUT6 #(
    .INIT(64'hffffffff000f00bb)
  ) __6578__ (
    .I5(__2649__),
    .I4(__2646__),
    .I3(__2645__),
    .I2(__2894__),
    .I1(__1802__),
    .I0(__375__),
    .O(__2895__)
  );
  LUT6 #(
    .INIT(64'h000a000c00000000)
  ) __6579__ (
    .I5(__936__),
    .I4(g3229),
    .I3(__1037__),
    .I2(__1036__),
    .I1(__926__),
    .I0(__927__),
    .O(__2896__)
  );
  LUT4 #(
    .INIT(16'h8040)
  ) __6580__ (
    .I3(__2230__),
    .I2(__988__),
    .I1(__2627__),
    .I0(__1674__),
    .O(__2897__)
  );
  LUT4 #(
    .INIT(16'h8040)
  ) __6581__ (
    .I3(__2222__),
    .I2(__988__),
    .I1(__2627__),
    .I0(__1674__),
    .O(__2898__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6582__ (
    .I1(__988__),
    .I0(__2627__),
    .O(__2899__)
  );
  LUT6 #(
    .INIT(64'h5a5aa55aa55a5a5a)
  ) __6583__ (
    .I5(__2219__),
    .I4(__2226__),
    .I3(__2899__),
    .I2(__2898__),
    .I1(__1805__),
    .I0(__2897__),
    .O(__2900__)
  );
  LUT6 #(
    .INIT(64'hf087000000000000)
  ) __6584__ (
    .I5(__988__),
    .I4(__2627__),
    .I3(__2225__),
    .I2(__1674__),
    .I1(__2876__),
    .I0(__2875__),
    .O(__2901__)
  );
  LUT4 #(
    .INIT(16'h8040)
  ) __6585__ (
    .I3(__2232__),
    .I2(__988__),
    .I1(__2627__),
    .I0(__1805__),
    .O(__2902__)
  );
  LUT6 #(
    .INIT(64'hf087000000000000)
  ) __6586__ (
    .I5(__988__),
    .I4(__2627__),
    .I3(__2228__),
    .I2(__1805__),
    .I1(__2876__),
    .I0(__2875__),
    .O(__2903__)
  );
  LUT6 #(
    .INIT(64'h9669699600000000)
  ) __6587__ (
    .I5(__1036__),
    .I4(__2903__),
    .I3(__2902__),
    .I2(__2901__),
    .I1(__2877__),
    .I0(__2900__),
    .O(__2904__)
  );
  LUT5 #(
    .INIT(32'ha9000000)
  ) __6588__ (
    .I4(__988__),
    .I3(__2627__),
    .I2(__2220__),
    .I1(__2636__),
    .I0(__1674__),
    .O(__2905__)
  );
  LUT5 #(
    .INIT(32'ha9000000)
  ) __6589__ (
    .I4(__988__),
    .I3(__2627__),
    .I2(__2218__),
    .I1(__2636__),
    .I0(__1805__),
    .O(__2906__)
  );
  LUT6 #(
    .INIT(64'hf8fffff8f8f8f8f8)
  ) __6590__ (
    .I5(__1037__),
    .I4(__2906__),
    .I3(__2905__),
    .I2(__2904__),
    .I1(__2627__),
    .I0(__2896__),
    .O(__2907__)
  );
  LUT5 #(
    .INIT(32'h0000125a)
  ) __6591__ (
    .I4(g3234),
    .I3(__1623__),
    .I2(__1503__),
    .I1(__215__),
    .I0(__2657__),
    .O(__2908__)
  );
  LUT6 #(
    .INIT(64'h3fffff3faaaaaaaa)
  ) __6592__ (
    .I5(__2134__),
    .I4(g3229),
    .I3(__1810__),
    .I2(__1809__),
    .I1(__1808__),
    .I0(__974__),
    .O(__2909__)
  );
  LUT6 #(
    .INIT(64'h0000baaaaaaaaaaa)
  ) __6593__ (
    .I5(__944__),
    .I4(__752__),
    .I3(__764__),
    .I2(__573__),
    .I1(__745__),
    .I0(__667__),
    .O(__2910__)
  );
  LUT4 #(
    .INIT(16'haccc)
  ) __6594__ (
    .I3(__589__),
    .I2(__603__),
    .I1(__785__),
    .I0(__1884__),
    .O(__2911__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __6595__ (
    .I3(__662__),
    .I2(__603__),
    .I1(__1455__),
    .I0(__1326__),
    .O(__2912__)
  );
  LUT5 #(
    .INIT(32'hccaa0f0f)
  ) __6596__ (
    .I4(__383__),
    .I3(__662__),
    .I2(__337__),
    .I1(__2161__),
    .I0(__362__),
    .O(__2913__)
  );
  LUT5 #(
    .INIT(32'hccaa0f0f)
  ) __6597__ (
    .I4(__1057__),
    .I3(__662__),
    .I2(__1027__),
    .I1(__2913__),
    .I0(__1056__),
    .O(__2914__)
  );
  LUT6 #(
    .INIT(64'hf000f0ccaaaaaaaa)
  ) __6598__ (
    .I5(__944__),
    .I4(__858__),
    .I3(__988__),
    .I2(__991__),
    .I1(__990__),
    .I0(__1379__),
    .O(__2915__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __6599__ (
    .I3(__663__),
    .I2(__603__),
    .I1(__1424__),
    .I0(__1318__),
    .O(__2916__)
  );
  LUT4 #(
    .INIT(16'haccc)
  ) __6600__ (
    .I3(__663__),
    .I2(__603__),
    .I1(__819__),
    .I0(__1751__),
    .O(__2917__)
  );
  LUT5 #(
    .INIT(32'h77f0f0f0)
  ) __6601__ (
    .I4(__663__),
    .I3(__603__),
    .I2(__1154__),
    .I1(__1591__),
    .I0(__1575__),
    .O(__2918__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6602__ (
    .I2(__1511__),
    .I1(__96__),
    .I0(__164__),
    .O(__2919__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __6603__ (
    .I3(__662__),
    .I2(__603__),
    .I1(__1459__),
    .I0(__1301__),
    .O(__2920__)
  );
  LUT6 #(
    .INIT(64'h00000000007f0080)
  ) __6604__ (
    .I5(__1497__),
    .I4(__1488__),
    .I3(__1611__),
    .I2(__1489__),
    .I1(__1490__),
    .I0(__2498__),
    .O(__2921__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __6605__ (
    .I3(__663__),
    .I2(__603__),
    .I1(__1436__),
    .I0(__849__),
    .O(__2922__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __6606__ (
    .I2(__589__),
    .I1(__2279__),
    .I0(__183__),
    .O(__2923__)
  );
  LUT6 #(
    .INIT(64'h8000000000000000)
  ) __6607__ (
    .I5(__2148__),
    .I4(__1174__),
    .I3(__1178__),
    .I2(__1176__),
    .I1(__1180__),
    .I0(__1175__),
    .O(__2924__)
  );
  LUT6 #(
    .INIT(64'h0078787878787878)
  ) __6608__ (
    .I5(__589__),
    .I4(__1598__),
    .I3(__603__),
    .I2(__730__),
    .I1(__1164__),
    .I0(__2924__),
    .O(__2925__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __6609__ (
    .I5(__858__),
    .I4(__936__),
    .I3(__927__),
    .I2(__924__),
    .I1(__892__),
    .I0(__914__),
    .O(__2926__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __6610__ (
    .I3(__589__),
    .I2(__603__),
    .I1(__1455__),
    .I0(__1325__),
    .O(__2927__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __6611__ (
    .I2(__944__),
    .I1(__357__),
    .I0(__356__),
    .O(__2928__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6612__ (
    .I2(__1479__),
    .I1(__1451__),
    .I0(__1461__),
    .O(__2929__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __6613__ (
    .I2(__663__),
    .I1(__2510__),
    .I0(__1192__),
    .O(__2930__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6614__ (
    .I2(__954__),
    .I1(__1784__),
    .I0(__1371__),
    .O(__2931__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6615__ (
    .I2(__662__),
    .I1(__2686__),
    .I0(__1269__),
    .O(__2932__)
  );
  LUT6 #(
    .INIT(64'hfa000f0fcccccccc)
  ) __6616__ (
    .I5(__589__),
    .I4(__603__),
    .I3(__2512__),
    .I2(__2277__),
    .I1(__615__),
    .I0(__2278__),
    .O(__2933__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __6617__ (
    .I2(__589__),
    .I1(__1657__),
    .I0(__1248__),
    .O(__2934__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __6618__ (
    .I2(__589__),
    .I1(__2597__),
    .I0(__519__),
    .O(__2935__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __6619__ (
    .I2(__662__),
    .I1(__2290__),
    .I0(__517__),
    .O(__2936__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __6620__ (
    .I1(__1532__),
    .I0(__1522__),
    .O(__2937__)
  );
  LUT4 #(
    .INIT(16'h0001)
  ) __6621__ (
    .I3(__1351__),
    .I2(__1350__),
    .I1(__1349__),
    .I0(__1352__),
    .O(__2938__)
  );
  LUT4 #(
    .INIT(16'h0001)
  ) __6622__ (
    .I3(__1355__),
    .I2(__1356__),
    .I1(__1353__),
    .I0(__1354__),
    .O(__2939__)
  );
  LUT5 #(
    .INIT(32'h00000010)
  ) __6623__ (
    .I4(__1352__),
    .I3(__1355__),
    .I2(__1354__),
    .I1(__1356__),
    .I0(__1353__),
    .O(__2940__)
  );
  LUT4 #(
    .INIT(16'h0008)
  ) __6624__ (
    .I3(__1351__),
    .I2(__1349__),
    .I1(__1350__),
    .I0(__2940__),
    .O(__2941__)
  );
  LUT3 #(
    .INIT(8'h10)
  ) __6625__ (
    .I2(__1350__),
    .I1(__1351__),
    .I0(__1349__),
    .O(__2942__)
  );
  LUT3 #(
    .INIT(8'h10)
  ) __6626__ (
    .I2(__1349__),
    .I1(__1351__),
    .I0(__1350__),
    .O(__2943__)
  );
  LUT4 #(
    .INIT(16'h0010)
  ) __6627__ (
    .I3(__1355__),
    .I2(__1354__),
    .I1(__1356__),
    .I0(__1353__),
    .O(__2944__)
  );
  LUT6 #(
    .INIT(64'h0777ffffffffffff)
  ) __6628__ (
    .I5(__1352__),
    .I4(__2944__),
    .I3(__1372__),
    .I2(__2943__),
    .I1(__2942__),
    .I0(__1371__),
    .O(__2945__)
  );
  LUT6 #(
    .INIT(64'h00bfbfbf00000000)
  ) __6629__ (
    .I5(__2945__),
    .I4(__1379__),
    .I3(__2941__),
    .I2(__2939__),
    .I1(__2938__),
    .I0(__2937__),
    .O(__2946__)
  );
  LUT6 #(
    .INIT(64'h0000000000000008)
  ) __6630__ (
    .I5(__1355__),
    .I4(__1356__),
    .I3(__1353__),
    .I2(__1354__),
    .I1(__1352__),
    .I0(__2942__),
    .O(__2947__)
  );
  LUT6 #(
    .INIT(64'h0000000000000008)
  ) __6631__ (
    .I5(__1351__),
    .I4(__1350__),
    .I3(__1349__),
    .I2(__1352__),
    .I1(__1381__),
    .I0(__2944__),
    .O(__2948__)
  );
  LUT3 #(
    .INIT(8'h08)
  ) __6632__ (
    .I2(__1350__),
    .I1(__1351__),
    .I0(__1349__),
    .O(__2949__)
  );
  LUT3 #(
    .INIT(8'h08)
  ) __6633__ (
    .I2(__1351__),
    .I1(__1350__),
    .I0(__1349__),
    .O(__2950__)
  );
  LUT6 #(
    .INIT(64'h0fff7777ffffffff)
  ) __6634__ (
    .I5(__2944__),
    .I4(__1352__),
    .I3(__2950__),
    .I2(__1370__),
    .I1(__1376__),
    .I0(__2949__),
    .O(__2951__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __6635__ (
    .I1(__1350__),
    .I0(__1349__),
    .O(__2952__)
  );
  LUT6 #(
    .INIT(64'hf53fffffffffffff)
  ) __6636__ (
    .I5(__2944__),
    .I4(__2952__),
    .I3(__1351__),
    .I2(__1352__),
    .I1(__1373__),
    .I0(__1377__),
    .O(__2953__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6637__ (
    .I1(__1350__),
    .I0(__1349__),
    .O(__2954__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __6638__ (
    .I1(__1349__),
    .I0(__1350__),
    .O(__2955__)
  );
  LUT6 #(
    .INIT(64'hffffffff13ff5fff)
  ) __6639__ (
    .I5(__1351__),
    .I4(__2955__),
    .I3(__2940__),
    .I2(__2954__),
    .I1(__1380__),
    .I0(__1378__),
    .O(__2956__)
  );
  LUT6 #(
    .INIT(64'h0b00000000000000)
  ) __6640__ (
    .I5(__2956__),
    .I4(__2953__),
    .I3(__2951__),
    .I2(__2948__),
    .I1(__2947__),
    .I0(__1346__),
    .O(__2957__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __6641__ (
    .I1(__1350__),
    .I0(__1349__),
    .O(__2958__)
  );
  LUT6 #(
    .INIT(64'h0777ffffffffffff)
  ) __6642__ (
    .I5(__1351__),
    .I4(__2940__),
    .I3(__1374__),
    .I2(__2954__),
    .I1(__2958__),
    .I0(__1375__),
    .O(__2959__)
  );
  LUT6 #(
    .INIT(64'h00001f5f0000ffff)
  ) __6643__ (
    .I5(__1351__),
    .I4(__2769__),
    .I3(__1352__),
    .I2(__2939__),
    .I1(__2958__),
    .I0(__2952__),
    .O(__2960__)
  );
  LUT4 #(
    .INIT(16'h7fff)
  ) __6644__ (
    .I3(__2960__),
    .I2(__2959__),
    .I1(__2957__),
    .I0(__2946__),
    .O(__2961__)
  );
  LUT5 #(
    .INIT(32'haa20cf45)
  ) __6645__ (
    .I4(g3229),
    .I3(__1810__),
    .I2(__1809__),
    .I1(__1808__),
    .I0(__2030__),
    .O(__2962__)
  );
  LUT4 #(
    .INIT(16'haccc)
  ) __6646__ (
    .I3(__858__),
    .I2(__2429__),
    .I1(__985__),
    .I0(__2962__),
    .O(__2963__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6647__ (
    .I2(__662__),
    .I1(__2412__),
    .I0(__532__),
    .O(__2964__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6648__ (
    .I2(__858__),
    .I1(__988__),
    .I0(__1369__),
    .O(__2965__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __6649__ (
    .I5(__858__),
    .I4(__936__),
    .I3(__927__),
    .I2(__924__),
    .I1(__907__),
    .I0(__920__),
    .O(__2966__)
  );
  LUT5 #(
    .INIT(32'h00f4f0f0)
  ) __6650__ (
    .I4(__589__),
    .I3(__2405__),
    .I2(__1171__),
    .I1(__603__),
    .I0(__2404__),
    .O(__2967__)
  );
  LUT5 #(
    .INIT(32'ha000cccc)
  ) __6651__ (
    .I4(__954__),
    .I3(__1036__),
    .I2(__1806__),
    .I1(__941__),
    .I0(__1805__),
    .O(__2968__)
  );
  LUT4 #(
    .INIT(16'haccc)
  ) __6652__ (
    .I3(__663__),
    .I2(__603__),
    .I1(__376__),
    .I0(__1712__),
    .O(__2969__)
  );
  LUT6 #(
    .INIT(64'h4f0f4f0000000000)
  ) __6653__ (
    .I5(__954__),
    .I4(__2056__),
    .I3(__2094__),
    .I2(__1647__),
    .I1(__266__),
    .I0(__1951__),
    .O(__2970__)
  );
  LUT6 #(
    .INIT(64'he4ee4e4e4eeee4e4)
  ) __6654__ (
    .I5(g3229),
    .I4(__1932__),
    .I3(__1929__),
    .I2(__1930__),
    .I1(__130__),
    .I0(__2970__),
    .O(__2971__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6655__ (
    .I2(__1479__),
    .I1(__1445__),
    .I0(__1464__),
    .O(__2972__)
  );
  LUT3 #(
    .INIT(8'h70)
  ) __6656__ (
    .I2(__2394__),
    .I1(__858__),
    .I0(__814__),
    .O(__2973__)
  );
  LUT6 #(
    .INIT(64'h5455555555555555)
  ) __6657__ (
    .I5(__1623__),
    .I4(__1506__),
    .I3(__1505__),
    .I2(__1508__),
    .I1(__1507__),
    .I0(__1649__),
    .O(__2974__)
  );
  LUT6 #(
    .INIT(64'h0f080f0f0f0f0f0f)
  ) __6658__ (
    .I5(__2395__),
    .I4(__2385__),
    .I3(__2380__),
    .I2(__2974__),
    .I1(__2973__),
    .I0(__2391__),
    .O(__2975__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __6659__ (
    .I2(__858__),
    .I1(__2975__),
    .I0(__806__),
    .O(__2976__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __6660__ (
    .I3(__589__),
    .I2(__603__),
    .I1(__1419__),
    .I0(__1322__),
    .O(__2977__)
  );
  LUT6 #(
    .INIT(64'h4000000000000000)
  ) __6661__ (
    .I5(__589__),
    .I4(__646__),
    .I3(__656__),
    .I2(__657__),
    .I1(__658__),
    .I0(__1598__),
    .O(__2978__)
  );
  LUT5 #(
    .INIT(32'h06666666)
  ) __6662__ (
    .I4(__589__),
    .I3(__1598__),
    .I2(__603__),
    .I1(__645__),
    .I0(__2978__),
    .O(__2979__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __6663__ (
    .I5(__944__),
    .I4(__936__),
    .I3(__927__),
    .I2(__924__),
    .I1(__881__),
    .I0(__911__),
    .O(__2980__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6664__ (
    .I2(__1479__),
    .I1(__1462__),
    .I0(__1413__),
    .O(__2981__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6665__ (
    .I2(__662__),
    .I1(__2364__),
    .I0(__1173__),
    .O(__2982__)
  );
  LUT6 #(
    .INIT(64'hbfffffffa0000000)
  ) __6666__ (
    .I5(__595__),
    .I4(__589__),
    .I3(__603__),
    .I2(__2462__),
    .I1(__2210__),
    .I0(__2209__),
    .O(__2983__)
  );
  LUT6 #(
    .INIT(64'h4545ff000505ff00)
  ) __6667__ (
    .I5(__858__),
    .I4(__954__),
    .I3(__972__),
    .I2(__2048__),
    .I1(__973__),
    .I0(__1624__),
    .O(__2984__)
  );
  LUT4 #(
    .INIT(16'haccc)
  ) __6668__ (
    .I3(__944__),
    .I2(__231__),
    .I1(__304__),
    .I0(__1800__),
    .O(__2985__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __6669__ (
    .I3(__662__),
    .I2(__2282__),
    .I1(__2140__),
    .I0(__753__),
    .O(__2986__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __6670__ (
    .I5(__764__),
    .I4(__573__),
    .I3(__954__),
    .I2(__745__),
    .I1(__686__),
    .I0(__741__),
    .O(__2987__)
  );
  LUT5 #(
    .INIT(32'h00f4f0f0)
  ) __6671__ (
    .I4(__663__),
    .I3(__2661__),
    .I2(__648__),
    .I1(__603__),
    .I0(__2660__),
    .O(__2988__)
  );
  LUT6 #(
    .INIT(64'hcc77f0f077ccf0f0)
  ) __6672__ (
    .I5(g3229),
    .I4(__2071__),
    .I3(__2070__),
    .I2(__630__),
    .I1(__2069__),
    .I0(__2581__),
    .O(__2989__)
  );
  LUT6 #(
    .INIT(64'hfd75a820df578a02)
  ) __6673__ (
    .I5(g3229),
    .I4(__634__),
    .I3(__2069__),
    .I2(__2070__),
    .I1(__2068__),
    .I0(__2582__),
    .O(__2990__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __6674__ (
    .I5(__858__),
    .I4(__242__),
    .I3(__370__),
    .I2(__229__),
    .I1(__363__),
    .I0(__367__),
    .O(__2991__)
  );
  LUT6 #(
    .INIT(64'h4000000000000000)
  ) __6675__ (
    .I5(__589__),
    .I4(__571__),
    .I3(__606__),
    .I2(__607__),
    .I1(__570__),
    .I0(__1598__),
    .O(__2992__)
  );
  LUT5 #(
    .INIT(32'h06666666)
  ) __6676__ (
    .I4(__589__),
    .I3(__1598__),
    .I2(__603__),
    .I1(__514__),
    .I0(__2992__),
    .O(__2993__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6677__ (
    .I2(__1479__),
    .I1(__1463__),
    .I0(__1412__),
    .O(__2994__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __6678__ (
    .I3(__662__),
    .I2(__2282__),
    .I1(__1617__),
    .I0(__1261__),
    .O(__2995__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __6679__ (
    .I2(__662__),
    .I1(__2889__),
    .I0(__715__),
    .O(__2996__)
  );
  LUT6 #(
    .INIT(64'h0000baaaaaaaaaaa)
  ) __6680__ (
    .I5(__954__),
    .I4(__925__),
    .I3(__936__),
    .I2(__927__),
    .I1(__924__),
    .I0(__852__),
    .O(__2997__)
  );
  LUT6 #(
    .INIT(64'h00f07878f0f0f0f0)
  ) __6681__ (
    .I5(__589__),
    .I4(__1598__),
    .I3(__603__),
    .I2(__1235__),
    .I1(__1236__),
    .I0(__1237__),
    .O(__2998__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __6682__ (
    .I1(__603__),
    .I0(__1899__),
    .O(__2999__)
  );
  LUT6 #(
    .INIT(64'hffff00ffd5ffd5d5)
  ) __6683__ (
    .I5(__1597__),
    .I4(__1596__),
    .I3(__1595__),
    .I2(__1898__),
    .I1(__1887__),
    .I0(__2999__),
    .O(__3000__)
  );
  LUT4 #(
    .INIT(16'h11f0)
  ) __6684__ (
    .I3(__589__),
    .I2(__850__),
    .I1(__2764__),
    .I0(__3000__),
    .O(__3001__)
  );
  LUT5 #(
    .INIT(32'haa20cf45)
  ) __6685__ (
    .I4(g3229),
    .I3(__1653__),
    .I2(__1651__),
    .I1(__1652__),
    .I0(__2269__),
    .O(__3002__)
  );
  LUT6 #(
    .INIT(64'h4f0f4f0000000000)
  ) __6686__ (
    .I5(__858__),
    .I4(__1649__),
    .I3(__1648__),
    .I2(__1647__),
    .I1(__968__),
    .I0(__1646__),
    .O(__3003__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6687__ (
    .I2(__3003__),
    .I1(__3002__),
    .I0(__866__),
    .O(__3004__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __6688__ (
    .I1(__603__),
    .I0(__1710__),
    .O(__3005__)
  );
  LUT6 #(
    .INIT(64'hffff00ffd5ffd5d5)
  ) __6689__ (
    .I5(__1682__),
    .I4(__1681__),
    .I3(__1680__),
    .I2(__1725__),
    .I1(__1720__),
    .I0(__3005__),
    .O(__3006__)
  );
  LUT5 #(
    .INIT(32'h00008000)
  ) __6690__ (
    .I4(__1731__),
    .I3(__1714__),
    .I2(__1709__),
    .I1(__1704__),
    .I0(__1701__),
    .O(__3007__)
  );
  LUT4 #(
    .INIT(16'h11f0)
  ) __6691__ (
    .I3(__589__),
    .I2(__161__),
    .I1(__3007__),
    .I0(__3006__),
    .O(__3008__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __6692__ (
    .I3(__663__),
    .I2(__603__),
    .I1(__1432__),
    .I0(__1297__),
    .O(__3009__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6693__ (
    .I2(__1479__),
    .I1(__1420__),
    .I0(__1476__),
    .O(__3010__)
  );
  LUT6 #(
    .INIT(64'hcc77f0f077ccf0f0)
  ) __6694__ (
    .I5(g3229),
    .I4(__2244__),
    .I3(__1979__),
    .I2(__289__),
    .I1(__1977__),
    .I0(__1976__),
    .O(__3011__)
  );
  LUT6 #(
    .INIT(64'h5555cffc55555555)
  ) __6695__ (
    .I5(__2015__),
    .I4(__2012__),
    .I3(__1881__),
    .I2(__2362__),
    .I1(__2008__),
    .I0(__1459__),
    .O(__3012__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __6696__ (
    .I2(__589__),
    .I1(__3012__),
    .I0(__1202__),
    .O(__3013__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __6697__ (
    .I5(__944__),
    .I4(__1003__),
    .I3(__858__),
    .I2(__1002__),
    .I1(__954__),
    .I0(__1004__),
    .O(__3014__)
  );
  LUT6 #(
    .INIT(64'h0100000100000000)
  ) __6698__ (
    .I5(__300__),
    .I4(__1982__),
    .I3(__1797__),
    .I2(__297__),
    .I1(g2637),
    .I0(__1784__),
    .O(__3015__)
  );
  LUT6 #(
    .INIT(64'h000000004fff0000)
  ) __6699__ (
    .I5(__354__),
    .I4(__356__),
    .I3(__300__),
    .I2(__1802__),
    .I1(__2647__),
    .I0(__2648__),
    .O(__3016__)
  );
  LUT6 #(
    .INIT(64'hffffffff000f00bb)
  ) __6700__ (
    .I5(__3016__),
    .I4(__2646__),
    .I3(__2645__),
    .I2(__3015__),
    .I1(__1802__),
    .I0(__240__),
    .O(__3017__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6701__ (
    .I2(__1479__),
    .I1(__1433__),
    .I0(__1470__),
    .O(__3018__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __6702__ (
    .I2(__663__),
    .I1(__2411__),
    .I0(__431__),
    .O(__3019__)
  );
  LUT5 #(
    .INIT(32'h00eef0f0)
  ) __6703__ (
    .I4(__662__),
    .I3(__1778__),
    .I2(__469__),
    .I1(__2733__),
    .I0(__2731__),
    .O(__3020__)
  );
  LUT6 #(
    .INIT(64'hd8fad850d850d8fa)
  ) __6704__ (
    .I5(g3229),
    .I4(__1653__),
    .I3(__1651__),
    .I2(__825__),
    .I1(__1652__),
    .I0(__3003__),
    .O(__3021__)
  );
  LUT4 #(
    .INIT(16'haccc)
  ) __6705__ (
    .I3(__954__),
    .I2(__925__),
    .I1(__879__),
    .I0(__1805__),
    .O(__3022__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __6706__ (
    .I2(g3229),
    .I1(__384__),
    .I0(__362__),
    .O(__3023__)
  );
  LUT4 #(
    .INIT(16'haccc)
  ) __6707__ (
    .I3(__954__),
    .I2(__925__),
    .I1(__876__),
    .I0(__1674__),
    .O(__3024__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __6708__ (
    .I3(__589__),
    .I2(__603__),
    .I1(__1411__),
    .I0(__639__),
    .O(__3025__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __6709__ (
    .I2(__662__),
    .I1(__2211__),
    .I0(__149__),
    .O(__3026__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __6710__ (
    .I2(__589__),
    .I1(__2889__),
    .I0(__714__),
    .O(__3027__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __6711__ (
    .I5(__858__),
    .I4(__936__),
    .I3(__927__),
    .I2(__924__),
    .I1(__898__),
    .I0(__916__),
    .O(__3028__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __6712__ (
    .I5(__764__),
    .I4(__573__),
    .I3(__954__),
    .I2(__745__),
    .I1(__680__),
    .I0(__749__),
    .O(__3029__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __6713__ (
    .I3(__662__),
    .I2(__603__),
    .I1(__1428__),
    .I0(__1303__),
    .O(__3030__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6714__ (
    .I2(__589__),
    .I1(__2784__),
    .I0(__1045__),
    .O(__3031__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __6715__ (
    .I5(__944__),
    .I4(__1000__),
    .I3(__858__),
    .I2(__999__),
    .I1(__954__),
    .I0(__1001__),
    .O(__3032__)
  );
  LUT6 #(
    .INIT(64'he4ee4e4e4eeee4e4)
  ) __6716__ (
    .I5(g3229),
    .I4(__1932__),
    .I3(__1929__),
    .I2(__1930__),
    .I1(__128__),
    .I0(__2095__),
    .O(__3033__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6717__ (
    .I2(__954__),
    .I1(__2178__),
    .I0(__1377__),
    .O(__3034__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __6718__ (
    .I5(__944__),
    .I4(__936__),
    .I3(__927__),
    .I2(__924__),
    .I1(__908__),
    .I0(__921__),
    .O(__3035__)
  );
  LUT5 #(
    .INIT(32'h4ecccccc)
  ) __6719__ (
    .I4(__589__),
    .I3(__1598__),
    .I2(__1419__),
    .I1(__1283__),
    .I0(__1635__),
    .O(__3036__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __6720__ (
    .I3(__663__),
    .I2(__603__),
    .I1(__1444__),
    .I0(__836__),
    .O(__3037__)
  );
  LUT5 #(
    .INIT(32'ha000cccc)
  ) __6721__ (
    .I4(__663__),
    .I3(__1682__),
    .I2(__1681__),
    .I1(__311__),
    .I0(__1680__),
    .O(__3038__)
  );
  LUT5 #(
    .INIT(32'h77f0f0f0)
  ) __6722__ (
    .I4(__589__),
    .I3(__603__),
    .I2(__1073__),
    .I1(__1972__),
    .I0(__2011__),
    .O(__3039__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6723__ (
    .I2(__2582__),
    .I1(__2788__),
    .I0(__637__),
    .O(__3040__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __6724__ (
    .I3(__589__),
    .I2(__603__),
    .I1(__1438__),
    .I0(__843__),
    .O(__3041__)
  );
  LUT6 #(
    .INIT(64'h000033330f0faf00)
  ) __6725__ (
    .I5(__354__),
    .I4(__356__),
    .I3(__242__),
    .I2(__1802__),
    .I1(__2815__),
    .I0(__236__),
    .O(__3042__)
  );
  LUT5 #(
    .INIT(32'hfcccaaaa)
  ) __6726__ (
    .I4(__858__),
    .I3(__862__),
    .I2(__868__),
    .I1(__1782__),
    .I0(__1375__),
    .O(__3043__)
  );
  LUT4 #(
    .INIT(16'haccc)
  ) __6727__ (
    .I3(__663__),
    .I2(__603__),
    .I1(__792__),
    .I0(__1884__),
    .O(__3044__)
  );
  LUT6 #(
    .INIT(64'hcc77f0f077ccf0f0)
  ) __6728__ (
    .I5(g3229),
    .I4(__1599__),
    .I3(__1602__),
    .I2(__1132__),
    .I1(__1600__),
    .I0(__1632__),
    .O(__3045__)
  );
  LUT5 #(
    .INIT(32'hcd000000)
  ) __6729__ (
    .I4(__663__),
    .I3(__603__),
    .I2(__1899__),
    .I1(__1922__),
    .I0(__1921__),
    .O(__3046__)
  );
  LUT6 #(
    .INIT(64'hffff0707ff00ff00)
  ) __6730__ (
    .I5(__3046__),
    .I4(__1597__),
    .I3(__1080__),
    .I2(__1916__),
    .I1(__1595__),
    .I0(__1915__),
    .O(__3047__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __6731__ (
    .I5(__858__),
    .I4(__242__),
    .I3(__370__),
    .I2(__229__),
    .I1(__177__),
    .I0(__222__),
    .O(__3048__)
  );
  LUT6 #(
    .INIT(64'h4f0f4f0000000000)
  ) __6732__ (
    .I5(__944__),
    .I4(__1982__),
    .I3(__1981__),
    .I2(__1647__),
    .I1(__354__),
    .I0(__1800__),
    .O(__3049__)
  );
  LUT6 #(
    .INIT(64'hcc77f0f077ccf0f0)
  ) __6733__ (
    .I5(g3229),
    .I4(__3049__),
    .I3(__1979__),
    .I2(__287__),
    .I1(__1977__),
    .I0(__1976__),
    .O(__3050__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6734__ (
    .I2(__663__),
    .I1(__2484__),
    .I0(__719__),
    .O(__3051__)
  );
  LUT6 #(
    .INIT(64'h4545ff000505ff00)
  ) __6735__ (
    .I5(__858__),
    .I4(__944__),
    .I3(__561__),
    .I2(__2394__),
    .I1(__814__),
    .I0(__1624__),
    .O(__3052__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __6736__ (
    .I3(__663__),
    .I2(__603__),
    .I1(__1409__),
    .I0(__538__),
    .O(__3053__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __6737__ (
    .I2(__663__),
    .I1(__3012__),
    .I0(__1205__),
    .O(__3054__)
  );
  LUT4 #(
    .INIT(16'hfbfe)
  ) __6738__ (
    .I3(__1493__),
    .I2(__1497__),
    .I1(__1494__),
    .I0(__1611__),
    .O(__3055__)
  );
  LUT6 #(
    .INIT(64'h0f007f00ff00ff00)
  ) __6739__ (
    .I5(__603__),
    .I4(__1710__),
    .I3(__1681__),
    .I2(__1680__),
    .I1(__1725__),
    .I0(__1720__),
    .O(__3056__)
  );
  LUT5 #(
    .INIT(32'hfcf9f0f0)
  ) __6740__ (
    .I4(__603__),
    .I3(__1710__),
    .I2(__1681__),
    .I1(__1680__),
    .I0(__2262__),
    .O(__3057__)
  );
  LUT5 #(
    .INIT(32'h000b0004)
  ) __6741__ (
    .I4(__1680__),
    .I3(__1682__),
    .I2(__3007__),
    .I1(__3057__),
    .I0(__3056__),
    .O(__3058__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6742__ (
    .I2(__663__),
    .I1(__3058__),
    .I0(__457__),
    .O(__3059__)
  );
  LUT6 #(
    .INIT(64'hfd75a820df578a02)
  ) __6743__ (
    .I5(g3229),
    .I4(__1212__),
    .I3(__2063__),
    .I2(__2065__),
    .I1(__2064__),
    .I0(__2701__),
    .O(__3060__)
  );
  LUT6 #(
    .INIT(64'h7878d27878787878)
  ) __6744__ (
    .I5(__1682__),
    .I4(__1681__),
    .I3(__1680__),
    .I2(__1692__),
    .I1(__1690__),
    .I0(__1960__),
    .O(__3061__)
  );
  LUT5 #(
    .INIT(32'hf011f0f0)
  ) __6745__ (
    .I4(__1732__),
    .I3(__1728__),
    .I2(__1414__),
    .I1(__1697__),
    .I0(__3061__),
    .O(__3062__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6746__ (
    .I2(__663__),
    .I1(__3062__),
    .I0(__584__),
    .O(__3063__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __6747__ (
    .I2(__663__),
    .I1(__1672__),
    .I0(__1001__),
    .O(__3064__)
  );
  LUT6 #(
    .INIT(64'hcc77f0f077ccf0f0)
  ) __6748__ (
    .I5(g3229),
    .I4(__2489__),
    .I3(__1810__),
    .I2(__979__),
    .I1(__1808__),
    .I0(__2030__),
    .O(__3065__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __6749__ (
    .I2(__1623__),
    .I1(__1505__),
    .I0(__215__),
    .O(__3066__)
  );
  LUT5 #(
    .INIT(32'h007d0080)
  ) __6750__ (
    .I4(__1508__),
    .I3(g3234),
    .I2(__1506__),
    .I1(__1507__),
    .I0(__3066__),
    .O(__3067__)
  );
  LUT5 #(
    .INIT(32'h00eef0f0)
  ) __6751__ (
    .I4(__663__),
    .I3(__1778__),
    .I2(__472__),
    .I1(__2733__),
    .I0(__2731__),
    .O(__3068__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __6752__ (
    .I2(__662__),
    .I1(__1957__),
    .I0(__474__),
    .O(__3069__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6753__ (
    .I2(__662__),
    .I1(__3062__),
    .I0(__610__),
    .O(__3070__)
  );
  LUT6 #(
    .INIT(64'h3fffff3faaaaaaaa)
  ) __6754__ (
    .I5(__2568__),
    .I4(g3229),
    .I3(__2065__),
    .I2(__2063__),
    .I1(__2064__),
    .I0(__1197__),
    .O(__3071__)
  );
  LUT6 #(
    .INIT(64'hf000b00000000000)
  ) __6755__ (
    .I5(__603__),
    .I4(__1710__),
    .I3(__1681__),
    .I2(__1680__),
    .I1(__1725__),
    .I0(__2262__),
    .O(__3072__)
  );
  LUT6 #(
    .INIT(64'hff5fffff2222ffff)
  ) __6756__ (
    .I5(__1681__),
    .I4(__1680__),
    .I3(__1727__),
    .I2(__1715__),
    .I1(__1725__),
    .I0(__1720__),
    .O(__3073__)
  );
  LUT6 #(
    .INIT(64'h00000000bfffffff)
  ) __6757__ (
    .I5(__1730__),
    .I4(__1714__),
    .I3(__1709__),
    .I2(__1704__),
    .I1(__1701__),
    .I0(__1727__),
    .O(__3074__)
  );
  LUT6 #(
    .INIT(64'hfafffaccfafffaff)
  ) __6758__ (
    .I5(__603__),
    .I4(__1710__),
    .I3(__1681__),
    .I2(__1680__),
    .I1(__1720__),
    .I0(__3074__),
    .O(__3075__)
  );
  LUT6 #(
    .INIT(64'h00ff000040400000)
  ) __6759__ (
    .I5(__1682__),
    .I4(__1681__),
    .I3(__1680__),
    .I2(__3075__),
    .I1(__3073__),
    .I0(__3072__),
    .O(__3076__)
  );
  LUT3 #(
    .INIT(8'h10)
  ) __6760__ (
    .I2(__603__),
    .I1(__1710__),
    .I0(__2262__),
    .O(__3077__)
  );
  LUT5 #(
    .INIT(32'h0000004f)
  ) __6761__ (
    .I4(__1682__),
    .I3(__1681__),
    .I2(__3075__),
    .I1(__3077__),
    .I0(__3073__),
    .O(__3078__)
  );
  LUT5 #(
    .INIT(32'h00eef0f0)
  ) __6762__ (
    .I4(__663__),
    .I3(__3007__),
    .I2(__160__),
    .I1(__3078__),
    .I0(__3076__),
    .O(__3079__)
  );
  LUT6 #(
    .INIT(64'h132033005fa0ff00)
  ) __6763__ (
    .I5(__954__),
    .I4(__913__),
    .I3(__911__),
    .I2(__912__),
    .I1(__925__),
    .I0(__1869__),
    .O(__3080__)
  );
  LUT6 #(
    .INIT(64'h0100000100000000)
  ) __6764__ (
    .I5(__868__),
    .I4(__1646__),
    .I3(__1830__),
    .I2(__1966__),
    .I1(g1943),
    .I0(__867__),
    .O(__3081__)
  );
  LUT5 #(
    .INIT(32'h003300af)
  ) __6765__ (
    .I4(__2348__),
    .I3(__2347__),
    .I2(__2346__),
    .I1(__3081__),
    .I0(__755__),
    .O(__3082__)
  );
  LUT3 #(
    .INIT(8'h07)
  ) __6766__ (
    .I2(__1816__),
    .I1(__2343__),
    .I0(__2342__),
    .O(__3083__)
  );
  LUT6 #(
    .INIT(64'haaaaaaaaeafabafa)
  ) __6767__ (
    .I5(__968__),
    .I4(__1646__),
    .I3(__2344__),
    .I2(__969__),
    .I1(__3083__),
    .I0(__3082__),
    .O(__3084__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __6768__ (
    .I3(__663__),
    .I2(__603__),
    .I1(__1457__),
    .I0(__1311__),
    .O(__3085__)
  );
  LUT6 #(
    .INIT(64'hfa000f0fcccccccc)
  ) __6769__ (
    .I5(__663__),
    .I4(__603__),
    .I3(__2462__),
    .I2(__2209__),
    .I1(__556__),
    .I0(__2210__),
    .O(__3086__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __6770__ (
    .I1(__1472__),
    .I0(__1471__),
    .O(__3087__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __6771__ (
    .I1(__1473__),
    .I0(__1470__),
    .O(__3088__)
  );
  LUT6 #(
    .INIT(64'h6996966996696996)
  ) __6772__ (
    .I5(__1475__),
    .I4(__1474__),
    .I3(__1476__),
    .I2(__1477__),
    .I1(__3088__),
    .I0(__3087__),
    .O(__3089__)
  );
  LUT5 #(
    .INIT(32'h3c33aaaa)
  ) __6773__ (
    .I4(__1479__),
    .I3(__1349__),
    .I2(g3231),
    .I1(__3089__),
    .I0(__1452__),
    .O(__3090__)
  );
  LUT5 #(
    .INIT(32'h3c33aaaa)
  ) __6774__ (
    .I4(__1479__),
    .I3(__1349__),
    .I2(g3231),
    .I1(__2830__),
    .I0(__1405__),
    .O(__3091__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __6775__ (
    .I5(__944__),
    .I4(__764__),
    .I3(__573__),
    .I2(__745__),
    .I1(__705__),
    .I0(__767__),
    .O(__3092__)
  );
  LUT4 #(
    .INIT(16'h125a)
  ) __6776__ (
    .I3(__954__),
    .I2(__750__),
    .I1(__752__),
    .I0(__1985__),
    .O(__3093__)
  );
  LUT6 #(
    .INIT(64'hd8fad850d850d8fa)
  ) __6777__ (
    .I5(g3229),
    .I4(__1930__),
    .I3(__1928__),
    .I2(__133__),
    .I1(__1932__),
    .I0(__2095__),
    .O(__3094__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __6778__ (
    .I2(__858__),
    .I1(__2126__),
    .I0(__946__),
    .O(__3095__)
  );
  LUT6 #(
    .INIT(64'hf000b00000000000)
  ) __6779__ (
    .I5(__1596__),
    .I4(__1899__),
    .I3(__1595__),
    .I2(__603__),
    .I1(__1898__),
    .I0(__1921__),
    .O(__3096__)
  );
  LUT6 #(
    .INIT(64'hf5ffffff2222ffff)
  ) __6780__ (
    .I5(__1596__),
    .I4(__1595__),
    .I3(__2011__),
    .I2(__2009__),
    .I1(__1898__),
    .I0(__1887__),
    .O(__3097__)
  );
  LUT6 #(
    .INIT(64'h00000000bfffffff)
  ) __6781__ (
    .I5(__2014__),
    .I4(__1914__),
    .I3(__1910__),
    .I2(__1907__),
    .I1(__1903__),
    .I0(__2009__),
    .O(__3098__)
  );
  LUT6 #(
    .INIT(64'hfafffaccfafffaff)
  ) __6782__ (
    .I5(__603__),
    .I4(__1899__),
    .I3(__1596__),
    .I2(__1595__),
    .I1(__1887__),
    .I0(__3098__),
    .O(__3099__)
  );
  LUT6 #(
    .INIT(64'h00ff000040400000)
  ) __6783__ (
    .I5(__1597__),
    .I4(__1596__),
    .I3(__1595__),
    .I2(__3099__),
    .I1(__3097__),
    .I0(__3096__),
    .O(__3100__)
  );
  LUT3 #(
    .INIT(8'h10)
  ) __6784__ (
    .I2(__603__),
    .I1(__1899__),
    .I0(__1921__),
    .O(__3101__)
  );
  LUT5 #(
    .INIT(32'h0000004f)
  ) __6785__ (
    .I4(__1597__),
    .I3(__1596__),
    .I2(__3099__),
    .I1(__3101__),
    .I0(__3097__),
    .O(__3102__)
  );
  LUT5 #(
    .INIT(32'h00eef0f0)
  ) __6786__ (
    .I4(__663__),
    .I3(__2764__),
    .I2(__743__),
    .I1(__3102__),
    .I0(__3100__),
    .O(__3103__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6787__ (
    .I2(__589__),
    .I1(__2686__),
    .I0(__1268__),
    .O(__3104__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6788__ (
    .I2(__589__),
    .I1(__2272__),
    .I0(__687__),
    .O(__3105__)
  );
  LUT5 #(
    .INIT(32'h00eef0f0)
  ) __6789__ (
    .I4(__662__),
    .I3(__2764__),
    .I2(__1088__),
    .I1(__3102__),
    .I0(__3100__),
    .O(__3106__)
  );
  LUT5 #(
    .INIT(32'hf8070000)
  ) __6790__ (
    .I4(__2669__),
    .I3(__2056__),
    .I2(__2193__),
    .I1(__2668__),
    .I0(__2667__),
    .O(__3107__)
  );
  LUT5 #(
    .INIT(32'hf8070000)
  ) __6791__ (
    .I4(__2669__),
    .I3(__2056__),
    .I2(__2197__),
    .I1(__2668__),
    .I0(__2667__),
    .O(__3108__)
  );
  LUT6 #(
    .INIT(64'h003f00bb003fffbb)
  ) __6792__ (
    .I5(__3108__),
    .I4(__2183__),
    .I3(__2182__),
    .I2(__3107__),
    .I1(__2179__),
    .I0(__75__),
    .O(__3109__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __6793__ (
    .I3(__662__),
    .I2(__603__),
    .I1(__1450__),
    .I0(__826__),
    .O(__3110__)
  );
  LUT4 #(
    .INIT(16'haccc)
  ) __6794__ (
    .I3(__954__),
    .I2(__875__),
    .I1(__654__),
    .I0(__1951__),
    .O(__3111__)
  );
  LUT4 #(
    .INIT(16'h11f0)
  ) __6795__ (
    .I3(__662__),
    .I2(__787__),
    .I1(__2764__),
    .I0(__3000__),
    .O(__3112__)
  );
  LUT6 #(
    .INIT(64'h3fffff3faaaaaaaa)
  ) __6796__ (
    .I5(__2427__),
    .I4(g3229),
    .I3(__2287__),
    .I2(__2286__),
    .I1(__2285__),
    .I0(__599__),
    .O(__3113__)
  );
  LUT4 #(
    .INIT(16'h0baa)
  ) __6797__ (
    .I3(__858__),
    .I2(__1624__),
    .I1(__1949__),
    .I0(__121__),
    .O(__3114__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6798__ (
    .I2(__1479__),
    .I1(__1441__),
    .I0(__1466__),
    .O(__3115__)
  );
  LUT5 #(
    .INIT(32'h0c66cccc)
  ) __6799__ (
    .I4(__589__),
    .I3(__1598__),
    .I2(__603__),
    .I1(__657__),
    .I0(__658__),
    .O(__3116__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __6800__ (
    .I5(__858__),
    .I4(__242__),
    .I3(__370__),
    .I2(__229__),
    .I1(__278__),
    .I0(__366__),
    .O(__3117__)
  );
  LUT6 #(
    .INIT(64'haa3aaaaaaaaaaaaa)
  ) __6801__ (
    .I5(__858__),
    .I4(__93__),
    .I3(__748__),
    .I2(__73__),
    .I1(__1051__),
    .I0(__1406__),
    .O(__3118__)
  );
  LUT5 #(
    .INIT(32'haa20cf45)
  ) __6802__ (
    .I4(g3229),
    .I3(__2287__),
    .I2(__2286__),
    .I1(__2285__),
    .I0(__2369__),
    .O(__3119__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6803__ (
    .I2(__2288__),
    .I1(__3119__),
    .I0(__563__),
    .O(__3120__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __6804__ (
    .I1(__944__),
    .I0(__229__),
    .O(__3121__)
  );
  LUT6 #(
    .INIT(64'h132033005fa0ff00)
  ) __6805__ (
    .I5(__954__),
    .I4(__366__),
    .I3(__227__),
    .I2(__367__),
    .I1(__231__),
    .I0(__3121__),
    .O(__3122__)
  );
  LUT6 #(
    .INIT(64'h0100000100000000)
  ) __6806__ (
    .I5(__142__),
    .I4(__2056__),
    .I3(__2184__),
    .I2(__2178__),
    .I1(__140__),
    .I0(g1249),
    .O(__3123__)
  );
  LUT6 #(
    .INIT(64'hffffffff000f00bb)
  ) __6807__ (
    .I5(__2307__),
    .I4(__2183__),
    .I3(__2182__),
    .I2(__3123__),
    .I1(__2179__),
    .I0(__90__),
    .O(__3124__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6808__ (
    .I2(__2134__),
    .I1(__2962__),
    .I0(__983__),
    .O(__3125__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __6809__ (
    .I2(__589__),
    .I1(__2211__),
    .I0(__148__),
    .O(__3126__)
  );
  LUT6 #(
    .INIT(64'h0000baaaaaaaaaaa)
  ) __6810__ (
    .I5(__954__),
    .I4(__875__),
    .I3(__93__),
    .I2(__73__),
    .I1(__748__),
    .I0(__1332__),
    .O(__3127__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __6811__ (
    .I2(__589__),
    .I1(__1606__),
    .I0(__198__),
    .O(__3128__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __6812__ (
    .I5(__944__),
    .I4(__764__),
    .I3(__573__),
    .I2(__745__),
    .I1(__679__),
    .I0(__749__),
    .O(__3129__)
  );
  LUT6 #(
    .INIT(64'h4000000000000000)
  ) __6813__ (
    .I5(__944__),
    .I4(__227__),
    .I3(__366__),
    .I2(__367__),
    .I1(__225__),
    .I0(__229__),
    .O(__3130__)
  );
  LUT6 #(
    .INIT(64'h132033005fa0ff00)
  ) __6814__ (
    .I5(__954__),
    .I4(__224__),
    .I3(__220__),
    .I2(__222__),
    .I1(__231__),
    .I0(__3130__),
    .O(__3131__)
  );
  LUT6 #(
    .INIT(64'h0078787878787878)
  ) __6815__ (
    .I5(__589__),
    .I4(__1598__),
    .I3(__603__),
    .I2(__644__),
    .I1(__645__),
    .I0(__2978__),
    .O(__3132__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6816__ (
    .I2(__663__),
    .I1(__2167__),
    .I0(__666__),
    .O(__3133__)
  );
  LUT6 #(
    .INIT(64'hbfffffffa0000000)
  ) __6817__ (
    .I5(__537__),
    .I4(__662__),
    .I3(__603__),
    .I2(__2512__),
    .I1(__2278__),
    .I0(__2277__),
    .O(__3134__)
  );
  LUT5 #(
    .INIT(32'h12305af0)
  ) __6818__ (
    .I4(__954__),
    .I3(__224__),
    .I2(__222__),
    .I1(__231__),
    .I0(__3130__),
    .O(__3135__)
  );
  LUT4 #(
    .INIT(16'h0baa)
  ) __6819__ (
    .I3(__858__),
    .I2(__1624__),
    .I1(__1627__),
    .I0(__115__),
    .O(__3136__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __6820__ (
    .I5(__954__),
    .I4(__936__),
    .I3(__927__),
    .I2(__924__),
    .I1(__885__),
    .I0(__912__),
    .O(__3137__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __6821__ (
    .I3(__662__),
    .I2(__603__),
    .I1(__1442__),
    .I0(__838__),
    .O(__3138__)
  );
  LUT6 #(
    .INIT(64'h0f0f4444ff00ff00)
  ) __6822__ (
    .I5(__663__),
    .I4(__2516__),
    .I3(__1217__),
    .I2(__2515__),
    .I1(__1458__),
    .I0(__2514__),
    .O(__3139__)
  );
  LUT5 #(
    .INIT(32'h12121012)
  ) __6823__ (
    .I4(__1507__),
    .I3(__1508__),
    .I2(__1506__),
    .I1(g3234),
    .I0(__3066__),
    .O(__3140__)
  );
  LUT5 #(
    .INIT(32'h00eef0f0)
  ) __6824__ (
    .I4(__589__),
    .I3(__3007__),
    .I2(__583__),
    .I1(__3078__),
    .I0(__3076__),
    .O(__3141__)
  );
  LUT5 #(
    .INIT(32'h80000000)
  ) __6825__ (
    .I4(__1501__),
    .I3(__1499__),
    .I2(__1500__),
    .I1(__1498__),
    .I0(__215__),
    .O(__3142__)
  );
  LUT5 #(
    .INIT(32'h0000125a)
  ) __6826__ (
    .I4(g3234),
    .I3(__1623__),
    .I2(__1502__),
    .I1(__215__),
    .I0(__3142__),
    .O(__3143__)
  );
  LUT6 #(
    .INIT(64'hcc77f0f077ccf0f0)
  ) __6827__ (
    .I5(g3229),
    .I4(__2870__),
    .I3(__1602__),
    .I2(__1134__),
    .I1(__1600__),
    .I0(__1632__),
    .O(__3144__)
  );
  LUT4 #(
    .INIT(16'h0baa)
  ) __6828__ (
    .I3(__858__),
    .I2(__1624__),
    .I1(__2394__),
    .I0(__814__),
    .O(__3145__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __6829__ (
    .I5(__954__),
    .I4(__242__),
    .I3(__370__),
    .I2(__229__),
    .I1(__166__),
    .I0(__220__),
    .O(__3146__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __6830__ (
    .I5(__954__),
    .I4(__242__),
    .I3(__370__),
    .I2(__229__),
    .I1(__137__),
    .I0(__219__),
    .O(__3147__)
  );
  LUT4 #(
    .INIT(16'haccc)
  ) __6831__ (
    .I3(__663__),
    .I2(__603__),
    .I1(__226__),
    .I0(__1705__),
    .O(__3148__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6832__ (
    .I2(__944__),
    .I1(__867__),
    .I0(__1385__),
    .O(__3149__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __6833__ (
    .I1(__797__),
    .I0(__2197__),
    .O(__3150__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __6834__ (
    .I1(__788__),
    .I0(__2184__),
    .O(__3151__)
  );
  LUT6 #(
    .INIT(64'h1428000000000000)
  ) __6835__ (
    .I5(__3151__),
    .I4(__3150__),
    .I3(__1055__),
    .I2(__1047__),
    .I1(__2196__),
    .I0(__2191__),
    .O(__3152__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6836__ (
    .I1(__796__),
    .I0(__2185__),
    .O(__3153__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __6837__ (
    .I1(__796__),
    .I0(__2185__),
    .O(__3154__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __6838__ (
    .I1(__2180__),
    .I0(__737__),
    .O(__3155__)
  );
  LUT4 #(
    .INIT(16'h7770)
  ) __6839__ (
    .I3(__802__),
    .I2(__2193__),
    .I1(__2180__),
    .I0(__737__),
    .O(__3156__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __6840__ (
    .I1(__1051__),
    .I0(__2187__),
    .O(__3157__)
  );
  LUT6 #(
    .INIT(64'h0110000000000000)
  ) __6841__ (
    .I5(__3157__),
    .I4(__3156__),
    .I3(__747__),
    .I2(__2190__),
    .I1(__3155__),
    .I0(__3154__),
    .O(__3158__)
  );
  LUT6 #(
    .INIT(64'h0007070000000000)
  ) __6842__ (
    .I5(__3158__),
    .I4(__799__),
    .I3(__2192__),
    .I2(__3153__),
    .I1(__802__),
    .I0(__2193__),
    .O(__3159__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __6843__ (
    .I1(__944__),
    .I0(__855__),
    .O(__3160__)
  );
  LUT6 #(
    .INIT(64'h00008acf00000000)
  ) __6844__ (
    .I5(__2188__),
    .I4(__3160__),
    .I3(__858__),
    .I2(__954__),
    .I1(__654__),
    .I0(__349__),
    .O(__3161__)
  );
  LUT4 #(
    .INIT(16'h0080)
  ) __6845__ (
    .I3(__748__),
    .I2(__944__),
    .I1(__93__),
    .I0(__73__),
    .O(__3162__)
  );
  LUT5 #(
    .INIT(32'h3f00aaaa)
  ) __6846__ (
    .I4(__3162__),
    .I3(__3161__),
    .I2(__3159__),
    .I1(__3152__),
    .I0(__1336__),
    .O(__3163__)
  );
  LUT6 #(
    .INIT(64'h0f005555cccccccc)
  ) __6847__ (
    .I5(__663__),
    .I4(__603__),
    .I3(__1617__),
    .I2(__1614__),
    .I1(__1107__),
    .I0(__1613__),
    .O(__3164__)
  );
  LUT6 #(
    .INIT(64'hd8fad850d850d8fa)
  ) __6848__ (
    .I5(g3229),
    .I4(__2070__),
    .I3(__2068__),
    .I2(__632__),
    .I1(__2069__),
    .I0(__2774__),
    .O(__3165__)
  );
  LUT6 #(
    .INIT(64'h0000077007700000)
  ) __6849__ (
    .I5(__1678__),
    .I4(__606__),
    .I3(__1685__),
    .I2(__567__),
    .I1(__1687__),
    .I0(__512__),
    .O(__3166__)
  );
  LUT6 #(
    .INIT(64'h00000eee0eee0000)
  ) __6850__ (
    .I5(__1692__),
    .I4(__604__),
    .I3(__1691__),
    .I2(__568__),
    .I1(__1687__),
    .I0(__512__),
    .O(__3167__)
  );
  LUT5 #(
    .INIT(32'heee0eeee)
  ) __6851__ (
    .I4(__1682__),
    .I3(__1681__),
    .I2(__1680__),
    .I1(__1689__),
    .I0(__514__),
    .O(__3168__)
  );
  LUT6 #(
    .INIT(64'h0000077707770000)
  ) __6852__ (
    .I5(__1686__),
    .I4(__570__),
    .I3(__1689__),
    .I2(__514__),
    .I1(__1677__),
    .I0(__607__),
    .O(__3169__)
  );
  LUT6 #(
    .INIT(64'h0e00000000000000)
  ) __6853__ (
    .I5(__3169__),
    .I4(__3168__),
    .I3(__3167__),
    .I2(__1598__),
    .I1(__1691__),
    .I0(__568__),
    .O(__3170__)
  );
  LUT4 #(
    .INIT(16'h0ee0)
  ) __6854__ (
    .I3(__1690__),
    .I2(__605__),
    .I1(__1677__),
    .I0(__607__),
    .O(__3171__)
  );
  LUT6 #(
    .INIT(64'h155555559fffffff)
  ) __6855__ (
    .I5(__1697__),
    .I4(__3171__),
    .I3(__3170__),
    .I2(__3166__),
    .I1(__571__),
    .I0(__1679__),
    .O(__3172__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __6856__ (
    .I3(__663__),
    .I2(__603__),
    .I1(__1458__),
    .I0(__1308__),
    .O(__3173__)
  );
  LUT6 #(
    .INIT(64'haa3aaaaaaaaaaaaa)
  ) __6857__ (
    .I5(__944__),
    .I4(__93__),
    .I3(__748__),
    .I2(__73__),
    .I1(__802__),
    .I0(__1403__),
    .O(__3174__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __6858__ (
    .I1(__1524__),
    .I0(__1523__),
    .O(__3175__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __6859__ (
    .I1(__1526__),
    .I0(__1525__),
    .O(__3176__)
  );
  LUT6 #(
    .INIT(64'h6996966996696996)
  ) __6860__ (
    .I5(__1530__),
    .I4(__1529__),
    .I3(__1528__),
    .I2(__1527__),
    .I1(__3176__),
    .I0(__3175__),
    .O(__3177__)
  );
  LUT3 #(
    .INIT(8'hb4)
  ) __6861__ (
    .I2(__3177__),
    .I1(__1350__),
    .I0(g3231),
    .O(__3178__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6862__ (
    .I2(__589__),
    .I1(__2155__),
    .I0(__523__),
    .O(__3179__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __6863__ (
    .I2(__954__),
    .I1(__2975__),
    .I0(__805__),
    .O(__3180__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __6864__ (
    .I5(__944__),
    .I4(__242__),
    .I3(__370__),
    .I2(__229__),
    .I1(__209__),
    .I0(__367__),
    .O(__3181__)
  );
  LUT6 #(
    .INIT(64'h4eeeeeeeeeee4eee)
  ) __6865__ (
    .I5(g3229),
    .I4(__1930__),
    .I3(__1932__),
    .I2(__1928__),
    .I1(__124__),
    .I0(__2970__),
    .O(__3182__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __6866__ (
    .I3(__663__),
    .I2(__603__),
    .I1(__1455__),
    .I0(__1327__),
    .O(__3183__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6867__ (
    .I2(__662__),
    .I1(__2090__),
    .I0(__548__),
    .O(__3184__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __6868__ (
    .I3(__663__),
    .I2(__603__),
    .I1(__1413__),
    .I0(__210__),
    .O(__3185__)
  );
  LUT6 #(
    .INIT(64'h3fffff3faaaaaaaa)
  ) __6869__ (
    .I5(__1633__),
    .I4(g3229),
    .I3(__1602__),
    .I2(__1601__),
    .I1(__1600__),
    .I0(__1130__),
    .O(__3186__)
  );
  LUT6 #(
    .INIT(64'h3fffff3faaaaaaaa)
  ) __6870__ (
    .I5(__2062__),
    .I4(g3229),
    .I3(__2065__),
    .I2(__2063__),
    .I1(__2064__),
    .I0(__1196__),
    .O(__3187__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6871__ (
    .I2(__1479__),
    .I1(__1468__),
    .I0(__1407__),
    .O(__3188__)
  );
  LUT6 #(
    .INIT(64'haa3aaaaaaaaaaaaa)
  ) __6872__ (
    .I5(__954__),
    .I4(__93__),
    .I3(__748__),
    .I2(__73__),
    .I1(__796__),
    .I0(__786__),
    .O(__3189__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6873__ (
    .I2(__663__),
    .I1(__2355__),
    .I0(__707__),
    .O(__3190__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __6874__ (
    .I5(__944__),
    .I4(__93__),
    .I3(__73__),
    .I2(__748__),
    .I1(__1392__),
    .I0(__737__),
    .O(__3191__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6875__ (
    .I2(__944__),
    .I1(__2397__),
    .I0(__807__),
    .O(__3192__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __6876__ (
    .I3(__662__),
    .I2(__603__),
    .I1(__1419__),
    .I0(__1323__),
    .O(__3193__)
  );
  LUT6 #(
    .INIT(64'hfa000f0fcccccccc)
  ) __6877__ (
    .I5(__663__),
    .I4(__603__),
    .I3(__2585__),
    .I2(__2508__),
    .I1(__1195__),
    .I0(__2509__),
    .O(__3194__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __6878__ (
    .I3(__589__),
    .I2(__603__),
    .I1(__1428__),
    .I0(__1302__),
    .O(__3195__)
  );
  LUT6 #(
    .INIT(64'h0100000100000000)
  ) __6879__ (
    .I5(__300__),
    .I4(__1800__),
    .I3(__1786__),
    .I2(__297__),
    .I1(g2637),
    .I0(__1784__),
    .O(__3196__)
  );
  LUT6 #(
    .INIT(64'hffffffff000f00bb)
  ) __6880__ (
    .I5(__3016__),
    .I4(__2646__),
    .I3(__2645__),
    .I2(__3196__),
    .I1(__1802__),
    .I0(__238__),
    .O(__3197__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __6881__ (
    .I1(__3089__),
    .I0(__1478__),
    .O(__3198__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6882__ (
    .I2(__589__),
    .I1(__2886__),
    .I0(__1245__),
    .O(__3199__)
  );
  LUT4 #(
    .INIT(16'haccc)
  ) __6883__ (
    .I3(__954__),
    .I2(__752__),
    .I1(__677__),
    .I0(__1646__),
    .O(__3200__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __6884__ (
    .I1(__2627__),
    .I0(__929__),
    .O(__3201__)
  );
  LUT6 #(
    .INIT(64'h00000f0f00ff4444)
  ) __6885__ (
    .I5(__1037__),
    .I4(__1036__),
    .I3(__2901__),
    .I2(__2905__),
    .I1(__936__),
    .I0(__3201__),
    .O(__3202__)
  );
  LUT4 #(
    .INIT(16'haccc)
  ) __6886__ (
    .I3(__954__),
    .I2(__231__),
    .I1(__292__),
    .I0(__1982__),
    .O(__3203__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __6887__ (
    .I5(__954__),
    .I4(__242__),
    .I3(__370__),
    .I2(__229__),
    .I1(__212__),
    .I0(__367__),
    .O(__3204__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6888__ (
    .I2(__3049__),
    .I1(__1980__),
    .I0(__294__),
    .O(__3205__)
  );
  LUT6 #(
    .INIT(64'haa3aaaaaaaaaaaaa)
  ) __6889__ (
    .I5(__954__),
    .I4(__93__),
    .I3(__748__),
    .I2(__73__),
    .I1(__1055__),
    .I0(__729__),
    .O(__3206__)
  );
  LUT5 #(
    .INIT(32'h0030aaaa)
  ) __6890__ (
    .I4(__589__),
    .I3(__1682__),
    .I2(__1681__),
    .I1(__1680__),
    .I0(__391__),
    .O(__3207__)
  );
  LUT5 #(
    .INIT(32'hcd000000)
  ) __6891__ (
    .I4(__663__),
    .I3(__603__),
    .I2(__1710__),
    .I1(__2263__),
    .I0(__2262__),
    .O(__3208__)
  );
  LUT6 #(
    .INIT(64'hffff0707ff00ff00)
  ) __6892__ (
    .I5(__3208__),
    .I4(__1682__),
    .I3(__118__),
    .I2(__2257__),
    .I1(__1680__),
    .I0(__2256__),
    .O(__3209__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6893__ (
    .I2(__662__),
    .I1(__2608__),
    .I0(__1272__),
    .O(__3210__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6894__ (
    .I2(__589__),
    .I1(__1733__),
    .I0(__614__),
    .O(__3211__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __6895__ (
    .I2(__662__),
    .I1(__2279__),
    .I0(__184__),
    .O(__3212__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __6896__ (
    .I5(__944__),
    .I4(__149__),
    .I3(__858__),
    .I2(__148__),
    .I1(__954__),
    .I0(__150__),
    .O(__3213__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __6897__ (
    .I3(__662__),
    .I2(__603__),
    .I1(__1408__),
    .I0(__427__),
    .O(__3214__)
  );
  LUT6 #(
    .INIT(64'h4545ff000505ff00)
  ) __6898__ (
    .I5(__858__),
    .I4(__944__),
    .I3(__113__),
    .I2(__1627__),
    .I1(__115__),
    .I0(__1624__),
    .O(__3215__)
  );
  LUT6 #(
    .INIT(64'haa3aaaaaaaaaaaaa)
  ) __6899__ (
    .I5(__858__),
    .I4(__93__),
    .I3(__748__),
    .I2(__73__),
    .I1(__799__),
    .I0(__1402__),
    .O(__3216__)
  );
  LUT6 #(
    .INIT(64'hcf300000aaaaaaaa)
  ) __6900__ (
    .I5(__589__),
    .I4(__1999__),
    .I3(__1759__),
    .I2(__1998__),
    .I1(__1992__),
    .I0(__414__),
    .O(__3217__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __6901__ (
    .I3(__589__),
    .I2(__603__),
    .I1(__1456__),
    .I0(__1312__),
    .O(__3218__)
  );
  LUT6 #(
    .INIT(64'h0000077007700000)
  ) __6902__ (
    .I5(__1539__),
    .I4(__1235__),
    .I3(__1536__),
    .I2(__1222__),
    .I1(__1540__),
    .I0(__1220__),
    .O(__3219__)
  );
  LUT6 #(
    .INIT(64'h00000eee0eee0000)
  ) __6903__ (
    .I5(__1550__),
    .I4(__1223__),
    .I3(__1549__),
    .I2(__1228__),
    .I1(__1540__),
    .I0(__1220__),
    .O(__3220__)
  );
  LUT5 #(
    .INIT(32'heee0eeee)
  ) __6904__ (
    .I4(__1543__),
    .I3(__1544__),
    .I2(__1542__),
    .I1(__1547__),
    .I0(__1232__),
    .O(__3221__)
  );
  LUT6 #(
    .INIT(64'h0000077707770000)
  ) __6905__ (
    .I5(__1537__),
    .I4(__1234__),
    .I3(__1547__),
    .I2(__1232__),
    .I1(__1546__),
    .I0(__1237__),
    .O(__3222__)
  );
  LUT6 #(
    .INIT(64'h0e00000000000000)
  ) __6906__ (
    .I5(__3222__),
    .I4(__3221__),
    .I3(__3220__),
    .I2(__1598__),
    .I1(__1549__),
    .I0(__1228__),
    .O(__3223__)
  );
  LUT4 #(
    .INIT(16'h0ee0)
  ) __6907__ (
    .I3(__1548__),
    .I2(__1224__),
    .I1(__1546__),
    .I0(__1237__),
    .O(__3224__)
  );
  LUT6 #(
    .INIT(64'h155555559fffffff)
  ) __6908__ (
    .I5(__1555__),
    .I4(__3224__),
    .I3(__3223__),
    .I2(__3219__),
    .I1(__1236__),
    .I0(__1538__),
    .O(__3225__)
  );
  LUT4 #(
    .INIT(16'h125a)
  ) __6909__ (
    .I3(__954__),
    .I2(__737__),
    .I1(__875__),
    .I0(__1668__),
    .O(__3226__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __6910__ (
    .I3(__589__),
    .I2(__603__),
    .I1(__1407__),
    .I0(__432__),
    .O(__3227__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __6911__ (
    .I3(__663__),
    .I2(__603__),
    .I1(__1412__),
    .I0(__638__),
    .O(__3228__)
  );
  LUT4 #(
    .INIT(16'h0008)
  ) __6912__ (
    .I3(__1430__),
    .I2(__1428__),
    .I1(__1426__),
    .I0(__1432__),
    .O(__3229__)
  );
  LUT5 #(
    .INIT(32'hb8f0f0f0)
  ) __6913__ (
    .I4(__662__),
    .I3(__1598__),
    .I2(__1287__),
    .I1(__1635__),
    .I0(__3229__),
    .O(__3230__)
  );
  LUT5 #(
    .INIT(32'hf8070000)
  ) __6914__ (
    .I4(__2344__),
    .I3(__1649__),
    .I2(__1823__),
    .I1(__2343__),
    .I0(__2342__),
    .O(__3231__)
  );
  LUT5 #(
    .INIT(32'hf8070000)
  ) __6915__ (
    .I4(__2344__),
    .I3(__1649__),
    .I2(__1818__),
    .I1(__2343__),
    .I0(__2342__),
    .O(__3232__)
  );
  LUT5 #(
    .INIT(32'h000000e0)
  ) __6916__ (
    .I4(__968__),
    .I3(__103__),
    .I2(__2346__),
    .I1(__764__),
    .I0(__969__),
    .O(__3233__)
  );
  LUT6 #(
    .INIT(64'h000000330f0f00aa)
  ) __6917__ (
    .I5(__968__),
    .I4(__969__),
    .I3(__3233__),
    .I2(__3232__),
    .I1(__3231__),
    .I0(__764__),
    .O(__3234__)
  );
  LUT2 #(
    .INIT(4'he)
  ) __6918__ (
    .I1(g51),
    .I0(__1495__),
    .O(__3235__)
  );
  LUT6 #(
    .INIT(64'h000a000c00000000)
  ) __6919__ (
    .I5(__93__),
    .I4(g3229),
    .I3(__266__),
    .I2(__269__),
    .I1(__72__),
    .I0(__73__),
    .O(__3236__)
  );
  LUT5 #(
    .INIT(32'h70077777)
  ) __6920__ (
    .I4(__269__),
    .I3(__2670__),
    .I2(__3108__),
    .I1(__2179__),
    .I0(__3236__),
    .O(__3237__)
  );
  LUT4 #(
    .INIT(16'h9669)
  ) __6921__ (
    .I3(__2711__),
    .I2(__2767__),
    .I1(__2666__),
    .I0(__3107__),
    .O(__3238__)
  );
  LUT5 #(
    .INIT(32'h28828228)
  ) __6922__ (
    .I4(__2056__),
    .I3(__2180__),
    .I2(__2191__),
    .I1(__1951__),
    .I0(__2669__),
    .O(__3239__)
  );
  LUT6 #(
    .INIT(64'h0100000100000000)
  ) __6923__ (
    .I5(__142__),
    .I4(__2185__),
    .I3(__1951__),
    .I2(__2178__),
    .I1(__140__),
    .I0(g1249),
    .O(__3240__)
  );
  LUT6 #(
    .INIT(64'hd77d7dd755555555)
  ) __6924__ (
    .I5(__266__),
    .I4(__3240__),
    .I3(__3123__),
    .I2(__3239__),
    .I1(__3238__),
    .I0(__3237__),
    .O(__3241__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __6925__ (
    .I3(__662__),
    .I2(__2282__),
    .I1(__1419__),
    .I0(__1284__),
    .O(__3242__)
  );
  LUT6 #(
    .INIT(64'h0000bfff00000000)
  ) __6926__ (
    .I5(g3233),
    .I4(g3230),
    .I3(__1352__),
    .I2(__2939__),
    .I1(__2942__),
    .I0(__1345__),
    .O(__3243__)
  );
  LUT5 #(
    .INIT(32'hcd000000)
  ) __6927__ (
    .I4(__663__),
    .I3(__603__),
    .I2(__1757__),
    .I1(__2314__),
    .I0(__1997__),
    .O(__3244__)
  );
  LUT6 #(
    .INIT(64'hffff0707ff00ff00)
  ) __6928__ (
    .I5(__3244__),
    .I4(__1761__),
    .I3(__411__),
    .I2(__2313__),
    .I1(__1759__),
    .I0(__2312__),
    .O(__3245__)
  );
  LUT5 #(
    .INIT(32'ha000cccc)
  ) __6929__ (
    .I4(__663__),
    .I3(__1543__),
    .I2(__1544__),
    .I1(__998__),
    .I0(__1542__),
    .O(__3246__)
  );
  LUT3 #(
    .INIT(8'hb4)
  ) __6930__ (
    .I2(__2335__),
    .I1(__1350__),
    .I0(g3231),
    .O(__3247__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __6931__ (
    .I3(__662__),
    .I2(__603__),
    .I1(__1417__),
    .I0(__1341__),
    .O(__3248__)
  );
  LUT5 #(
    .INIT(32'h00f4f0f0)
  ) __6932__ (
    .I4(__663__),
    .I3(__2405__),
    .I2(__1177__),
    .I1(__603__),
    .I0(__2404__),
    .O(__3249__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6933__ (
    .I2(__2173__),
    .I1(__2676__),
    .I0(__139__),
    .O(__3250__)
  );
  LUT6 #(
    .INIT(64'h4545ff000505ff00)
  ) __6934__ (
    .I5(__858__),
    .I4(__944__),
    .I3(__810__),
    .I2(__1665__),
    .I1(__812__),
    .I0(__1624__),
    .O(__3251__)
  );
  LUT4 #(
    .INIT(16'haccc)
  ) __6935__ (
    .I3(__954__),
    .I2(__752__),
    .I1(__674__),
    .I0(__1649__),
    .O(__3252__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6936__ (
    .I2(__663__),
    .I1(__2364__),
    .I0(__1165__),
    .O(__3253__)
  );
  LUT4 #(
    .INIT(16'h25aa)
  ) __6937__ (
    .I3(__589__),
    .I2(__1598__),
    .I1(__603__),
    .I0(__1180__),
    .O(__3254__)
  );
  LUT4 #(
    .INIT(16'haccc)
  ) __6938__ (
    .I3(__662__),
    .I2(__603__),
    .I1(__593__),
    .I0(__1705__),
    .O(__3255__)
  );
  LUT6 #(
    .INIT(64'h0078787878787878)
  ) __6939__ (
    .I5(__589__),
    .I4(__1598__),
    .I3(__603__),
    .I2(__605__),
    .I1(__568__),
    .I0(__2149__),
    .O(__3256__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6940__ (
    .I2(__944__),
    .I1(__1036__),
    .I0(__925__),
    .O(__3257__)
  );
  LUT5 #(
    .INIT(32'ha000cccc)
  ) __6941__ (
    .I4(__944__),
    .I3(__1036__),
    .I2(__1806__),
    .I1(__940__),
    .I0(__1805__),
    .O(__3258__)
  );
  LUT6 #(
    .INIT(64'h0f005555cccccccc)
  ) __6942__ (
    .I5(__663__),
    .I4(__603__),
    .I3(__2089__),
    .I2(__2084__),
    .I1(__551__),
    .I0(__2085__),
    .O(__3259__)
  );
  LUT4 #(
    .INIT(16'h11f0)
  ) __6943__ (
    .I3(__662__),
    .I2(__1169__),
    .I1(__2621__),
    .I0(__2620__),
    .O(__3260__)
  );
  LUT6 #(
    .INIT(64'hbfffffffa0000000)
  ) __6944__ (
    .I5(__1120__),
    .I4(__589__),
    .I3(__603__),
    .I2(__2417__),
    .I1(__2247__),
    .I0(__2248__),
    .O(__3261__)
  );
  LUT5 #(
    .INIT(32'h00000080)
  ) __6945__ (
    .I4(__1351__),
    .I3(__1350__),
    .I2(__1349__),
    .I1(__1352__),
    .I0(__2944__),
    .O(__3262__)
  );
  LUT6 #(
    .INIT(64'hf53fffffffffffff)
  ) __6946__ (
    .I5(__2944__),
    .I4(__2952__),
    .I3(__1351__),
    .I2(__1352__),
    .I1(__1385__),
    .I0(__1389__),
    .O(__3263__)
  );
  LUT6 #(
    .INIT(64'h0000000000004ccc)
  ) __6947__ (
    .I5(__2769__),
    .I4(__2947__),
    .I3(__2944__),
    .I2(__1397__),
    .I1(__3263__),
    .I0(__2938__),
    .O(__3264__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __6948__ (
    .I1(__1481__),
    .I0(__1482__),
    .O(__3265__)
  );
  LUT3 #(
    .INIT(8'h01)
  ) __6949__ (
    .I2(__1351__),
    .I1(__1350__),
    .I0(__1349__),
    .O(__3266__)
  );
  LUT3 #(
    .INIT(8'h08)
  ) __6950__ (
    .I2(__1349__),
    .I1(__1351__),
    .I0(__1350__),
    .O(__3267__)
  );
  LUT5 #(
    .INIT(32'h53ffffff)
  ) __6951__ (
    .I4(__2942__),
    .I3(__2944__),
    .I2(__1352__),
    .I1(__1395__),
    .I0(__1383__),
    .O(__3268__)
  );
  LUT6 #(
    .INIT(64'h0f00bb00ff00ff00)
  ) __6952__ (
    .I5(__2939__),
    .I4(__1352__),
    .I3(__3268__),
    .I2(__3267__),
    .I1(__3266__),
    .I0(__3265__),
    .O(__3269__)
  );
  LUT5 #(
    .INIT(32'h00000080)
  ) __6953__ (
    .I4(__1351__),
    .I3(__1350__),
    .I2(__1349__),
    .I1(__2940__),
    .I0(__1396__),
    .O(__3270__)
  );
  LUT6 #(
    .INIT(64'h05030f0f0f0f0f0f)
  ) __6954__ (
    .I5(__2944__),
    .I4(__2950__),
    .I3(__1352__),
    .I2(__3270__),
    .I1(__1394__),
    .I0(__1382__),
    .O(__3271__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __6955__ (
    .I2(__1351__),
    .I1(__1350__),
    .I0(__1349__),
    .O(__3272__)
  );
  LUT5 #(
    .INIT(32'h00008000)
  ) __6956__ (
    .I4(__1350__),
    .I3(__1351__),
    .I2(__1349__),
    .I1(__1388__),
    .I0(__2940__),
    .O(__3273__)
  );
  LUT6 #(
    .INIT(64'h000000000777ffff)
  ) __6957__ (
    .I5(__3273__),
    .I4(__2940__),
    .I3(__1386__),
    .I2(__3272__),
    .I1(__3267__),
    .I0(__1387__),
    .O(__3274__)
  );
  LUT6 #(
    .INIT(64'h8fffffffffffffff)
  ) __6958__ (
    .I5(__3274__),
    .I4(__3271__),
    .I3(__3269__),
    .I2(__3264__),
    .I1(__3262__),
    .I0(__1384__),
    .O(__3275__)
  );
  LUT6 #(
    .INIT(64'h0000baaaaaaaaaaa)
  ) __6959__ (
    .I5(__944__),
    .I4(__925__),
    .I3(__936__),
    .I2(__927__),
    .I1(__924__),
    .I0(__851__),
    .O(__3276__)
  );
  LUT6 #(
    .INIT(64'h0000baaaaaaaaaaa)
  ) __6960__ (
    .I5(__858__),
    .I4(__925__),
    .I3(__936__),
    .I2(__927__),
    .I1(__924__),
    .I0(__854__),
    .O(__3277__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __6961__ (
    .I3(__662__),
    .I2(__2282__),
    .I1(__1436__),
    .I0(__776__),
    .O(__3278__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __6962__ (
    .I3(__589__),
    .I2(__603__),
    .I1(__1410__),
    .I0(__665__),
    .O(__3279__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6963__ (
    .I2(__1650__),
    .I1(__3002__),
    .I0(__577__),
    .O(__3280__)
  );
  LUT6 #(
    .INIT(64'h4545ff000505ff00)
  ) __6964__ (
    .I5(__858__),
    .I4(__954__),
    .I3(__813__),
    .I2(__2394__),
    .I1(__814__),
    .I0(__1624__),
    .O(__3281__)
  );
  LUT4 #(
    .INIT(16'haccc)
  ) __6965__ (
    .I3(__858__),
    .I2(__231__),
    .I1(__152__),
    .I0(__1800__),
    .O(__3282__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6966__ (
    .I2(__1479__),
    .I1(__1470__),
    .I0(__1460__),
    .O(__3283__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __6967__ (
    .I2(__944__),
    .I1(__2975__),
    .I0(__804__),
    .O(__3284__)
  );
  LUT6 #(
    .INIT(64'hf000f0ccaaaaaaaa)
  ) __6968__ (
    .I5(__954__),
    .I4(__858__),
    .I3(__988__),
    .I2(__991__),
    .I1(__990__),
    .I0(__1380__),
    .O(__3285__)
  );
  LUT4 #(
    .INIT(16'haccc)
  ) __6969__ (
    .I3(__662__),
    .I2(__603__),
    .I1(__822__),
    .I0(__1742__),
    .O(__3286__)
  );
  LUT6 #(
    .INIT(64'h0f005555cccccccc)
  ) __6970__ (
    .I5(__662__),
    .I4(__603__),
    .I3(__2140__),
    .I2(__2137__),
    .I1(__527__),
    .I0(__2136__),
    .O(__3287__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6971__ (
    .I2(__944__),
    .I1(__1647__),
    .I0(__924__),
    .O(__3288__)
  );
  LUT6 #(
    .INIT(64'hffffffff000f00bb)
  ) __6972__ (
    .I5(__2200__),
    .I4(__2183__),
    .I3(__2182__),
    .I2(__3240__),
    .I1(__2179__),
    .I0(__85__),
    .O(__3289__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6973__ (
    .I2(__2568__),
    .I1(__2881__),
    .I0(__1215__),
    .O(__3290__)
  );
  LUT5 #(
    .INIT(32'ha000cccc)
  ) __6974__ (
    .I4(__663__),
    .I3(__1761__),
    .I2(__1760__),
    .I1(__181__),
    .I0(__1759__),
    .O(__3291__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __6975__ (
    .I5(__764__),
    .I4(__573__),
    .I3(__954__),
    .I2(__745__),
    .I1(__690__),
    .I0(__772__),
    .O(__3292__)
  );
  LUT5 #(
    .INIT(32'h007f0080)
  ) __6976__ (
    .I4(__1161__),
    .I3(__2151__),
    .I2(__730__),
    .I1(__1164__),
    .I0(__2924__),
    .O(__3293__)
  );
  LUT5 #(
    .INIT(32'hccaa0f0f)
  ) __6977__ (
    .I4(__501__),
    .I3(__662__),
    .I2(__499__),
    .I1(__2914__),
    .I0(__500__),
    .O(__3294__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __6978__ (
    .I3(__663__),
    .I2(__2282__),
    .I1(__1617__),
    .I0(__1262__),
    .O(__3295__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __6979__ (
    .I5(__858__),
    .I4(__93__),
    .I3(__73__),
    .I2(__748__),
    .I1(__798__),
    .I0(__797__),
    .O(__3296__)
  );
  LUT6 #(
    .INIT(64'h132033005fa0ff00)
  ) __6980__ (
    .I5(__954__),
    .I4(__770__),
    .I3(__749__),
    .I2(__741__),
    .I1(__752__),
    .I0(__1986__),
    .O(__3297__)
  );
  LUT5 #(
    .INIT(32'hcd000000)
  ) __6981__ (
    .I4(__662__),
    .I3(__603__),
    .I2(__1757__),
    .I1(__2314__),
    .I0(__1997__),
    .O(__3298__)
  );
  LUT6 #(
    .INIT(64'hffff0707ff00ff00)
  ) __6982__ (
    .I5(__3298__),
    .I4(__1761__),
    .I3(__408__),
    .I2(__2313__),
    .I1(__1759__),
    .I0(__2312__),
    .O(__3299__)
  );
  LUT6 #(
    .INIT(64'haaaacaaaaaaaaaaa)
  ) __6983__ (
    .I5(__954__),
    .I4(__229__),
    .I3(__242__),
    .I2(__370__),
    .I1(__2425__),
    .I0(__248__),
    .O(__3300__)
  );
  LUT6 #(
    .INIT(64'h00007fff00008000)
  ) __6984__ (
    .I5(__1222__),
    .I4(__2151__),
    .I3(__1228__),
    .I2(__2713__),
    .I1(__1224__),
    .I0(__1223__),
    .O(__3301__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __6985__ (
    .I5(__944__),
    .I4(__242__),
    .I3(__370__),
    .I2(__229__),
    .I1(__180__),
    .I0(__224__),
    .O(__3302__)
  );
  LUT3 #(
    .INIT(8'h06)
  ) __6986__ (
    .I2(g3234),
    .I1(__1498__),
    .I0(__215__),
    .O(__3303__)
  );
  LUT4 #(
    .INIT(16'h0008)
  ) __6987__ (
    .I3(__1458__),
    .I2(__1459__),
    .I1(__1460__),
    .I0(__1457__),
    .O(__3304__)
  );
  LUT5 #(
    .INIT(32'hb8f0f0f0)
  ) __6988__ (
    .I4(__662__),
    .I3(__1598__),
    .I2(__1264__),
    .I1(__1635__),
    .I0(__3304__),
    .O(__3305__)
  );
  LUT5 #(
    .INIT(32'hf0f06633)
  ) __6989__ (
    .I4(__1479__),
    .I3(__1349__),
    .I2(__1416__),
    .I1(__3089__),
    .I0(g3231),
    .O(__3306__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6990__ (
    .I2(__1479__),
    .I1(__1464__),
    .I0(__1411__),
    .O(__3307__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6991__ (
    .I2(__663__),
    .I1(__2886__),
    .I0(__1247__),
    .O(__3308__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __6992__ (
    .I5(__764__),
    .I4(__573__),
    .I3(__954__),
    .I2(__745__),
    .I1(__746__),
    .I0(__760__),
    .O(__3309__)
  );
  LUT4 #(
    .INIT(16'he7ee)
  ) __6993__ (
    .I3(__2089__),
    .I2(__2084__),
    .I1(__2085__),
    .I0(__1957__),
    .O(__3310__)
  );
  LUT6 #(
    .INIT(64'h108000c000000000)
  ) __6994__ (
    .I5(__603__),
    .I4(__2089__),
    .I3(__1957__),
    .I2(__2086__),
    .I1(__2085__),
    .I0(__2084__),
    .O(__3311__)
  );
  LUT5 #(
    .INIT(32'h00f4f0f0)
  ) __6995__ (
    .I4(__663__),
    .I3(__3311__),
    .I2(__546__),
    .I1(__603__),
    .I0(__3310__),
    .O(__3312__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __6996__ (
    .I2(__663__),
    .I1(__2279__),
    .I0(__185__),
    .O(__3313__)
  );
  LUT4 #(
    .INIT(16'h11f0)
  ) __6997__ (
    .I3(__663__),
    .I2(__1170__),
    .I1(__2621__),
    .I0(__2620__),
    .O(__3314__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6998__ (
    .I2(__663__),
    .I1(__2765__),
    .I0(__1084__),
    .O(__3315__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __6999__ (
    .I2(__589__),
    .I1(__2249__),
    .I0(__429__),
    .O(__3316__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __7000__ (
    .I3(__589__),
    .I2(__603__),
    .I1(__1424__),
    .I0(__1316__),
    .O(__3317__)
  );
  LUT5 #(
    .INIT(32'h0c66cccc)
  ) __7001__ (
    .I4(__589__),
    .I3(__1598__),
    .I2(__603__),
    .I1(__571__),
    .I0(__607__),
    .O(__3318__)
  );
  LUT2 #(
    .INIT(4'h7)
  ) __7002__ (
    .I1(__1597__),
    .I0(__1595__),
    .O(__3319__)
  );
  LUT6 #(
    .INIT(64'h5555fccf55555555)
  ) __7003__ (
    .I5(__2015__),
    .I4(__2012__),
    .I3(__1877__),
    .I2(__3319__),
    .I1(__2008__),
    .I0(__1453__),
    .O(__3320__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __7004__ (
    .I2(__589__),
    .I1(__3320__),
    .I0(__1243__),
    .O(__3321__)
  );
  LUT6 #(
    .INIT(64'h0f0f4444ff00ff00)
  ) __7005__ (
    .I5(__662__),
    .I4(__2867__),
    .I3(__450__),
    .I2(__2866__),
    .I1(__1412__),
    .I0(__2865__),
    .O(__3322__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7006__ (
    .I2(__663__),
    .I1(__1865__),
    .I0(__725__),
    .O(__3323__)
  );
  LUT6 #(
    .INIT(64'h1113020013130000)
  ) __7007__ (
    .I5(__1499__),
    .I4(__1500__),
    .I3(__1498__),
    .I2(__1623__),
    .I1(g3234),
    .I0(__215__),
    .O(__3324__)
  );
  LUT4 #(
    .INIT(16'haccc)
  ) __7008__ (
    .I3(__662__),
    .I2(__603__),
    .I1(__1293__),
    .I0(__1565__),
    .O(__3325__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __7009__ (
    .I2(__663__),
    .I1(__2357__),
    .I0(__710__),
    .O(__3326__)
  );
  LUT5 #(
    .INIT(32'ha000cccc)
  ) __7010__ (
    .I4(__858__),
    .I3(__1951__),
    .I2(__2094__),
    .I1(__106__),
    .I0(__266__),
    .O(__3327__)
  );
  LUT6 #(
    .INIT(64'h0000000000008000)
  ) __7011__ (
    .I5(__1351__),
    .I4(__1350__),
    .I3(__1349__),
    .I2(__1352__),
    .I1(__2944__),
    .I0(__1359__),
    .O(__3328__)
  );
  LUT6 #(
    .INIT(64'h05030f0f0f0f0f0f)
  ) __7012__ (
    .I5(__1352__),
    .I4(__2939__),
    .I3(__1351__),
    .I2(__2769__),
    .I1(__2958__),
    .I0(__2952__),
    .O(__3329__)
  );
  LUT6 #(
    .INIT(64'hf53fffffffffffff)
  ) __7013__ (
    .I5(__2944__),
    .I4(__2952__),
    .I3(__1351__),
    .I2(__1352__),
    .I1(__1360__),
    .I0(__1365__),
    .O(__3330__)
  );
  LUT6 #(
    .INIT(64'h0fff7777ffffffff)
  ) __7014__ (
    .I5(__2940__),
    .I4(__1351__),
    .I3(__2954__),
    .I2(__1361__),
    .I1(__2955__),
    .I0(__1368__),
    .O(__3331__)
  );
  LUT6 #(
    .INIT(64'h0777ffffffffffff)
  ) __7015__ (
    .I5(__1351__),
    .I4(__2940__),
    .I3(__1362__),
    .I2(__2958__),
    .I1(__2955__),
    .I0(__1363__),
    .O(__3332__)
  );
  LUT6 #(
    .INIT(64'h0777ffffffffffff)
  ) __7016__ (
    .I5(__1352__),
    .I4(__2944__),
    .I3(__2942__),
    .I2(__1358__),
    .I1(__1357__),
    .I0(__2950__),
    .O(__3333__)
  );
  LUT6 #(
    .INIT(64'h0000000000000008)
  ) __7017__ (
    .I5(__1351__),
    .I4(__1350__),
    .I3(__1349__),
    .I2(__1352__),
    .I1(__2944__),
    .I0(__1369__),
    .O(__3334__)
  );
  LUT5 #(
    .INIT(32'h00008000)
  ) __7018__ (
    .I4(__1351__),
    .I3(__1350__),
    .I2(__1349__),
    .I1(__1366__),
    .I0(__2940__),
    .O(__3335__)
  );
  LUT5 #(
    .INIT(32'h00000080)
  ) __7019__ (
    .I4(__3335__),
    .I3(__3334__),
    .I2(__3333__),
    .I1(__3332__),
    .I0(__3331__),
    .O(__3336__)
  );
  LUT6 #(
    .INIT(64'hf8ffffffffffffff)
  ) __7020__ (
    .I5(__3336__),
    .I4(__3330__),
    .I3(__3329__),
    .I2(__3328__),
    .I1(__2941__),
    .I0(__1367__),
    .O(__3337__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7021__ (
    .I2(__589__),
    .I1(__2690__),
    .I0(__1238__),
    .O(__3338__)
  );
  LUT6 #(
    .INIT(64'hd8fad850d850d8fa)
  ) __7022__ (
    .I5(g3229),
    .I4(__1979__),
    .I3(__1978__),
    .I2(__290__),
    .I1(__1977__),
    .I0(__3049__),
    .O(__3339__)
  );
  LUT6 #(
    .INIT(64'hbfffffffa0000000)
  ) __7023__ (
    .I5(__596__),
    .I4(__662__),
    .I3(__603__),
    .I2(__2462__),
    .I1(__2210__),
    .I0(__2209__),
    .O(__3340__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __7024__ (
    .I1(__1469__),
    .I0(__2830__),
    .O(__3341__)
  );
  LUT6 #(
    .INIT(64'h1320330031003300)
  ) __7025__ (
    .I5(__1484__),
    .I4(__1486__),
    .I3(__1483__),
    .I2(__1485__),
    .I1(__1497__),
    .I0(__1611__),
    .O(__3342__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7026__ (
    .I2(__944__),
    .I1(__1037__),
    .I0(__1036__),
    .O(__3343__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __7027__ (
    .I2(__589__),
    .I1(__2019__),
    .I0(__738__),
    .O(__3344__)
  );
  LUT6 #(
    .INIT(64'h0000baaaaaaaaaaa)
  ) __7028__ (
    .I5(__858__),
    .I4(__752__),
    .I3(__764__),
    .I2(__573__),
    .I1(__745__),
    .I0(__669__),
    .O(__3345__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __7029__ (
    .I1(__1531__),
    .I0(__3177__),
    .O(__3346__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7030__ (
    .I2(__954__),
    .I1(__2120__),
    .I0(__275__),
    .O(__3347__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __7031__ (
    .I2(__662__),
    .I1(__3012__),
    .I0(__1203__),
    .O(__3348__)
  );
  LUT4 #(
    .INIT(16'h0080)
  ) __7032__ (
    .I3(__924__),
    .I2(__858__),
    .I1(__936__),
    .I0(__927__),
    .O(__3349__)
  );
  LUT5 #(
    .INIT(32'h3f00aaaa)
  ) __7033__ (
    .I4(__3349__),
    .I3(__2240__),
    .I2(__2237__),
    .I1(__2224__),
    .I0(__871__),
    .O(__3350__)
  );
  LUT5 #(
    .INIT(32'h0000efff)
  ) __7034__ (
    .I4(g3234),
    .I3(__1508__),
    .I2(__3066__),
    .I1(__1506__),
    .I0(__1507__),
    .O(__3351__)
  );
  LUT4 #(
    .INIT(16'h7df5)
  ) __7035__ (
    .I3(__1623__),
    .I2(__1505__),
    .I1(__215__),
    .I0(__3351__),
    .O(__3352__)
  );
  LUT6 #(
    .INIT(64'h0100000100000000)
  ) __7036__ (
    .I5(__868__),
    .I4(__1828__),
    .I3(__1649__),
    .I2(__1966__),
    .I1(g1943),
    .I0(__867__),
    .O(__3353__)
  );
  LUT6 #(
    .INIT(64'h000000004fff0000)
  ) __7037__ (
    .I5(__968__),
    .I4(__969__),
    .I3(__868__),
    .I2(__2346__),
    .I1(__2551__),
    .I0(__2552__),
    .O(__3354__)
  );
  LUT6 #(
    .INIT(64'hffffffff000f00bb)
  ) __7038__ (
    .I5(__3354__),
    .I4(__2348__),
    .I3(__2347__),
    .I2(__3353__),
    .I1(__2346__),
    .I0(__763__),
    .O(__3355__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __7039__ (
    .I1(__2627__),
    .I0(__928__),
    .O(__3356__)
  );
  LUT6 #(
    .INIT(64'h00000f0f00ff4444)
  ) __7040__ (
    .I5(__1037__),
    .I4(__1036__),
    .I3(__2902__),
    .I2(__2906__),
    .I1(__936__),
    .I0(__3356__),
    .O(__3357__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7041__ (
    .I2(__589__),
    .I1(__2608__),
    .I0(__1271__),
    .O(__3358__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __7042__ (
    .I5(__944__),
    .I4(__764__),
    .I3(__573__),
    .I2(__745__),
    .I1(__685__),
    .I0(__741__),
    .O(__3359__)
  );
  LUT5 #(
    .INIT(32'h00f4f0f0)
  ) __7043__ (
    .I4(__662__),
    .I3(__2143__),
    .I2(__521__),
    .I1(__603__),
    .I0(__2141__),
    .O(__3360__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7044__ (
    .I2(__954__),
    .I1(__2051__),
    .I0(__949__),
    .O(__3361__)
  );
  LUT6 #(
    .INIT(64'h0f0f4444ff00ff00)
  ) __7045__ (
    .I5(__662__),
    .I4(__2653__),
    .I3(__1252__),
    .I2(__2652__),
    .I1(__1428__),
    .I0(__2651__),
    .O(__3362__)
  );
  LUT6 #(
    .INIT(64'h4150c3f05050f0f0)
  ) __7046__ (
    .I5(__944__),
    .I4(__954__),
    .I3(__747__),
    .I2(__802__),
    .I1(__748__),
    .I0(__875__),
    .O(__3363__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7047__ (
    .I2(__1511__),
    .I1(__77__),
    .I0(__218__),
    .O(__3364__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __7048__ (
    .I3(__589__),
    .I2(__2282__),
    .I1(__1617__),
    .I0(__1227__),
    .O(__3365__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7049__ (
    .I2(__944__),
    .I1(__1784__),
    .I0(__1370__),
    .O(__3366__)
  );
  LUT6 #(
    .INIT(64'haa3aaaaaaaaaaaaa)
  ) __7050__ (
    .I5(__954__),
    .I4(__93__),
    .I3(__748__),
    .I2(__73__),
    .I1(__747__),
    .I0(__1050__),
    .O(__3367__)
  );
  LUT6 #(
    .INIT(64'hcc77f0f077ccf0f0)
  ) __7051__ (
    .I5(g3229),
    .I4(__2134__),
    .I3(__1810__),
    .I2(__977__),
    .I1(__1808__),
    .I0(__2030__),
    .O(__3368__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __7052__ (
    .I3(__662__),
    .I2(__603__),
    .I1(__1438__),
    .I0(__844__),
    .O(__3369__)
  );
  LUT4 #(
    .INIT(16'h8000)
  ) __7053__ (
    .I3(__224__),
    .I2(__220__),
    .I1(__222__),
    .I0(__3130__),
    .O(__3370__)
  );
  LUT5 #(
    .INIT(32'h12305af0)
  ) __7054__ (
    .I4(__954__),
    .I3(__219__),
    .I2(__365__),
    .I1(__231__),
    .I0(__3370__),
    .O(__3371__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7055__ (
    .I2(__662__),
    .I1(__2709__),
    .I0(__1265__),
    .O(__3372__)
  );
  LUT5 #(
    .INIT(32'hf000aaaa)
  ) __7056__ (
    .I4(__858__),
    .I3(__988__),
    .I2(__991__),
    .I1(__990__),
    .I0(__1381__),
    .O(__3373__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __7057__ (
    .I5(__858__),
    .I4(__93__),
    .I3(__73__),
    .I2(__748__),
    .I1(__459__),
    .I0(__737__),
    .O(__3374__)
  );
  LUT5 #(
    .INIT(32'h4ecccccc)
  ) __7058__ (
    .I4(__663__),
    .I3(__1598__),
    .I2(__1454__),
    .I1(__1230__),
    .I0(__1635__),
    .O(__3375__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7059__ (
    .I2(__589__),
    .I1(__2709__),
    .I0(__1257__),
    .O(__3376__)
  );
  LUT4 #(
    .INIT(16'haccc)
  ) __7060__ (
    .I3(__662__),
    .I2(__603__),
    .I1(__800__),
    .I0(__1884__),
    .O(__3377__)
  );
  LUT6 #(
    .INIT(64'h4545ff000505ff00)
  ) __7061__ (
    .I5(__858__),
    .I4(__944__),
    .I3(__382__),
    .I2(__1844__),
    .I1(__279__),
    .I0(__1624__),
    .O(__3378__)
  );
  LUT6 #(
    .INIT(64'h4eeeeeeeeeee4eee)
  ) __7062__ (
    .I5(g3229),
    .I4(__1653__),
    .I3(__1652__),
    .I2(__1651__),
    .I1(__818__),
    .I0(__3003__),
    .O(__3379__)
  );
  LUT6 #(
    .INIT(64'h0f005555cccccccc)
  ) __7063__ (
    .I5(__663__),
    .I4(__603__),
    .I3(__2140__),
    .I2(__2137__),
    .I1(__528__),
    .I0(__2136__),
    .O(__3380__)
  );
  LUT4 #(
    .INIT(16'h8000)
  ) __7064__ (
    .I3(__2960__),
    .I2(__2959__),
    .I1(__2957__),
    .I0(__2946__),
    .O(__3381__)
  );
  LUT5 #(
    .INIT(32'h77f0f0f0)
  ) __7065__ (
    .I4(__663__),
    .I3(__603__),
    .I2(__406__),
    .I1(__1777__),
    .I0(__1858__),
    .O(__3382__)
  );
  LUT6 #(
    .INIT(64'hfa000f0fcccccccc)
  ) __7066__ (
    .I5(__589__),
    .I4(__603__),
    .I3(__2462__),
    .I2(__2209__),
    .I1(__598__),
    .I0(__2210__),
    .O(__3383__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __7067__ (
    .I3(__662__),
    .I2(__603__),
    .I1(__1453__),
    .I0(__1337__),
    .O(__3384__)
  );
  LUT4 #(
    .INIT(16'h0080)
  ) __7068__ (
    .I3(__748__),
    .I2(__954__),
    .I1(__93__),
    .I0(__73__),
    .O(__3385__)
  );
  LUT5 #(
    .INIT(32'h3f00aaaa)
  ) __7069__ (
    .I4(__3385__),
    .I3(__3161__),
    .I2(__3159__),
    .I1(__3152__),
    .I0(__1338__),
    .O(__3386__)
  );
  LUT6 #(
    .INIT(64'hd8fad850d850d8fa)
  ) __7070__ (
    .I5(g3229),
    .I4(__1930__),
    .I3(__1928__),
    .I2(__134__),
    .I1(__1932__),
    .I0(__2970__),
    .O(__3387__)
  );
  LUT6 #(
    .INIT(64'hcf300000aaaaaaaa)
  ) __7071__ (
    .I5(__662__),
    .I4(__1999__),
    .I3(__1759__),
    .I2(__1998__),
    .I1(__1992__),
    .I0(__415__),
    .O(__3388__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7072__ (
    .I2(__663__),
    .I1(__2016__),
    .I0(__736__),
    .O(__3389__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7073__ (
    .I2(__589__),
    .I1(__2167__),
    .I0(__659__),
    .O(__3390__)
  );
  LUT6 #(
    .INIT(64'h0000baaaaaaaaaaa)
  ) __7074__ (
    .I5(__954__),
    .I4(__231__),
    .I3(__242__),
    .I2(__370__),
    .I1(__229__),
    .I0(__228__),
    .O(__3391__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __7075__ (
    .I5(__858__),
    .I4(__93__),
    .I3(__73__),
    .I2(__748__),
    .I1(__1040__),
    .I0(__1047__),
    .O(__3392__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __7076__ (
    .I2(__663__),
    .I1(__3320__),
    .I0(__1226__),
    .O(__3393__)
  );
  LUT5 #(
    .INIT(32'ha000cccc)
  ) __7077__ (
    .I4(__944__),
    .I3(__968__),
    .I2(__1646__),
    .I1(__853__),
    .I0(__1648__),
    .O(__3394__)
  );
  LUT6 #(
    .INIT(64'h4545ff000505ff00)
  ) __7078__ (
    .I5(__858__),
    .I4(__954__),
    .I3(__281__),
    .I2(__2117__),
    .I1(__282__),
    .I0(__1624__),
    .O(__3395__)
  );
  LUT6 #(
    .INIT(64'h0f0f4444ff00ff00)
  ) __7079__ (
    .I5(__589__),
    .I4(__2867__),
    .I3(__449__),
    .I2(__2866__),
    .I1(__1412__),
    .I0(__2865__),
    .O(__3396__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __7080__ (
    .I3(__663__),
    .I2(__2282__),
    .I1(__1436__),
    .I0(__777__),
    .O(__3397__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7081__ (
    .I2(__1479__),
    .I1(__1447__),
    .I0(__1463__),
    .O(__3398__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __7082__ (
    .I2(__944__),
    .I1(__445__),
    .I0(__969__),
    .O(__3399__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __7083__ (
    .I2(__663__),
    .I1(__1593__),
    .I0(__1256__),
    .O(__3400__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __7084__ (
    .I5(__944__),
    .I4(__188__),
    .I3(__858__),
    .I2(__187__),
    .I1(__954__),
    .I0(__190__),
    .O(__3401__)
  );
  LUT6 #(
    .INIT(64'hbfffffffa0000000)
  ) __7085__ (
    .I5(__539__),
    .I4(__663__),
    .I3(__603__),
    .I2(__2512__),
    .I1(__2278__),
    .I0(__2277__),
    .O(__3402__)
  );
  LUT5 #(
    .INIT(32'h00eef0f0)
  ) __7086__ (
    .I4(__662__),
    .I3(__3007__),
    .I2(__159__),
    .I1(__3078__),
    .I0(__3076__),
    .O(__3403__)
  );
  LUT6 #(
    .INIT(64'h0f005555cccccccc)
  ) __7087__ (
    .I5(__589__),
    .I4(__603__),
    .I3(__2140__),
    .I2(__2137__),
    .I1(__526__),
    .I0(__2136__),
    .O(__3404__)
  );
  LUT6 #(
    .INIT(64'hfa000f0fcccccccc)
  ) __7088__ (
    .I5(__663__),
    .I4(__603__),
    .I3(__2417__),
    .I2(__2248__),
    .I1(__1128__),
    .I0(__2247__),
    .O(__3405__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7089__ (
    .I2(__2774__),
    .I1(__2788__),
    .I0(__635__),
    .O(__3406__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7090__ (
    .I2(__1812__),
    .I1(__3002__),
    .I0(__859__),
    .O(__3407__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7091__ (
    .I2(__944__),
    .I1(__300__),
    .I0(__1357__),
    .O(__3408__)
  );
  LUT5 #(
    .INIT(32'ha000cccc)
  ) __7092__ (
    .I4(__589__),
    .I3(__1543__),
    .I2(__1544__),
    .I1(__996__),
    .I0(__1542__),
    .O(__3409__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7093__ (
    .I2(__2701__),
    .I1(__2881__),
    .I0(__1219__),
    .O(__3410__)
  );
  LUT5 #(
    .INIT(32'h0030aaaa)
  ) __7094__ (
    .I4(__589__),
    .I3(__1761__),
    .I2(__1760__),
    .I1(__1759__),
    .I0(__187__),
    .O(__3411__)
  );
  LUT6 #(
    .INIT(64'h000000004fff0000)
  ) __7095__ (
    .I5(__1036__),
    .I4(__1037__),
    .I3(__988__),
    .I2(__2627__),
    .I1(__2631__),
    .I0(__2636__),
    .O(__3412__)
  );
  LUT6 #(
    .INIT(64'hffffffff000f00bb)
  ) __7096__ (
    .I5(__3412__),
    .I4(__2630__),
    .I3(__2629__),
    .I2(__2897__),
    .I1(__2627__),
    .I0(__935__),
    .O(__3413__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __7097__ (
    .I5(__954__),
    .I4(__242__),
    .I3(__370__),
    .I2(__229__),
    .I1(__174__),
    .I0(__222__),
    .O(__3414__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __7098__ (
    .I5(__858__),
    .I4(__242__),
    .I3(__370__),
    .I2(__229__),
    .I1(__189__),
    .I0(__224__),
    .O(__3415__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7099__ (
    .I1(__954__),
    .I0(__231__),
    .O(__3416__)
  );
  LUT6 #(
    .INIT(64'h00007fff00008000)
  ) __7100__ (
    .I5(__219__),
    .I4(__3416__),
    .I3(__224__),
    .I2(__220__),
    .I1(__222__),
    .I0(__3130__),
    .O(__3417__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __7101__ (
    .I3(__589__),
    .I2(__603__),
    .I1(__1453__),
    .I0(__1335__),
    .O(__3418__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __7102__ (
    .I3(__663__),
    .I2(__603__),
    .I1(__1460__),
    .I0(__735__),
    .O(__3419__)
  );
  LUT5 #(
    .INIT(32'h12123030)
  ) __7103__ (
    .I4(__1506__),
    .I3(__1508__),
    .I2(__1507__),
    .I1(g3234),
    .I0(__3066__),
    .O(__3420__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7104__ (
    .I2(__589__),
    .I1(__2791__),
    .I0(__1198__),
    .O(__3421__)
  );
  LUT6 #(
    .INIT(64'he4ee4e4e4eeee4e4)
  ) __7105__ (
    .I5(g3229),
    .I4(__1652__),
    .I3(__2269__),
    .I2(__1653__),
    .I1(__821__),
    .I0(__3003__),
    .O(__3422__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __7106__ (
    .I5(__764__),
    .I4(__573__),
    .I3(__858__),
    .I2(__745__),
    .I1(__698__),
    .I0(__750__),
    .O(__3423__)
  );
  LUT5 #(
    .INIT(32'h0030aaaa)
  ) __7107__ (
    .I4(__663__),
    .I3(__1544__),
    .I2(__1543__),
    .I1(__1542__),
    .I0(__1007__),
    .O(__3424__)
  );
  LUT5 #(
    .INIT(32'h00eef0f0)
  ) __7108__ (
    .I4(__662__),
    .I3(__2621__),
    .I2(__1166__),
    .I1(__2725__),
    .I0(__2723__),
    .O(__3425__)
  );
  LUT4 #(
    .INIT(16'haccc)
  ) __7109__ (
    .I3(__663__),
    .I2(__603__),
    .I1(__823__),
    .I0(__1742__),
    .O(__3426__)
  );
  LUT6 #(
    .INIT(64'haa3aaaaaaaaaaaaa)
  ) __7110__ (
    .I5(__858__),
    .I4(__93__),
    .I3(__748__),
    .I2(__73__),
    .I1(__802__),
    .I0(__192__),
    .O(__3427__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __7111__ (
    .I1(__217__),
    .I0(g3234),
    .O(__3428__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7112__ (
    .I2(__663__),
    .I1(__2571__),
    .I0(__1204__),
    .O(__3429__)
  );
  LUT5 #(
    .INIT(32'h0030aaaa)
  ) __7113__ (
    .I4(__663__),
    .I3(__1761__),
    .I2(__1760__),
    .I1(__1759__),
    .I0(__190__),
    .O(__3430__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __7114__ (
    .I5(__944__),
    .I4(__936__),
    .I3(__927__),
    .I2(__924__),
    .I1(__905__),
    .I0(__920__),
    .O(__3431__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7115__ (
    .I2(__662__),
    .I1(__2475__),
    .I0(__535__),
    .O(__3432__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __7116__ (
    .I5(__944__),
    .I4(__242__),
    .I3(__370__),
    .I2(__229__),
    .I1(__153__),
    .I0(__216__),
    .O(__3433__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __7117__ (
    .I3(__589__),
    .I2(__603__),
    .I1(__1446__),
    .I0(__831__),
    .O(__3434__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7118__ (
    .I2(__2370__),
    .I1(__3119__),
    .I0(__578__),
    .O(__3435__)
  );
  LUT6 #(
    .INIT(64'hcc77f0f077ccf0f0)
  ) __7119__ (
    .I5(g3229),
    .I4(__1983__),
    .I3(__1979__),
    .I2(__288__),
    .I1(__1977__),
    .I0(__1976__),
    .O(__3436__)
  );
  LUT6 #(
    .INIT(64'h3fffff3faaaaaaaa)
  ) __7120__ (
    .I5(__3049__),
    .I4(g3229),
    .I3(__1979__),
    .I2(__1978__),
    .I1(__1977__),
    .I0(__283__),
    .O(__3437__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7121__ (
    .I2(__858__),
    .I1(__986__),
    .I0(__1397__),
    .O(__3438__)
  );
  LUT4 #(
    .INIT(16'h125a)
  ) __7122__ (
    .I3(__954__),
    .I2(__224__),
    .I1(__231__),
    .I0(__3130__),
    .O(__3439__)
  );
  LUT6 #(
    .INIT(64'h00007fff00008000)
  ) __7123__ (
    .I5(__1234__),
    .I4(__2151__),
    .I3(__2148__),
    .I2(__1236__),
    .I1(__1235__),
    .I0(__1237__),
    .O(__3440__)
  );
  LUT2 #(
    .INIT(4'he)
  ) __7124__ (
    .I1(g3234),
    .I0(__233__),
    .O(__3441__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __7125__ (
    .I5(__944__),
    .I4(__764__),
    .I3(__573__),
    .I2(__745__),
    .I1(__696__),
    .I0(__750__),
    .O(__3442__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __7126__ (
    .I3(__589__),
    .I2(__603__),
    .I1(__1442__),
    .I0(__837__),
    .O(__3443__)
  );
  LUT4 #(
    .INIT(16'haccc)
  ) __7127__ (
    .I3(__944__),
    .I2(__875__),
    .I1(__1348__),
    .I0(__2056__),
    .O(__3444__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7128__ (
    .I2(__1479__),
    .I1(__1471__),
    .I0(__1459__),
    .O(__3445__)
  );
  LUT5 #(
    .INIT(32'h4ecccccc)
  ) __7129__ (
    .I4(__662__),
    .I3(__1598__),
    .I2(__1438__),
    .I1(__779__),
    .I0(__1635__),
    .O(__3446__)
  );
  LUT5 #(
    .INIT(32'h00f4f0f0)
  ) __7130__ (
    .I4(__589__),
    .I3(__3311__),
    .I2(__544__),
    .I1(__603__),
    .I0(__3310__),
    .O(__3447__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __7131__ (
    .I5(__858__),
    .I4(__936__),
    .I3(__927__),
    .I2(__924__),
    .I1(__910__),
    .I0(__921__),
    .O(__3448__)
  );
  LUT6 #(
    .INIT(64'h0000ffff00001f3f)
  ) __7132__ (
    .I5(__1351__),
    .I4(__2769__),
    .I3(__1352__),
    .I2(__2939__),
    .I1(__2952__),
    .I0(__2955__),
    .O(__3449__)
  );
  LUT4 #(
    .INIT(16'h0008)
  ) __7133__ (
    .I3(__1350__),
    .I2(__1349__),
    .I1(__1351__),
    .I0(__1352__),
    .O(__3450__)
  );
  LUT5 #(
    .INIT(32'haaaaaa2a)
  ) __7134__ (
    .I4(__1532__),
    .I3(__1522__),
    .I2(__2944__),
    .I1(__3450__),
    .I0(__3449__),
    .O(__3451__)
  );
  LUT6 #(
    .INIT(64'hffff0000007f0000)
  ) __7135__ (
    .I5(__1347__),
    .I4(__3451__),
    .I3(__2947__),
    .I2(__1352__),
    .I1(__2944__),
    .I0(__2949__),
    .O(__3452__)
  );
  LUT6 #(
    .INIT(64'h4150c3f05050f0f0)
  ) __7136__ (
    .I5(__944__),
    .I4(__954__),
    .I3(__367__),
    .I2(__366__),
    .I1(__229__),
    .I0(__231__),
    .O(__3453__)
  );
  LUT4 #(
    .INIT(16'h125a)
  ) __7137__ (
    .I3(__954__),
    .I2(__918__),
    .I1(__925__),
    .I0(__2746__),
    .O(__3454__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7138__ (
    .I2(__589__),
    .I1(__2090__),
    .I0(__547__),
    .O(__3455__)
  );
  LUT6 #(
    .INIT(64'haa3aaaaaaaaaaaaa)
  ) __7139__ (
    .I5(__944__),
    .I4(__93__),
    .I3(__748__),
    .I2(__73__),
    .I1(__796__),
    .I0(__1391__),
    .O(__3456__)
  );
  LUT5 #(
    .INIT(32'h00008000)
  ) __7140__ (
    .I4(__229__),
    .I3(__944__),
    .I2(__227__),
    .I1(__366__),
    .I0(__367__),
    .O(__3457__)
  );
  LUT4 #(
    .INIT(16'h125a)
  ) __7141__ (
    .I3(__954__),
    .I2(__225__),
    .I1(__231__),
    .I0(__3457__),
    .O(__3458__)
  );
  LUT5 #(
    .INIT(32'hf8070000)
  ) __7142__ (
    .I4(__2344__),
    .I3(__1649__),
    .I2(__1832__),
    .I1(__2343__),
    .I0(__2342__),
    .O(__3459__)
  );
  LUT6 #(
    .INIT(64'h000033330f0faf00)
  ) __7143__ (
    .I5(__968__),
    .I4(__969__),
    .I3(__764__),
    .I2(__2346__),
    .I1(__3459__),
    .I0(__758__),
    .O(__3460__)
  );
  LUT6 #(
    .INIT(64'hcc77f0f077ccf0f0)
  ) __7144__ (
    .I5(g3229),
    .I4(__2062__),
    .I3(__2065__),
    .I2(__1206__),
    .I1(__2063__),
    .I0(__2679__),
    .O(__3461__)
  );
  LUT6 #(
    .INIT(64'h0100000100000000)
  ) __7145__ (
    .I5(__868__),
    .I4(__1649__),
    .I3(__1820__),
    .I2(__1966__),
    .I1(g1943),
    .I0(__867__),
    .O(__3462__)
  );
  LUT6 #(
    .INIT(64'hffffffff000f00bb)
  ) __7146__ (
    .I5(__2553__),
    .I4(__2348__),
    .I3(__2347__),
    .I2(__3462__),
    .I1(__2346__),
    .I0(__761__),
    .O(__3463__)
  );
  LUT5 #(
    .INIT(32'h44ff00f0)
  ) __7147__ (
    .I4(__1648__),
    .I3(__1647__),
    .I2(__1649__),
    .I1(__968__),
    .I0(__1646__),
    .O(__3464__)
  );
  LUT5 #(
    .INIT(32'h0030aaaa)
  ) __7148__ (
    .I4(__662__),
    .I3(__1681__),
    .I2(__1682__),
    .I1(__1680__),
    .I0(__422__),
    .O(__3465__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7149__ (
    .I2(__662__),
    .I1(__2791__),
    .I0(__1200__),
    .O(__3466__)
  );
  LUT6 #(
    .INIT(64'haa3aaaaaaaaaaaaa)
  ) __7150__ (
    .I5(__944__),
    .I4(__93__),
    .I3(__748__),
    .I2(__73__),
    .I1(__1055__),
    .I0(__794__),
    .O(__3467__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __7151__ (
    .I5(__764__),
    .I4(__573__),
    .I3(__954__),
    .I2(__745__),
    .I1(__701__),
    .I0(__766__),
    .O(__3468__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7152__ (
    .I2(__1511__),
    .I1(__86__),
    .I0(__207__),
    .O(__3469__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7153__ (
    .I2(__1479__),
    .I1(__1465__),
    .I0(__1410__),
    .O(__3470__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __7154__ (
    .I3(__662__),
    .I2(__603__),
    .I1(__1446__),
    .I0(__832__),
    .O(__3471__)
  );
  LUT6 #(
    .INIT(64'hbfffffffa0000000)
  ) __7155__ (
    .I5(__1187__),
    .I4(__589__),
    .I3(__603__),
    .I2(__2585__),
    .I1(__2509__),
    .I0(__2508__),
    .O(__3472__)
  );
  LUT6 #(
    .INIT(64'he4ee4e4e4eeee4e4)
  ) __7156__ (
    .I5(g3229),
    .I4(__1652__),
    .I3(__2269__),
    .I2(__1653__),
    .I1(__564__),
    .I0(__1650__),
    .O(__3473__)
  );
  LUT4 #(
    .INIT(16'h11f0)
  ) __7157__ (
    .I3(__662__),
    .I2(__460__),
    .I1(__3007__),
    .I0(__3006__),
    .O(__3474__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7158__ (
    .I2(__662__),
    .I1(__2367__),
    .I0(__721__),
    .O(__3475__)
  );
  LUT6 #(
    .INIT(64'hd8fad850d850d8fa)
  ) __7159__ (
    .I5(g3229),
    .I4(__1810__),
    .I3(__1809__),
    .I2(__982__),
    .I1(__1808__),
    .I0(__2489__),
    .O(__3476__)
  );
  LUT6 #(
    .INIT(64'h00007fff00008000)
  ) __7160__ (
    .I5(__641__),
    .I4(__2151__),
    .I3(__642__),
    .I2(__643__),
    .I1(__644__),
    .I0(__2591__),
    .O(__3477__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __7161__ (
    .I5(__954__),
    .I4(__242__),
    .I3(__370__),
    .I2(__229__),
    .I1(__157__),
    .I0(__365__),
    .O(__3478__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __7162__ (
    .I3(__589__),
    .I2(__2282__),
    .I1(__1643__),
    .I0(__1277__),
    .O(__3479__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __7163__ (
    .I3(__662__),
    .I2(__603__),
    .I1(__1410__),
    .I0(__453__),
    .O(__3480__)
  );
  LUT6 #(
    .INIT(64'h3fffff3faaaaaaaa)
  ) __7164__ (
    .I5(__2370__),
    .I4(g3229),
    .I3(__2287__),
    .I2(__2286__),
    .I1(__2285__),
    .I0(__557__),
    .O(__3481__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __7165__ (
    .I1(__1496__),
    .I0(g51),
    .O(__3482__)
  );
  LUT6 #(
    .INIT(64'h00007fff00008000)
  ) __7166__ (
    .I5(__570__),
    .I4(__2151__),
    .I3(__2148__),
    .I2(__571__),
    .I1(__606__),
    .I0(__607__),
    .O(__3483__)
  );
  LUT4 #(
    .INIT(16'h11f0)
  ) __7167__ (
    .I3(__663__),
    .I2(__543__),
    .I1(__3007__),
    .I0(__3006__),
    .O(__3484__)
  );
  LUT4 #(
    .INIT(16'haccc)
  ) __7168__ (
    .I3(__858__),
    .I2(__925__),
    .I1(__880__),
    .I0(__1805__),
    .O(__3485__)
  );
  LUT6 #(
    .INIT(64'h3fffff3faaaaaaaa)
  ) __7169__ (
    .I5(__2701__),
    .I4(g3229),
    .I3(__2065__),
    .I2(__2063__),
    .I1(__2064__),
    .I0(__1199__),
    .O(__3486__)
  );
  LUT6 #(
    .INIT(64'hbfffffffa0000000)
  ) __7170__ (
    .I5(__1123__),
    .I4(__663__),
    .I3(__603__),
    .I2(__2417__),
    .I1(__2247__),
    .I0(__2248__),
    .O(__3487__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __7171__ (
    .I2(__944__),
    .I1(__1038__),
    .I0(__1037__),
    .O(__3488__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7172__ (
    .I2(__944__),
    .I1(__140__),
    .I0(__1388__),
    .O(__3489__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __7173__ (
    .I5(__764__),
    .I4(__573__),
    .I3(__858__),
    .I2(__745__),
    .I1(__706__),
    .I0(__767__),
    .O(__3490__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7174__ (
    .I2(__1479__),
    .I1(__1475__),
    .I0(__1455__),
    .O(__3491__)
  );
  LUT5 #(
    .INIT(32'h0030aaaa)
  ) __7175__ (
    .I4(__589__),
    .I3(__1760__),
    .I2(__1761__),
    .I1(__1759__),
    .I0(__191__),
    .O(__3492__)
  );
  LUT5 #(
    .INIT(32'h0030aaaa)
  ) __7176__ (
    .I4(__662__),
    .I3(__1761__),
    .I2(__1760__),
    .I1(__1759__),
    .I0(__188__),
    .O(__3493__)
  );
  LUT5 #(
    .INIT(32'h0030aaaa)
  ) __7177__ (
    .I4(__662__),
    .I3(__1597__),
    .I2(__1596__),
    .I1(__1595__),
    .I0(__435__),
    .O(__3494__)
  );
  LUT4 #(
    .INIT(16'haccc)
  ) __7178__ (
    .I3(__944__),
    .I2(__231__),
    .I1(__285__),
    .I0(__1982__),
    .O(__3495__)
  );
  LUT5 #(
    .INIT(32'h06666666)
  ) __7179__ (
    .I4(__589__),
    .I3(__1598__),
    .I2(__603__),
    .I1(__1174__),
    .I0(__1874__),
    .O(__3496__)
  );
  LUT5 #(
    .INIT(32'h00f4f0f0)
  ) __7180__ (
    .I4(__662__),
    .I3(__2661__),
    .I2(__647__),
    .I1(__603__),
    .I0(__2660__),
    .O(__3497__)
  );
  LUT6 #(
    .INIT(64'h0000bfff00000000)
  ) __7181__ (
    .I5(g3233),
    .I4(g3230),
    .I3(__1352__),
    .I2(__2939__),
    .I1(__2942__),
    .I0(__1344__),
    .O(__3498__)
  );
  LUT4 #(
    .INIT(16'haccc)
  ) __7182__ (
    .I3(__944__),
    .I2(__925__),
    .I1(__878__),
    .I0(__1805__),
    .O(__3499__)
  );
  LUT5 #(
    .INIT(32'h00008000)
  ) __7183__ (
    .I4(__748__),
    .I3(__944__),
    .I2(__799__),
    .I1(__747__),
    .I0(__802__),
    .O(__3500__)
  );
  LUT4 #(
    .INIT(16'h125a)
  ) __7184__ (
    .I3(__954__),
    .I2(__1051__),
    .I1(__875__),
    .I0(__3500__),
    .O(__3501__)
  );
  LUT6 #(
    .INIT(64'h00f07878f0f0f0f0)
  ) __7185__ (
    .I5(__589__),
    .I4(__1598__),
    .I3(__603__),
    .I2(__606__),
    .I1(__571__),
    .I0(__607__),
    .O(__3502__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __7186__ (
    .I3(__663__),
    .I2(__603__),
    .I1(__1410__),
    .I0(__655__),
    .O(__3503__)
  );
  LUT5 #(
    .INIT(32'h77f0f0f0)
  ) __7187__ (
    .I4(__589__),
    .I3(__603__),
    .I2(__467__),
    .I1(__1731__),
    .I0(__1715__),
    .O(__3504__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __7188__ (
    .I3(__662__),
    .I2(__603__),
    .I1(__1456__),
    .I0(__1117__),
    .O(__3505__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __7189__ (
    .I2(g3229),
    .I1(__1112__),
    .I0(__1110__),
    .O(__3506__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7190__ (
    .I2(__954__),
    .I1(__142__),
    .I0(__1365__),
    .O(__3507__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __7191__ (
    .I3(__589__),
    .I2(__603__),
    .I1(__1422__),
    .I0(__1319__),
    .O(__3508__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7192__ (
    .I2(__589__),
    .I1(__2571__),
    .I0(__1160__),
    .O(__3509__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7193__ (
    .I2(__663__),
    .I1(__2743__),
    .I0(__428__),
    .O(__3510__)
  );
  LUT5 #(
    .INIT(32'hb8f0f0f0)
  ) __7194__ (
    .I4(__662__),
    .I3(__1598__),
    .I2(__783__),
    .I1(__1635__),
    .I0(__2455__),
    .O(__3511__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __7195__ (
    .I2(__662__),
    .I1(__2327__),
    .I0(__1218__),
    .O(__3512__)
  );
  LUT6 #(
    .INIT(64'h0000077007700000)
  ) __7196__ (
    .I5(__1886__),
    .I4(__1176__),
    .I3(__1883__),
    .I2(__1048__),
    .I1(__1892__),
    .I0(__1043__),
    .O(__3513__)
  );
  LUT6 #(
    .INIT(64'h00000eee0eee0000)
  ) __7197__ (
    .I5(__1890__),
    .I4(__1161__),
    .I3(__1888__),
    .I2(__1164__),
    .I1(__1892__),
    .I0(__1043__),
    .O(__3514__)
  );
  LUT5 #(
    .INIT(32'heee0eeee)
  ) __7198__ (
    .I4(__1597__),
    .I3(__1596__),
    .I2(__1595__),
    .I1(__1879__),
    .I0(__1174__),
    .O(__3515__)
  );
  LUT6 #(
    .INIT(64'h0000077707770000)
  ) __7199__ (
    .I5(__1895__),
    .I4(__1175__),
    .I3(__1879__),
    .I2(__1174__),
    .I1(__1877__),
    .I0(__1180__),
    .O(__3516__)
  );
  LUT6 #(
    .INIT(64'h0e00000000000000)
  ) __7200__ (
    .I5(__3516__),
    .I4(__3515__),
    .I3(__3514__),
    .I2(__1598__),
    .I1(__1888__),
    .I0(__1164__),
    .O(__3517__)
  );
  LUT4 #(
    .INIT(16'h0ee0)
  ) __7201__ (
    .I3(__1881__),
    .I2(__730__),
    .I1(__1877__),
    .I0(__1180__),
    .O(__3518__)
  );
  LUT6 #(
    .INIT(64'h155555559fffffff)
  ) __7202__ (
    .I5(__2008__),
    .I4(__3518__),
    .I3(__3517__),
    .I2(__3513__),
    .I1(__1178__),
    .I0(__1897__),
    .O(__3519__)
  );
  LUT5 #(
    .INIT(32'ha000cccc)
  ) __7203__ (
    .I4(__662__),
    .I3(__1682__),
    .I2(__1681__),
    .I1(__309__),
    .I0(__1680__),
    .O(__3520__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7204__ (
    .I2(__858__),
    .I1(__142__),
    .I0(__1366__),
    .O(__3521__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7205__ (
    .I2(__663__),
    .I1(__2641__),
    .I0(__1162__),
    .O(__3522__)
  );
  LUT5 #(
    .INIT(32'h00eef0f0)
  ) __7206__ (
    .I4(__589__),
    .I3(__2621__),
    .I2(__1163__),
    .I1(__2725__),
    .I0(__2723__),
    .O(__3523__)
  );
  LUT6 #(
    .INIT(64'hd8fad850d850d8fa)
  ) __7207__ (
    .I5(g3229),
    .I4(__1602__),
    .I3(__1601__),
    .I2(__1136__),
    .I1(__1600__),
    .I0(__1633__),
    .O(__3524__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __7208__ (
    .I3(__589__),
    .I2(__603__),
    .I1(__1458__),
    .I0(__1306__),
    .O(__3525__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __7209__ (
    .I2(__663__),
    .I1(__1640__),
    .I0(__1010__),
    .O(__3526__)
  );
  LUT5 #(
    .INIT(32'h12305af0)
  ) __7210__ (
    .I4(__954__),
    .I3(__767__),
    .I2(__766__),
    .I1(__752__),
    .I0(__2613__),
    .O(__3527__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __7211__ (
    .I3(__589__),
    .I2(__603__),
    .I1(__1408__),
    .I0(__425__),
    .O(__3528__)
  );
  LUT6 #(
    .INIT(64'h0f005555cccccccc)
  ) __7212__ (
    .I5(__663__),
    .I4(__603__),
    .I3(__1643__),
    .I2(__1637__),
    .I1(__1186__),
    .I0(__1638__),
    .O(__3529__)
  );
  LUT6 #(
    .INIT(64'ha3aaaaaaaaaaaaaa)
  ) __7213__ (
    .I5(__954__),
    .I4(__93__),
    .I3(__73__),
    .I2(__748__),
    .I1(__788__),
    .I0(__801__),
    .O(__3530__)
  );
  LUT4 #(
    .INIT(16'h11f0)
  ) __7214__ (
    .I3(__663__),
    .I2(__791__),
    .I1(__2764__),
    .I0(__3000__),
    .O(__3531__)
  );
  LUT6 #(
    .INIT(64'h00007fff00008000)
  ) __7215__ (
    .I5(__1048__),
    .I4(__2151__),
    .I3(__730__),
    .I2(__1161__),
    .I1(__1164__),
    .I0(__2924__),
    .O(__3532__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7216__ (
    .I2(__589__),
    .I1(__2367__),
    .I0(__720__),
    .O(__3533__)
  );
  LUT4 #(
    .INIT(16'haccc)
  ) __7217__ (
    .I3(__944__),
    .I2(__875__),
    .I1(__855__),
    .I0(__1951__),
    .O(__3534__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __7218__ (
    .I3(__662__),
    .I2(__603__),
    .I1(__1444__),
    .I0(__835__),
    .O(__3535__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __7219__ (
    .I3(__662__),
    .I2(__603__),
    .I1(__1414__),
    .I0(__235__),
    .O(__3536__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __7220__ (
    .I3(__662__),
    .I2(__603__),
    .I1(__1411__),
    .I0(__440__),
    .O(__3537__)
  );
  LUT6 #(
    .INIT(64'h55555d5500000800)
  ) __7221__ (
    .I5(__590__),
    .I4(__1413__),
    .I3(__1411__),
    .I2(__1412__),
    .I1(__1414__),
    .I0(__2407__),
    .O(__3538__)
  );
  LUT6 #(
    .INIT(64'hd8fad850d850d8fa)
  ) __7222__ (
    .I5(g3229),
    .I4(__1979__),
    .I3(__1978__),
    .I2(__291__),
    .I1(__1977__),
    .I0(__1983__),
    .O(__3539__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __7223__ (
    .I2(__944__),
    .I1(__273__),
    .I0(__269__),
    .O(__3540__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __7224__ (
    .I5(__954__),
    .I4(__936__),
    .I3(__927__),
    .I2(__924__),
    .I1(__900__),
    .I0(__917__),
    .O(__3541__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7225__ (
    .I2(__662__),
    .I1(__3058__),
    .I0(__355__),
    .O(__3542__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __7226__ (
    .I2(__662__),
    .I1(__2357__),
    .I0(__709__),
    .O(__3543__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __7227__ (
    .I5(__858__),
    .I4(__936__),
    .I3(__927__),
    .I2(__924__),
    .I1(__889__),
    .I0(__913__),
    .O(__3544__)
  );
  LUT6 #(
    .INIT(64'h0f005555cccccccc)
  ) __7228__ (
    .I5(__662__),
    .I4(__603__),
    .I3(__1643__),
    .I2(__1637__),
    .I1(__1185__),
    .I0(__1638__),
    .O(__3545__)
  );
  LUT6 #(
    .INIT(64'h4545ff000505ff00)
  ) __7229__ (
    .I5(__858__),
    .I4(__944__),
    .I3(__116__),
    .I2(__1949__),
    .I1(__121__),
    .I0(__1624__),
    .O(__3546__)
  );
  LUT6 #(
    .INIT(64'hbfffffffa0000000)
  ) __7230__ (
    .I5(__552__),
    .I4(__663__),
    .I3(__603__),
    .I2(__2462__),
    .I1(__2210__),
    .I0(__2209__),
    .O(__3547__)
  );
  LUT4 #(
    .INIT(16'h8040)
  ) __7231__ (
    .I3(__2226__),
    .I2(__988__),
    .I1(__2627__),
    .I0(__1805__),
    .O(__3548__)
  );
  LUT6 #(
    .INIT(64'hffffffff000f00bb)
  ) __7232__ (
    .I5(__3412__),
    .I4(__2630__),
    .I3(__2629__),
    .I2(__3548__),
    .I1(__2627__),
    .I0(__932__),
    .O(__3549__)
  );
  LUT6 #(
    .INIT(64'h0000baaaaaaaaaaa)
  ) __7233__ (
    .I5(__858__),
    .I4(__231__),
    .I3(__242__),
    .I2(__370__),
    .I1(__229__),
    .I0(__213__),
    .O(__3550__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __7234__ (
    .I2(__663__),
    .I1(__2019__),
    .I0(__742__),
    .O(__3551__)
  );
  LUT4 #(
    .INIT(16'haccc)
  ) __7235__ (
    .I3(__662__),
    .I2(__603__),
    .I1(__342__),
    .I0(__1893__),
    .O(__3552__)
  );
  LUT5 #(
    .INIT(32'h00f4f0f0)
  ) __7236__ (
    .I4(__589__),
    .I3(__2143__),
    .I2(__509__),
    .I1(__603__),
    .I0(__2141__),
    .O(__3553__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __7237__ (
    .I5(__944__),
    .I4(__200__),
    .I3(__858__),
    .I2(__198__),
    .I1(__954__),
    .I0(__203__),
    .O(__3554__)
  );
  LUT5 #(
    .INIT(32'h00000001)
  ) __7238__ (
    .I4(__297__),
    .I3(g2637),
    .I2(__1784__),
    .I1(__2646__),
    .I0(__371__),
    .O(__3555__)
  );
  LUT6 #(
    .INIT(64'h000000330f0f00aa)
  ) __7239__ (
    .I5(__354__),
    .I4(__356__),
    .I3(__3555__),
    .I2(__2810__),
    .I1(__2816__),
    .I0(__242__),
    .O(__3556__)
  );
  LUT6 #(
    .INIT(64'h0f0f4444ff00ff00)
  ) __7240__ (
    .I5(__662__),
    .I4(__2516__),
    .I3(__1216__),
    .I2(__2515__),
    .I1(__1458__),
    .I0(__2514__),
    .O(__3557__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __7241__ (
    .I3(__589__),
    .I2(__603__),
    .I1(__1414__),
    .I0(__591__),
    .O(__3558__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __7242__ (
    .I2(__944__),
    .I1(__2126__),
    .I0(__943__),
    .O(__3559__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __7243__ (
    .I2(__663__),
    .I1(__2290__),
    .I0(__611__),
    .O(__3560__)
  );
  LUT6 #(
    .INIT(64'h3fffff3faaaaaaaa)
  ) __7244__ (
    .I5(__1983__),
    .I4(g3229),
    .I3(__1979__),
    .I2(__1978__),
    .I1(__1977__),
    .I0(__284__),
    .O(__3561__)
  );
  LUT6 #(
    .INIT(64'h0100000100000000)
  ) __7245__ (
    .I5(__868__),
    .I4(__1646__),
    .I3(__1824__),
    .I2(__1966__),
    .I1(g1943),
    .I0(__867__),
    .O(__3562__)
  );
  LUT6 #(
    .INIT(64'hffffffff000f00bb)
  ) __7246__ (
    .I5(__3354__),
    .I4(__2348__),
    .I3(__2347__),
    .I2(__3562__),
    .I1(__2346__),
    .I0(__759__),
    .O(__3563__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __7247__ (
    .I2(__589__),
    .I1(__2411__),
    .I0(__438__),
    .O(__3564__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7248__ (
    .I2(__954__),
    .I1(__867__),
    .I0(__1386__),
    .O(__3565__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __7249__ (
    .I3(__662__),
    .I2(__603__),
    .I1(__1432__),
    .I0(__1296__),
    .O(__3566__)
  );
  LUT5 #(
    .INIT(32'h00eef0f0)
  ) __7250__ (
    .I4(__589__),
    .I3(__2764__),
    .I2(__1086__),
    .I1(__3102__),
    .I0(__3100__),
    .O(__3567__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __7251__ (
    .I3(__589__),
    .I2(__2282__),
    .I1(__2089__),
    .I0(__463__),
    .O(__3568__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __7252__ (
    .I2(__644__),
    .I1(__645__),
    .I0(__2978__),
    .O(__3569__)
  );
  LUT6 #(
    .INIT(64'h00007fff00008000)
  ) __7253__ (
    .I5(__640__),
    .I4(__2151__),
    .I3(__642__),
    .I2(__643__),
    .I1(__3569__),
    .I0(__641__),
    .O(__3570__)
  );
  LUT6 #(
    .INIT(64'h00007fff00008000)
  ) __7254__ (
    .I5(__567__),
    .I4(__2151__),
    .I3(__605__),
    .I2(__604__),
    .I1(__568__),
    .I0(__2149__),
    .O(__3571__)
  );
  LUT5 #(
    .INIT(32'h0030aaaa)
  ) __7255__ (
    .I4(__663__),
    .I3(__1596__),
    .I2(__1597__),
    .I1(__1595__),
    .I0(__426__),
    .O(__3572__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __7256__ (
    .I2(__858__),
    .I1(__2058__),
    .I0(__109__),
    .O(__3573__)
  );
  LUT5 #(
    .INIT(32'h007f0080)
  ) __7257__ (
    .I4(__642__),
    .I3(__2151__),
    .I2(__643__),
    .I1(__644__),
    .I0(__2591__),
    .O(__3574__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __7258__ (
    .I5(__944__),
    .I4(__242__),
    .I3(__370__),
    .I2(__229__),
    .I1(__170__),
    .I0(__220__),
    .O(__3575__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __7259__ (
    .I5(__954__),
    .I4(__242__),
    .I3(__370__),
    .I2(__229__),
    .I1(__197__),
    .I0(__225__),
    .O(__3576__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7260__ (
    .I2(__858__),
    .I1(__1784__),
    .I0(__1372__),
    .O(__3577__)
  );
  LUT6 #(
    .INIT(64'haa3aaaaaaaaaaaaa)
  ) __7261__ (
    .I5(__944__),
    .I4(__93__),
    .I3(__748__),
    .I2(__73__),
    .I1(__747__),
    .I0(__789__),
    .O(__3578__)
  );
  LUT4 #(
    .INIT(16'haccc)
  ) __7262__ (
    .I3(__589__),
    .I2(__603__),
    .I1(__374__),
    .I0(__1712__),
    .O(__3579__)
  );
  LUT4 #(
    .INIT(16'haccc)
  ) __7263__ (
    .I3(__662__),
    .I2(__603__),
    .I1(__817__),
    .I0(__1751__),
    .O(__3580__)
  );
  LUT5 #(
    .INIT(32'h00f4f0f0)
  ) __7264__ (
    .I4(__662__),
    .I3(__3311__),
    .I2(__545__),
    .I1(__603__),
    .I0(__3310__),
    .O(__3581__)
  );
  LUT5 #(
    .INIT(32'h4ecccccc)
  ) __7265__ (
    .I4(__662__),
    .I3(__1598__),
    .I2(__1408__),
    .I1(__585__),
    .I0(__1635__),
    .O(__3582__)
  );
  LUT6 #(
    .INIT(64'h132033005fa0ff00)
  ) __7266__ (
    .I5(__954__),
    .I4(__365__),
    .I3(__216__),
    .I2(__219__),
    .I1(__231__),
    .I0(__3370__),
    .O(__3583__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7267__ (
    .I2(__2970__),
    .I1(__2676__),
    .I0(__138__),
    .O(__3584__)
  );
  LUT6 #(
    .INIT(64'hbfffffffa0000000)
  ) __7268__ (
    .I5(__529__),
    .I4(__589__),
    .I3(__603__),
    .I2(__2512__),
    .I1(__2278__),
    .I0(__2277__),
    .O(__3585__)
  );
  LUT5 #(
    .INIT(32'h0030aaaa)
  ) __7269__ (
    .I4(__662__),
    .I3(__1760__),
    .I2(__1761__),
    .I1(__1759__),
    .I0(__195__),
    .O(__3586__)
  );
  LUT5 #(
    .INIT(32'h0030aaaa)
  ) __7270__ (
    .I4(__663__),
    .I3(__1543__),
    .I2(__1544__),
    .I1(__1542__),
    .I0(__1004__),
    .O(__3587__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7271__ (
    .I2(__858__),
    .I1(__140__),
    .I0(__1394__),
    .O(__3588__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __7272__ (
    .I5(__858__),
    .I4(__242__),
    .I3(__370__),
    .I2(__229__),
    .I1(__338__),
    .I0(__365__),
    .O(__3589__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __7273__ (
    .I2(__662__),
    .I1(__3320__),
    .I0(__1225__),
    .O(__3590__)
  );
  LUT6 #(
    .INIT(64'h000033330f0faf00)
  ) __7274__ (
    .I5(__1036__),
    .I4(__1037__),
    .I3(__936__),
    .I2(__2627__),
    .I1(__2903__),
    .I0(__930__),
    .O(__3591__)
  );
  LUT5 #(
    .INIT(32'ha000cccc)
  ) __7275__ (
    .I4(__944__),
    .I3(__1981__),
    .I2(__354__),
    .I1(__145__),
    .I0(__1800__),
    .O(__3592__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __7276__ (
    .I3(__662__),
    .I2(__2282__),
    .I1(__2089__),
    .I0(__464__),
    .O(__3593__)
  );
  LUT6 #(
    .INIT(64'h0f0f4444ff00ff00)
  ) __7277__ (
    .I5(__589__),
    .I4(__2526__),
    .I3(__711__),
    .I2(__2525__),
    .I1(__1446__),
    .I0(__2524__),
    .O(__3594__)
  );
  LUT5 #(
    .INIT(32'ha000cccc)
  ) __7278__ (
    .I4(__662__),
    .I3(__1543__),
    .I2(__1544__),
    .I1(__997__),
    .I0(__1542__),
    .O(__3595__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7279__ (
    .I2(__944__),
    .I1(__986__),
    .I0(__1395__),
    .O(__3596__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7280__ (
    .I2(__858__),
    .I1(__868__),
    .I0(__1362__),
    .O(__3597__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __7281__ (
    .I5(__954__),
    .I4(__936__),
    .I3(__927__),
    .I2(__924__),
    .I1(__894__),
    .I0(__915__),
    .O(__3598__)
  );
  LUT5 #(
    .INIT(32'h77f0f0f0)
  ) __7282__ (
    .I4(__589__),
    .I3(__603__),
    .I2(__404__),
    .I1(__1777__),
    .I0(__1858__),
    .O(__3599__)
  );
  LUT6 #(
    .INIT(64'hcc77f0f077ccf0f0)
  ) __7283__ (
    .I5(g3229),
    .I4(__1807__),
    .I3(__1810__),
    .I2(__978__),
    .I1(__1808__),
    .I0(__2030__),
    .O(__3600__)
  );
  LUT6 #(
    .INIT(64'haaaacaaaaaaaaaaa)
  ) __7284__ (
    .I5(__944__),
    .I4(__229__),
    .I3(__242__),
    .I2(__370__),
    .I1(__2425__),
    .I0(__147__),
    .O(__3601__)
  );
  LUT4 #(
    .INIT(16'haccc)
  ) __7285__ (
    .I3(__944__),
    .I2(__752__),
    .I1(__676__),
    .I0(__1646__),
    .O(__3602__)
  );
  LUT6 #(
    .INIT(64'haa000000000f33ff)
  ) __7286__ (
    .I5(__1351__),
    .I4(__1350__),
    .I3(__1349__),
    .I2(__2937__),
    .I1(__3265__),
    .I0(__1381__),
    .O(__3603__)
  );
  LUT5 #(
    .INIT(32'h4ecccccc)
  ) __7287__ (
    .I4(__662__),
    .I3(__1598__),
    .I2(__1407__),
    .I1(__437__),
    .I0(__1635__),
    .O(__3604__)
  );
  LUT6 #(
    .INIT(64'h0f005555cccccccc)
  ) __7288__ (
    .I5(__662__),
    .I4(__603__),
    .I3(__2089__),
    .I2(__2084__),
    .I1(__550__),
    .I0(__2085__),
    .O(__3605__)
  );
  LUT6 #(
    .INIT(64'h55555d5500000800)
  ) __7289__ (
    .I5(__1231__),
    .I4(__1458__),
    .I3(__1460__),
    .I2(__1459__),
    .I1(__1457__),
    .I0(__1964__),
    .O(__3606__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __7290__ (
    .I3(__589__),
    .I2(__603__),
    .I1(__1409__),
    .I0(__471__),
    .O(__3607__)
  );
  LUT6 #(
    .INIT(64'hd8fad850d850d8fa)
  ) __7291__ (
    .I5(g3229),
    .I4(__1653__),
    .I3(__1651__),
    .I2(__864__),
    .I1(__1652__),
    .I0(__1650__),
    .O(__3608__)
  );
  LUT5 #(
    .INIT(32'h4ecccccc)
  ) __7292__ (
    .I4(__589__),
    .I3(__1598__),
    .I2(__1453__),
    .I1(__1258__),
    .I0(__1635__),
    .O(__3609__)
  );
  LUT5 #(
    .INIT(32'h44ff00f0)
  ) __7293__ (
    .I4(__1981__),
    .I3(__1647__),
    .I2(__1982__),
    .I1(__354__),
    .I0(__1800__),
    .O(__3610__)
  );
  LUT6 #(
    .INIT(64'h5455555555555555)
  ) __7294__ (
    .I5(__1483__),
    .I4(__1486__),
    .I3(__1611__),
    .I2(__1484__),
    .I1(__1485__),
    .I0(__1497__),
    .O(__3611__)
  );
  LUT3 #(
    .INIT(8'h6f)
  ) __7295__ (
    .I2(__3611__),
    .I1(__1486__),
    .I0(__1611__),
    .O(__3612__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7296__ (
    .I2(__663__),
    .I1(__2475__),
    .I0(__1221__),
    .O(__3613__)
  );
  LUT6 #(
    .INIT(64'h000f00ab000fffab)
  ) __7297__ (
    .I5(__2812__),
    .I4(__2646__),
    .I3(__2645__),
    .I2(__2818__),
    .I1(__1802__),
    .I0(__372__),
    .O(__3614__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7298__ (
    .I2(__858__),
    .I1(__2397__),
    .I0(__809__),
    .O(__3615__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7299__ (
    .I2(__1807__),
    .I1(__2962__),
    .I0(__984__),
    .O(__3616__)
  );
  LUT6 #(
    .INIT(64'hd8fad850d850d8fa)
  ) __7300__ (
    .I5(g3229),
    .I4(__1979__),
    .I3(__1978__),
    .I2(__293__),
    .I1(__1977__),
    .I0(__2244__),
    .O(__3617__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __7301__ (
    .I3(__589__),
    .I2(__603__),
    .I1(__1430__),
    .I0(__1298__),
    .O(__3618__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __7302__ (
    .I3(__663__),
    .I2(__603__),
    .I1(__1440__),
    .I0(__842__),
    .O(__3619__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7303__ (
    .I2(__954__),
    .I1(__140__),
    .I0(__1389__),
    .O(__3620__)
  );
  LUT6 #(
    .INIT(64'h0078787878787878)
  ) __7304__ (
    .I5(__589__),
    .I4(__1598__),
    .I3(__603__),
    .I2(__1228__),
    .I1(__1232__),
    .I0(__2075__),
    .O(__3621__)
  );
  LUT6 #(
    .INIT(64'hfa000f0fcccccccc)
  ) __7305__ (
    .I5(__589__),
    .I4(__603__),
    .I3(__2417__),
    .I2(__2248__),
    .I1(__1126__),
    .I0(__2247__),
    .O(__3622__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7306__ (
    .I2(__2244__),
    .I1(__1980__),
    .I0(__296__),
    .O(__3623__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __7307__ (
    .I5(__858__),
    .I4(__242__),
    .I3(__370__),
    .I2(__229__),
    .I1(__154__),
    .I0(__216__),
    .O(__3624__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __7308__ (
    .I5(__954__),
    .I4(__242__),
    .I3(__370__),
    .I2(__229__),
    .I1(__186__),
    .I0(__224__),
    .O(__3625__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __7309__ (
    .I5(__944__),
    .I4(__242__),
    .I3(__370__),
    .I2(__229__),
    .I1(__201__),
    .I0(__227__),
    .O(__3626__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7310__ (
    .I2(__589__),
    .I1(__2016__),
    .I0(__793__),
    .O(__3627__)
  );
  LUT6 #(
    .INIT(64'h55555d5500000800)
  ) __7311__ (
    .I5(__781__),
    .I4(__1448__),
    .I3(__1444__),
    .I2(__1446__),
    .I1(__1450__),
    .I0(__1964__),
    .O(__3628__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7312__ (
    .I2(__858__),
    .I1(__1953__),
    .I0(__112__),
    .O(__3629__)
  );
  LUT6 #(
    .INIT(64'hcc77f0f077ccf0f0)
  ) __7313__ (
    .I5(g3229),
    .I4(__2774__),
    .I3(__2070__),
    .I2(__629__),
    .I1(__2069__),
    .I0(__2581__),
    .O(__3630__)
  );
  LUT6 #(
    .INIT(64'hffffffff000f00bb)
  ) __7314__ (
    .I5(__2637__),
    .I4(__2630__),
    .I3(__2629__),
    .I2(__2898__),
    .I1(__2627__),
    .I0(__933__),
    .O(__3631__)
  );
  LUT4 #(
    .INIT(16'h0080)
  ) __7315__ (
    .I3(__748__),
    .I2(__858__),
    .I1(__93__),
    .I0(__73__),
    .O(__3632__)
  );
  LUT5 #(
    .INIT(32'h3f00aaaa)
  ) __7316__ (
    .I4(__3632__),
    .I3(__3161__),
    .I2(__3159__),
    .I1(__3152__),
    .I0(__1340__),
    .O(__3633__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7317__ (
    .I2(__589__),
    .I1(__3058__),
    .I0(__451__),
    .O(__3634__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7318__ (
    .I2(__1511__),
    .I1(__129__),
    .I0(__171__),
    .O(__3635__)
  );
  LUT6 #(
    .INIT(64'h000a000c00000000)
  ) __7319__ (
    .I5(__764__),
    .I4(g3229),
    .I3(__968__),
    .I2(__969__),
    .I1(__754__),
    .I0(__573__),
    .O(__3636__)
  );
  LUT3 #(
    .INIT(8'h07)
  ) __7320__ (
    .I2(__1818__),
    .I1(__2343__),
    .I0(__2342__),
    .O(__3637__)
  );
  LUT6 #(
    .INIT(64'h6996000000000000)
  ) __7321__ (
    .I5(__2344__),
    .I4(__969__),
    .I3(__1646__),
    .I2(__1649__),
    .I1(__3083__),
    .I0(__3637__),
    .O(__3638__)
  );
  LUT3 #(
    .INIT(8'h07)
  ) __7322__ (
    .I2(__1823__),
    .I1(__2343__),
    .I0(__2342__),
    .O(__3639__)
  );
  LUT3 #(
    .INIT(8'h07)
  ) __7323__ (
    .I2(__1832__),
    .I1(__2343__),
    .I0(__2342__),
    .O(__3640__)
  );
  LUT4 #(
    .INIT(16'hf807)
  ) __7324__ (
    .I3(__1646__),
    .I2(__1826__),
    .I1(__2343__),
    .I0(__2342__),
    .O(__3641__)
  );
  LUT5 #(
    .INIT(32'h7dd78228)
  ) __7325__ (
    .I4(__3081__),
    .I3(__3641__),
    .I2(__3640__),
    .I1(__3639__),
    .I0(__2344__),
    .O(__3642__)
  );
  LUT4 #(
    .INIT(16'h6996)
  ) __7326__ (
    .I3(__2550__),
    .I2(__3562__),
    .I1(__3353__),
    .I0(__3462__),
    .O(__3643__)
  );
  LUT6 #(
    .INIT(64'hf8fffff8f8f8f8f8)
  ) __7327__ (
    .I5(__968__),
    .I4(__3643__),
    .I3(__3642__),
    .I2(__3638__),
    .I1(__3636__),
    .I0(__2346__),
    .O(__3644__)
  );
  LUT6 #(
    .INIT(64'h3fffff3faaaaaaaa)
  ) __7328__ (
    .I5(__2870__),
    .I4(g3229),
    .I3(__1602__),
    .I2(__1601__),
    .I1(__1600__),
    .I0(__1131__),
    .O(__3645__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7329__ (
    .I2(__2870__),
    .I1(__2617__),
    .I0(__1139__),
    .O(__3646__)
  );
  LUT4 #(
    .INIT(16'h0baa)
  ) __7330__ (
    .I3(__858__),
    .I2(__1624__),
    .I1(__2117__),
    .I0(__282__),
    .O(__3647__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __7331__ (
    .I2(__589__),
    .I1(__2510__),
    .I0(__1190__),
    .O(__3648__)
  );
  LUT6 #(
    .INIT(64'h0f005555cccccccc)
  ) __7332__ (
    .I5(__589__),
    .I4(__603__),
    .I3(__1643__),
    .I2(__1637__),
    .I1(__1184__),
    .I0(__1638__),
    .O(__3649__)
  );
  LUT5 #(
    .INIT(32'h77f0f0f0)
  ) __7333__ (
    .I4(__662__),
    .I3(__603__),
    .I2(__405__),
    .I1(__1777__),
    .I0(__1858__),
    .O(__3650__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7334__ (
    .I2(__944__),
    .I1(__2178__),
    .I0(__1376__),
    .O(__3651__)
  );
  LUT6 #(
    .INIT(64'h3fffff3faaaaaaaa)
  ) __7335__ (
    .I5(__2582__),
    .I4(g3229),
    .I3(__2070__),
    .I2(__2069__),
    .I1(__2068__),
    .I0(__628__),
    .O(__3652__)
  );
  LUT6 #(
    .INIT(64'h55555d5500000800)
  ) __7336__ (
    .I5(__1288__),
    .I4(__1430__),
    .I3(__1426__),
    .I2(__1428__),
    .I1(__1432__),
    .I0(__2407__),
    .O(__3653__)
  );
  LUT5 #(
    .INIT(32'hfcccaaaa)
  ) __7337__ (
    .I4(__954__),
    .I3(__862__),
    .I2(__868__),
    .I1(__1782__),
    .I0(__1374__),
    .O(__3654__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __7338__ (
    .I5(__944__),
    .I4(__936__),
    .I3(__927__),
    .I2(__924__),
    .I1(__893__),
    .I0(__915__),
    .O(__3655__)
  );
  LUT4 #(
    .INIT(16'haccc)
  ) __7339__ (
    .I3(__589__),
    .I2(__603__),
    .I1(__586__),
    .I0(__1705__),
    .O(__3656__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7340__ (
    .I2(__1479__),
    .I1(__1429__),
    .I0(__1472__),
    .O(__3657__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7341__ (
    .I2(__944__),
    .I1(__297__),
    .I0(__1382__),
    .O(__3658__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7342__ (
    .I2(__1479__),
    .I1(__1467__),
    .I0(__1408__),
    .O(__3659__)
  );
  LUT6 #(
    .INIT(64'hd8fad850d850d8fa)
  ) __7343__ (
    .I5(g3229),
    .I4(__2287__),
    .I3(__2286__),
    .I2(__211__),
    .I1(__2285__),
    .I0(__2370__),
    .O(__3660__)
  );
  LUT4 #(
    .INIT(16'haccc)
  ) __7344__ (
    .I3(__858__),
    .I2(__231__),
    .I1(__298__),
    .I0(__1982__),
    .O(__3661__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __7345__ (
    .I5(__944__),
    .I4(__936__),
    .I3(__927__),
    .I2(__924__),
    .I1(__902__),
    .I0(__918__),
    .O(__3662__)
  );
  LUT6 #(
    .INIT(64'hd8fad850d850d8fa)
  ) __7346__ (
    .I5(g3229),
    .I4(__2287__),
    .I3(__2286__),
    .I2(__602__),
    .I1(__2285__),
    .I0(__2288__),
    .O(__3663__)
  );
  LUT4 #(
    .INIT(16'h3aaa)
  ) __7347__ (
    .I3(__663__),
    .I2(__603__),
    .I1(__1450__),
    .I0(__827__),
    .O(__3664__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7348__ (
    .I2(__589__),
    .I1(__3062__),
    .I0(__575__),
    .O(__3665__)
  );
  LUT6 #(
    .INIT(64'hb0bb0000b0bbb0bb)
  ) __7349__ (
    .I5(__944__),
    .I4(__151__),
    .I3(__858__),
    .I2(__391__),
    .I1(__954__),
    .I0(__380__),
    .O(__3666__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7350__ (
    .I2(__1511__),
    .I1(__99__),
    .I0(__175__),
    .O(__3667__)
  );
  LUT5 #(
    .INIT(32'h4ecccccc)
  ) __7351__ (
    .I4(__589__),
    .I3(__1598__),
    .I2(__1438__),
    .I1(__778__),
    .I0(__1635__),
    .O(__3668__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7352__ (
    .I2(__1479__),
    .I1(__1461__),
    .I0(__1414__),
    .O(__3669__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7353__ (
    .I2(__662__),
    .I1(__2690__),
    .I0(__1239__),
    .O(__3670__)
  );
  LUT6 #(
    .INIT(64'h132033005fa0ff00)
  ) __7354__ (
    .I5(__954__),
    .I4(__765__),
    .I3(__772__),
    .I2(__750__),
    .I1(__752__),
    .I0(__1985__),
    .O(__3671__)
  );
  LUT5 #(
    .INIT(32'h00008000)
  ) __7355__ (
    .I4(__1598__),
    .I3(__589__),
    .I2(__656__),
    .I1(__657__),
    .I0(__658__),
    .O(__3672__)
  );
  LUT5 #(
    .INIT(32'h06666666)
  ) __7356__ (
    .I4(__589__),
    .I3(__1598__),
    .I2(__603__),
    .I1(__646__),
    .I0(__3672__),
    .O(__3673__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7357__ (
    .I2(__589__),
    .I1(__2743__),
    .I0(__613__),
    .O(__3674__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7358__ (
    .I2(__2427__),
    .I1(__3119__),
    .I0(__562__),
    .O(__3675__)
  );
  LUT5 #(
    .INIT(32'h77f0f0f0)
  ) __7359__ (
    .I4(__663__),
    .I3(__603__),
    .I2(__1075__),
    .I1(__1972__),
    .I0(__2011__),
    .O(__3676__)
  );
  LUT4 #(
    .INIT(16'haccc)
  ) __7360__ (
    .I3(__954__),
    .I2(__875__),
    .I1(__1343__),
    .I0(__2056__),
    .O(__3677__)
  );
  LUT6 #(
    .INIT(64'h132033005fa0ff00)
  ) __7361__ (
    .I5(__954__),
    .I4(__788__),
    .I3(__1055__),
    .I2(__796__),
    .I1(__875__),
    .I0(__1667__),
    .O(__3678__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7362__ (
    .I2(__662__),
    .I1(__2272__),
    .I0(__695__),
    .O(__3679__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __7363__ (
    .I5(__764__),
    .I4(__573__),
    .I3(__954__),
    .I2(__745__),
    .I1(__507__),
    .I0(__768__),
    .O(__3680__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7364__ (
    .I2(__1599__),
    .I1(__2617__),
    .I0(__1138__),
    .O(__3681__)
  );
  LUT6 #(
    .INIT(64'hc5cccccccccccccc)
  ) __7365__ (
    .I5(__944__),
    .I4(__764__),
    .I3(__573__),
    .I2(__745__),
    .I1(__682__),
    .I0(__770__),
    .O(__3682__)
  );
  assign g4590 = __1445__;
  assign g25420 = __2769__;
  assign g25442 = __2769__;
  assign g25489 = __3603__;
  assign g8021 = __1497__;
  assign g7334 = __1437__;
  assign g24734 = __68__;
  assign g8258 = __1533__;
  assign g8273 = __1514__;
  assign g5437 = __663__;
  assign g5472 = __663__;
  assign g5511 = __663__;
  assign g5555 = __663__;
  assign g6231 = __663__;
  assign g6368 = __663__;
  assign g6573 = __663__;
  assign g6837 = __663__;
  assign g7909 = __663__;
  assign g7961 = __663__;
  assign g8012 = __663__;
  assign g8087 = __663__;
  assign g8261 = __1529__;
  assign g8023 = __1427__;
  assign g26104 = __3275__;
  assign g5629 = __858__;
  assign g5657 = __858__;
  assign g5695 = __858__;
  assign g5747 = __858__;
  assign g6485 = __858__;
  assign g6677 = __858__;
  assign g6750 = __858__;
  assign g6979 = __858__;
  assign g7052 = __858__;
  assign g7229 = __858__;
  assign g7302 = __858__;
  assign g7425 = __858__;
  assign g8106 = __858__;
  assign g8096 = __1416__;
  assign g3993 = __1423__;
  assign g8259 = __1530__;
  assign g4088 = __1431__;
  assign g16355 = __94__;
  assign g8249 = __1433__;
  assign g16496 = __2584__;
  assign g16437 = __244__;
  assign g8251 = __1451__;
  assign g4090 = __1449__;
  assign g6442 = __1441__;
  assign g8266 = __1523__;
  assign g8271 = __1519__;
  assign g4323 = __1447__;
  assign g8263 = __1527__;
  assign g4321 = __1429__;
  assign g4450 = __1418__;
  assign g16297 = __937__;
  assign g8267 = __1521__;
  assign g8275 = __1512__;
  assign g4200 = __1420__;
  assign g8269 = __1517__;
  assign g7519 = __1435__;
  assign g16399 = __771__;
  assign g25435 = __69__;
  assign g5549 = __581__;
  assign g5595 = __581__;
  assign g5612 = __581__;
  assign g5637 = __581__;
  assign g8274 = __1513__;
  assign g6225 = __1443__;
  assign g8270 = __1518__;
  assign g8264 = __1525__;
  assign g8272 = __1515__;
  assign g5648 = __954__;
  assign g5686 = __954__;
  assign g5738 = __954__;
  assign g5796 = __954__;
  assign g6642 = __954__;
  assign g6911 = __954__;
  assign g6944 = __954__;
  assign g7161 = __954__;
  assign g7194 = __954__;
  assign g7357 = __954__;
  assign g7390 = __954__;
  assign g7487 = __954__;
  assign g8030 = __954__;
  assign g8268 = __1516__;
  assign g26149 = __3337__;
  assign g5388 = __1509__;
  assign g8265 = __1524__;
  assign g27380 = __70__;
  assign g6313 = __662__;
  assign g6447 = __662__;
  assign g6518 = __662__;
  assign g6712 = __662__;
  assign g6782 = __662__;
  assign g7014 = __662__;
  assign g7084 = __662__;
  assign g7264 = __662__;
  assign g7956 = __662__;
  assign g8007 = __662__;
  assign g8082 = __662__;
  assign g8167 = __662__;
  assign g26135 = __2961__;
  assign g8262 = __1526__;
  assign g8260 = __1528__;
  assign g6895 = __1439__;
  assign g8175 = __1425__;
endmodule
