module s38584 (
  CK,
  g100,
  g113,
  g114,
  g115,
  g116,
  g120,
  g124,
  g125,
  g126,
  g127,
  g134,
  g135,
  g35,
  g36,
  g44,
  g5,
  g53,
  g54,
  g56,
  g57,
  g64,
  g6744,
  g6745,
  g6746,
  g6747,
  g6748,
  g6749,
  g6750,
  g6751,
  g6752,
  g6753,
  g72,
  g73,
  g84,
  g90,
  g91,
  g92,
  g99,
  g20652,
  g29214,
  g16624,
  g17845,
  g13881,
  g33636,
  g17320,
  g14673,
  g16874,
  g28030,
  g9680,
  g12833,
  g9251,
  g28041,
  g21245,
  g29220,
  g21270,
  g29217,
  g11349,
  g13272,
  g13906,
  g17604,
  g12184,
  g18095,
  g14779,
  g8291,
  g17787,
  g13085,
  g14694,
  g23002,
  g30327,
  g20763,
  g29211,
  g14451,
  g17674,
  g12350,
  g10527,
  g25114,
  g31860,
  g34917,
  g14147,
  g34921,
  g8235,
  g18099,
  g8344,
  g18092,
  g14201,
  g34927,
  g16659,
  g9615,
  g24162,
  g16722,
  g24183,
  g14518,
  g17404,
  g24185,
  g17400,
  g34425,
  g34839,
  g34956,
  g34923,
  g17739,
  g24168,
  g7243,
  g16656,
  g16775,
  g34925,
  g24181,
  g8784,
  g24151,
  g25582,
  g25583,
  g25584,
  g25585,
  g25586,
  g25587,
  g25588,
  g25589,
  g25590,
  g32429,
  g32454,
  g33945,
  g33946,
  g33947,
  g33948,
  g33949,
  g33950,
  g34232,
  g34233,
  g34234,
  g34235,
  g34236,
  g34237,
  g34238,
  g34239,
  g34240,
  g16603,
  g17813,
  g13926,
  g17577,
  g8920,
  g21727,
  g17711,
  g17649,
  g19357,
  g7260,
  g25259,
  g31862,
  g8132,
  g27831,
  g33533,
  g8786,
  g20049,
  g29210,
  g24163,
  g24176,
  g8398,
  g24182,
  g7245,
  g24171,
  g24178,
  g12919,
  g17639,
  g11418,
  g21176,
  g29216,
  g9019,
  g8839,
  g9741,
  g16748,
  g14738,
  g26876,
  g8788,
  g16924,
  g9555,
  g33435,
  g9817,
  g17715,
  g20901,
  g29215,
  g25167,
  g31863,
  g17871,
  g23683,
  g30332,
  g24165,
  g17778,
  g24177,
  g31521,
  g34435,
  g14662,
  g32185,
  g16627,
  g9048,
  g18101,
  g14635,
  g16955,
  g16686,
  g33894,
  g34788,
  g28042,
  g8917,
  g8787,
  g14217,
  g10306,
  g10500,
  g24179,
  g17291,
  g17722,
  g9617,
  g34201,
  g13039,
  g24170,
  g20899,
  g29212,
  g13895,
  g20557,
  g29213,
  g17423,
  g9743,
  g17607,
  g13068,
  g8719,
  g17760,
  g18881,
  g29218,
  g24175,
  g8916,
  g14125,
  g26875,
  g31656,
  g34436,
  g17819,
  g13865,
  g7540,
  g21698,
  g8783,
  g12923,
  g7946,
  g18094,
  g14189,
  g21292,
  g29221,
  g18098,
  g34972,
  g11388,
  g13049,
  g18100,
  g24167,
  g8358,
  g14749,
  g11770,
  g8178,
  g14167,
  g8342,
  g8475,
  g14421,
  g8277,
  g19334,
  g34383,
  g34919,
  g17580,
  g12368,
  g28753,
  g33959,
  g33874,
  g17316,
  g8353,
  g17685,
  g16718,
  g34913,
  g10122,
  g8283,
  g33935,
  g12832,
  g12470,
  g24174,
  g33079,
  g17678,
  g20654,
  g29219,
  g14597,
  g9553,
  g24164,
  g8279,
  g8416,
  g24161,
  g24169,
  g17646,
  g18097,
  g25219,
  g31861,
  g17743,
  g33659,
  g24172,
  g31793,
  g8870,
  g12238,
  g12422,
  g8789,
  g7257,
  g17764,
  g13099,
  g34221,
  g8785,
  g16744,
  g14828,
  g24173,
  g12300,
  g14705,
  g8215,
  g11447,
  g17519,
  g8918,
  g17688,
  g31665,
  g34437,
  g24180,
  g23759,
  g30331,
  g13966,
  g26801,
  g32975,
  g24184,
  g8403,
  g23652,
  g30330,
  g11678,
  g24166,
  g26877,
  g9682,
  g7916,
  g9497,
  g13259,
  g23612,
  g30329,
  g14096,
  g34915,
  g16693,
  g8915,
  g8919,
  g23190,
  g34597,
  g18096
);
  input CK;
  wire CK;
  input g100;
  wire g100;
  input g113;
  wire g113;
  input g114;
  wire g114;
  input g115;
  wire g115;
  input g116;
  wire g116;
  input g120;
  wire g120;
  input g124;
  wire g124;
  input g125;
  wire g125;
  input g126;
  wire g126;
  input g127;
  wire g127;
  input g134;
  wire g134;
  input g135;
  wire g135;
  input g35;
  wire g35;
  input g36;
  wire g36;
  input g44;
  wire g44;
  input g5;
  wire g5;
  input g53;
  wire g53;
  input g54;
  wire g54;
  input g56;
  wire g56;
  input g57;
  wire g57;
  input g64;
  wire g64;
  input g6744;
  wire g6744;
  input g6745;
  wire g6745;
  input g6746;
  wire g6746;
  input g6747;
  wire g6747;
  input g6748;
  wire g6748;
  input g6749;
  wire g6749;
  input g6750;
  wire g6750;
  input g6751;
  wire g6751;
  input g6752;
  wire g6752;
  input g6753;
  wire g6753;
  input g72;
  wire g72;
  input g73;
  wire g73;
  input g84;
  wire g84;
  input g90;
  wire g90;
  input g91;
  wire g91;
  input g92;
  wire g92;
  input g99;
  wire g99;
  output g20652;
  wire g20652;
  output g29214;
  wire g29214;
  output g16624;
  wire g16624;
  output g17845;
  wire g17845;
  output g13881;
  wire g13881;
  output g33636;
  wire g33636;
  output g17320;
  wire g17320;
  output g14673;
  wire g14673;
  output g16874;
  wire g16874;
  output g28030;
  wire g28030;
  output g9680;
  wire g9680;
  output g12833;
  wire g12833;
  output g9251;
  wire g9251;
  output g28041;
  wire g28041;
  output g21245;
  wire g21245;
  output g29220;
  wire g29220;
  output g21270;
  wire g21270;
  output g29217;
  wire g29217;
  output g11349;
  wire g11349;
  output g13272;
  wire g13272;
  output g13906;
  wire g13906;
  output g17604;
  wire g17604;
  output g12184;
  wire g12184;
  output g18095;
  wire g18095;
  output g14779;
  wire g14779;
  output g8291;
  wire g8291;
  output g17787;
  wire g17787;
  output g13085;
  wire g13085;
  output g14694;
  wire g14694;
  output g23002;
  wire g23002;
  output g30327;
  wire g30327;
  output g20763;
  wire g20763;
  output g29211;
  wire g29211;
  output g14451;
  wire g14451;
  output g17674;
  wire g17674;
  output g12350;
  wire g12350;
  output g10527;
  wire g10527;
  output g25114;
  wire g25114;
  output g31860;
  wire g31860;
  output g34917;
  wire g34917;
  output g14147;
  wire g14147;
  output g34921;
  wire g34921;
  output g8235;
  wire g8235;
  output g18099;
  wire g18099;
  output g8344;
  wire g8344;
  output g18092;
  wire g18092;
  output g14201;
  wire g14201;
  output g34927;
  wire g34927;
  output g16659;
  wire g16659;
  output g9615;
  wire g9615;
  output g24162;
  wire g24162;
  output g16722;
  wire g16722;
  output g24183;
  wire g24183;
  output g14518;
  wire g14518;
  output g17404;
  wire g17404;
  output g24185;
  wire g24185;
  output g17400;
  wire g17400;
  output g34425;
  wire g34425;
  output g34839;
  wire g34839;
  output g34956;
  wire g34956;
  output g34923;
  wire g34923;
  output g17739;
  wire g17739;
  output g24168;
  wire g24168;
  output g7243;
  wire g7243;
  output g16656;
  wire g16656;
  output g16775;
  wire g16775;
  output g34925;
  wire g34925;
  output g24181;
  wire g24181;
  output g8784;
  wire g8784;
  output g24151;
  wire g24151;
  output g25582;
  wire g25582;
  output g25583;
  wire g25583;
  output g25584;
  wire g25584;
  output g25585;
  wire g25585;
  output g25586;
  wire g25586;
  output g25587;
  wire g25587;
  output g25588;
  wire g25588;
  output g25589;
  wire g25589;
  output g25590;
  wire g25590;
  output g32429;
  wire g32429;
  output g32454;
  wire g32454;
  output g33945;
  wire g33945;
  output g33946;
  wire g33946;
  output g33947;
  wire g33947;
  output g33948;
  wire g33948;
  output g33949;
  wire g33949;
  output g33950;
  wire g33950;
  output g34232;
  wire g34232;
  output g34233;
  wire g34233;
  output g34234;
  wire g34234;
  output g34235;
  wire g34235;
  output g34236;
  wire g34236;
  output g34237;
  wire g34237;
  output g34238;
  wire g34238;
  output g34239;
  wire g34239;
  output g34240;
  wire g34240;
  output g16603;
  wire g16603;
  output g17813;
  wire g17813;
  output g13926;
  wire g13926;
  output g17577;
  wire g17577;
  output g8920;
  wire g8920;
  output g21727;
  wire g21727;
  output g17711;
  wire g17711;
  output g17649;
  wire g17649;
  output g19357;
  wire g19357;
  output g7260;
  wire g7260;
  output g25259;
  wire g25259;
  output g31862;
  wire g31862;
  output g8132;
  wire g8132;
  output g27831;
  wire g27831;
  output g33533;
  wire g33533;
  output g8786;
  wire g8786;
  output g20049;
  wire g20049;
  output g29210;
  wire g29210;
  output g24163;
  wire g24163;
  output g24176;
  wire g24176;
  output g8398;
  wire g8398;
  output g24182;
  wire g24182;
  output g7245;
  wire g7245;
  output g24171;
  wire g24171;
  output g24178;
  wire g24178;
  output g12919;
  wire g12919;
  output g17639;
  wire g17639;
  output g11418;
  wire g11418;
  output g21176;
  wire g21176;
  output g29216;
  wire g29216;
  output g9019;
  wire g9019;
  output g8839;
  wire g8839;
  output g9741;
  wire g9741;
  output g16748;
  wire g16748;
  output g14738;
  wire g14738;
  output g26876;
  wire g26876;
  output g8788;
  wire g8788;
  output g16924;
  wire g16924;
  output g9555;
  wire g9555;
  output g33435;
  wire g33435;
  output g9817;
  wire g9817;
  output g17715;
  wire g17715;
  output g20901;
  wire g20901;
  output g29215;
  wire g29215;
  output g25167;
  wire g25167;
  output g31863;
  wire g31863;
  output g17871;
  wire g17871;
  output g23683;
  wire g23683;
  output g30332;
  wire g30332;
  output g24165;
  wire g24165;
  output g17778;
  wire g17778;
  output g24177;
  wire g24177;
  output g31521;
  wire g31521;
  output g34435;
  wire g34435;
  output g14662;
  wire g14662;
  output g32185;
  wire g32185;
  output g16627;
  wire g16627;
  output g9048;
  wire g9048;
  output g18101;
  wire g18101;
  output g14635;
  wire g14635;
  output g16955;
  wire g16955;
  output g16686;
  wire g16686;
  output g33894;
  wire g33894;
  output g34788;
  wire g34788;
  output g28042;
  wire g28042;
  output g8917;
  wire g8917;
  output g8787;
  wire g8787;
  output g14217;
  wire g14217;
  output g10306;
  wire g10306;
  output g10500;
  wire g10500;
  output g24179;
  wire g24179;
  output g17291;
  wire g17291;
  output g17722;
  wire g17722;
  output g9617;
  wire g9617;
  output g34201;
  wire g34201;
  output g13039;
  wire g13039;
  output g24170;
  wire g24170;
  output g20899;
  wire g20899;
  output g29212;
  wire g29212;
  output g13895;
  wire g13895;
  output g20557;
  wire g20557;
  output g29213;
  wire g29213;
  output g17423;
  wire g17423;
  output g9743;
  wire g9743;
  output g17607;
  wire g17607;
  output g13068;
  wire g13068;
  output g8719;
  wire g8719;
  output g17760;
  wire g17760;
  output g18881;
  wire g18881;
  output g29218;
  wire g29218;
  output g24175;
  wire g24175;
  output g8916;
  wire g8916;
  output g14125;
  wire g14125;
  output g26875;
  wire g26875;
  output g31656;
  wire g31656;
  output g34436;
  wire g34436;
  output g17819;
  wire g17819;
  output g13865;
  wire g13865;
  output g7540;
  wire g7540;
  output g21698;
  wire g21698;
  output g8783;
  wire g8783;
  output g12923;
  wire g12923;
  output g7946;
  wire g7946;
  output g18094;
  wire g18094;
  output g14189;
  wire g14189;
  output g21292;
  wire g21292;
  output g29221;
  wire g29221;
  output g18098;
  wire g18098;
  output g34972;
  wire g34972;
  output g11388;
  wire g11388;
  output g13049;
  wire g13049;
  output g18100;
  wire g18100;
  output g24167;
  wire g24167;
  output g8358;
  wire g8358;
  output g14749;
  wire g14749;
  output g11770;
  wire g11770;
  output g8178;
  wire g8178;
  output g14167;
  wire g14167;
  output g8342;
  wire g8342;
  output g8475;
  wire g8475;
  output g14421;
  wire g14421;
  output g8277;
  wire g8277;
  output g19334;
  wire g19334;
  output g34383;
  wire g34383;
  output g34919;
  wire g34919;
  output g17580;
  wire g17580;
  output g12368;
  wire g12368;
  output g28753;
  wire g28753;
  output g33959;
  wire g33959;
  output g33874;
  wire g33874;
  output g17316;
  wire g17316;
  output g8353;
  wire g8353;
  output g17685;
  wire g17685;
  output g16718;
  wire g16718;
  output g34913;
  wire g34913;
  output g10122;
  wire g10122;
  output g8283;
  wire g8283;
  output g33935;
  wire g33935;
  output g12832;
  wire g12832;
  output g12470;
  wire g12470;
  output g24174;
  wire g24174;
  output g33079;
  wire g33079;
  output g17678;
  wire g17678;
  output g20654;
  wire g20654;
  output g29219;
  wire g29219;
  output g14597;
  wire g14597;
  output g9553;
  wire g9553;
  output g24164;
  wire g24164;
  output g8279;
  wire g8279;
  output g8416;
  wire g8416;
  output g24161;
  wire g24161;
  output g24169;
  wire g24169;
  output g17646;
  wire g17646;
  output g18097;
  wire g18097;
  output g25219;
  wire g25219;
  output g31861;
  wire g31861;
  output g17743;
  wire g17743;
  output g33659;
  wire g33659;
  output g24172;
  wire g24172;
  output g31793;
  wire g31793;
  output g8870;
  wire g8870;
  output g12238;
  wire g12238;
  output g12422;
  wire g12422;
  output g8789;
  wire g8789;
  output g7257;
  wire g7257;
  output g17764;
  wire g17764;
  output g13099;
  wire g13099;
  output g34221;
  wire g34221;
  output g8785;
  wire g8785;
  output g16744;
  wire g16744;
  output g14828;
  wire g14828;
  output g24173;
  wire g24173;
  output g12300;
  wire g12300;
  output g14705;
  wire g14705;
  output g8215;
  wire g8215;
  output g11447;
  wire g11447;
  output g17519;
  wire g17519;
  output g8918;
  wire g8918;
  output g17688;
  wire g17688;
  output g31665;
  wire g31665;
  output g34437;
  wire g34437;
  output g24180;
  wire g24180;
  output g23759;
  wire g23759;
  output g30331;
  wire g30331;
  output g13966;
  wire g13966;
  output g26801;
  wire g26801;
  output g32975;
  wire g32975;
  output g24184;
  wire g24184;
  output g8403;
  wire g8403;
  output g23652;
  wire g23652;
  output g30330;
  wire g30330;
  output g11678;
  wire g11678;
  output g24166;
  wire g24166;
  output g26877;
  wire g26877;
  output g9682;
  wire g9682;
  output g7916;
  wire g7916;
  output g9497;
  wire g9497;
  output g13259;
  wire g13259;
  output g23612;
  wire g23612;
  output g30329;
  wire g30329;
  output g14096;
  wire g14096;
  output g34915;
  wire g34915;
  output g16693;
  wire g16693;
  output g8915;
  wire g8915;
  output g8919;
  wire g8919;
  output g23190;
  wire g23190;
  output g34597;
  wire g34597;
  output g18096;
  wire g18096;
  wire __0__;
  wire __1__;
  wire __2__;
  wire __3__;
  wire __4__;
  wire __5__;
  wire __6__;
  wire __7__;
  wire __8__;
  wire __9__;
  wire __10__;
  wire __11__;
  wire __12__;
  wire __13__;
  wire __14__;
  wire __15__;
  wire __16__;
  wire __17__;
  wire __18__;
  wire __19__;
  wire __20__;
  wire __21__;
  wire __22__;
  wire __23__;
  wire __24__;
  wire __25__;
  wire __26__;
  wire __27__;
  wire __28__;
  wire __29__;
  wire __30__;
  wire __31__;
  wire __32__;
  wire __33__;
  wire __34__;
  wire __35__;
  wire __36__;
  wire __37__;
  wire __38__;
  wire __39__;
  wire __40__;
  wire __41__;
  wire __42__;
  wire __43__;
  wire __44__;
  wire __45__;
  wire __46__;
  wire __47__;
  wire __48__;
  wire __49__;
  wire __50__;
  wire __51__;
  wire __52__;
  wire __53__;
  wire __54__;
  wire __55__;
  wire __56__;
  wire __57__;
  wire __58__;
  wire __59__;
  wire __60__;
  wire __61__;
  wire __62__;
  wire __63__;
  wire __64__;
  wire __65__;
  wire __66__;
  wire __67__;
  wire __68__;
  wire __69__;
  wire __70__;
  wire __71__;
  wire __72__;
  wire __73__;
  wire __74__;
  wire __75__;
  wire __76__;
  wire __77__;
  wire __78__;
  wire __79__;
  wire __80__;
  wire __81__;
  wire __82__;
  wire __83__;
  wire __84__;
  wire __85__;
  wire __86__;
  wire __87__;
  wire __88__;
  wire __89__;
  wire __90__;
  wire __91__;
  wire __92__;
  wire __93__;
  wire __94__;
  wire __95__;
  wire __96__;
  wire __97__;
  wire __98__;
  wire __99__;
  wire __100__;
  wire __101__;
  wire __102__;
  wire __103__;
  wire __104__;
  wire __105__;
  wire __106__;
  wire __107__;
  wire __108__;
  wire __109__;
  wire __110__;
  wire __111__;
  wire __112__;
  wire __113__;
  wire __114__;
  wire __115__;
  wire __116__;
  wire __117__;
  wire __118__;
  wire __119__;
  wire __120__;
  wire __121__;
  wire __122__;
  wire __123__;
  wire __124__;
  wire __125__;
  wire __126__;
  wire __127__;
  wire __128__;
  wire __129__;
  wire __130__;
  wire __131__;
  wire __132__;
  wire __133__;
  wire __134__;
  wire __135__;
  wire __136__;
  wire __137__;
  wire __138__;
  wire __139__;
  wire __140__;
  wire __141__;
  wire __142__;
  wire __143__;
  wire __144__;
  wire __145__;
  wire __146__;
  wire __147__;
  wire __148__;
  wire __149__;
  wire __150__;
  wire __151__;
  wire __152__;
  wire __153__;
  wire __154__;
  wire __155__;
  wire __156__;
  wire __157__;
  wire __158__;
  wire __159__;
  wire __160__;
  wire __161__;
  wire __162__;
  wire __163__;
  wire __164__;
  wire __165__;
  wire __166__;
  wire __167__;
  wire __168__;
  wire __169__;
  wire __170__;
  wire __171__;
  wire __172__;
  wire __173__;
  wire __174__;
  wire __175__;
  wire __176__;
  wire __177__;
  wire __178__;
  wire __179__;
  wire __180__;
  wire __181__;
  wire __182__;
  wire __183__;
  wire __184__;
  wire __185__;
  wire __186__;
  wire __187__;
  wire __188__;
  wire __189__;
  wire __190__;
  wire __191__;
  wire __192__;
  wire __193__;
  wire __194__;
  wire __195__;
  wire __196__;
  wire __197__;
  wire __198__;
  wire __199__;
  wire __200__;
  wire __201__;
  wire __202__;
  wire __203__;
  wire __204__;
  wire __205__;
  wire __206__;
  wire __207__;
  wire __208__;
  wire __209__;
  wire __210__;
  wire __211__;
  wire __212__;
  wire __213__;
  wire __214__;
  wire __215__;
  wire __216__;
  wire __217__;
  wire __218__;
  wire __219__;
  wire __220__;
  wire __221__;
  wire __222__;
  wire __223__;
  wire __224__;
  wire __225__;
  wire __226__;
  wire __227__;
  wire __228__;
  wire __229__;
  wire __230__;
  wire __231__;
  wire __232__;
  wire __233__;
  wire __234__;
  wire __235__;
  wire __236__;
  wire __237__;
  wire __238__;
  wire __239__;
  wire __240__;
  wire __241__;
  wire __242__;
  wire __243__;
  wire __244__;
  wire __245__;
  wire __246__;
  wire __247__;
  wire __248__;
  wire __249__;
  wire __250__;
  wire __251__;
  wire __252__;
  wire __253__;
  wire __254__;
  wire __255__;
  wire __256__;
  wire __257__;
  wire __258__;
  wire __259__;
  wire __260__;
  wire __261__;
  wire __262__;
  wire __263__;
  wire __264__;
  wire __265__;
  wire __266__;
  wire __267__;
  wire __268__;
  wire __269__;
  wire __270__;
  wire __271__;
  wire __272__;
  wire __273__;
  wire __274__;
  wire __275__;
  wire __276__;
  wire __277__;
  wire __278__;
  wire __279__;
  wire __280__;
  wire __281__;
  wire __282__;
  wire __283__;
  wire __284__;
  wire __285__;
  wire __286__;
  wire __287__;
  wire __288__;
  wire __289__;
  wire __290__;
  wire __291__;
  wire __292__;
  wire __293__;
  wire __294__;
  wire __295__;
  wire __296__;
  wire __297__;
  wire __298__;
  wire __299__;
  wire __300__;
  wire __301__;
  wire __302__;
  wire __303__;
  wire __304__;
  wire __305__;
  wire __306__;
  wire __307__;
  wire __308__;
  wire __309__;
  wire __310__;
  wire __311__;
  wire __312__;
  wire __313__;
  wire __314__;
  wire __315__;
  wire __316__;
  wire __317__;
  wire __318__;
  wire __319__;
  wire __320__;
  wire __321__;
  wire __322__;
  wire __323__;
  wire __324__;
  wire __325__;
  wire __326__;
  wire __327__;
  wire __328__;
  wire __329__;
  wire __330__;
  wire __331__;
  wire __332__;
  wire __333__;
  wire __334__;
  wire __335__;
  wire __336__;
  wire __337__;
  wire __338__;
  wire __339__;
  wire __340__;
  wire __341__;
  wire __342__;
  wire __343__;
  wire __344__;
  wire __345__;
  wire __346__;
  wire __347__;
  wire __348__;
  wire __349__;
  wire __350__;
  wire __351__;
  wire __352__;
  wire __353__;
  wire __354__;
  wire __355__;
  wire __356__;
  wire __357__;
  wire __358__;
  wire __359__;
  wire __360__;
  wire __361__;
  wire __362__;
  wire __363__;
  wire __364__;
  wire __365__;
  wire __366__;
  wire __367__;
  wire __368__;
  wire __369__;
  wire __370__;
  wire __371__;
  wire __372__;
  wire __373__;
  wire __374__;
  wire __375__;
  wire __376__;
  wire __377__;
  wire __378__;
  wire __379__;
  wire __380__;
  wire __381__;
  wire __382__;
  wire __383__;
  wire __384__;
  wire __385__;
  wire __386__;
  wire __387__;
  wire __388__;
  wire __389__;
  wire __390__;
  wire __391__;
  wire __392__;
  wire __393__;
  wire __394__;
  wire __395__;
  wire __396__;
  wire __397__;
  wire __398__;
  wire __399__;
  wire __400__;
  wire __401__;
  wire __402__;
  wire __403__;
  wire __404__;
  wire __405__;
  wire __406__;
  wire __407__;
  wire __408__;
  wire __409__;
  wire __410__;
  wire __411__;
  wire __412__;
  wire __413__;
  wire __414__;
  wire __415__;
  wire __416__;
  wire __417__;
  wire __418__;
  wire __419__;
  wire __420__;
  wire __421__;
  wire __422__;
  wire __423__;
  wire __424__;
  wire __425__;
  wire __426__;
  wire __427__;
  wire __428__;
  wire __429__;
  wire __430__;
  wire __431__;
  wire __432__;
  wire __433__;
  wire __434__;
  wire __435__;
  wire __436__;
  wire __437__;
  wire __438__;
  wire __439__;
  wire __440__;
  wire __441__;
  wire __442__;
  wire __443__;
  wire __444__;
  wire __445__;
  wire __446__;
  wire __447__;
  wire __448__;
  wire __449__;
  wire __450__;
  wire __451__;
  wire __452__;
  wire __453__;
  wire __454__;
  wire __455__;
  wire __456__;
  wire __457__;
  wire __458__;
  wire __459__;
  wire __460__;
  wire __461__;
  wire __462__;
  wire __463__;
  wire __464__;
  wire __465__;
  wire __466__;
  wire __467__;
  wire __468__;
  wire __469__;
  wire __470__;
  wire __471__;
  wire __472__;
  wire __473__;
  wire __474__;
  wire __475__;
  wire __476__;
  wire __477__;
  wire __478__;
  wire __479__;
  wire __480__;
  wire __481__;
  wire __482__;
  wire __483__;
  wire __484__;
  wire __485__;
  wire __486__;
  wire __487__;
  wire __488__;
  wire __489__;
  wire __490__;
  wire __491__;
  wire __492__;
  wire __493__;
  wire __494__;
  wire __495__;
  wire __496__;
  wire __497__;
  wire __498__;
  wire __499__;
  wire __500__;
  wire __501__;
  wire __502__;
  wire __503__;
  wire __504__;
  wire __505__;
  wire __506__;
  wire __507__;
  wire __508__;
  wire __509__;
  wire __510__;
  wire __511__;
  wire __512__;
  wire __513__;
  wire __514__;
  wire __515__;
  wire __516__;
  wire __517__;
  wire __518__;
  wire __519__;
  wire __520__;
  wire __521__;
  wire __522__;
  wire __523__;
  wire __524__;
  wire __525__;
  wire __526__;
  wire __527__;
  wire __528__;
  wire __529__;
  wire __530__;
  wire __531__;
  wire __532__;
  wire __533__;
  wire __534__;
  wire __535__;
  wire __536__;
  wire __537__;
  wire __538__;
  wire __539__;
  wire __540__;
  wire __541__;
  wire __542__;
  wire __543__;
  wire __544__;
  wire __545__;
  wire __546__;
  wire __547__;
  wire __548__;
  wire __549__;
  wire __550__;
  wire __551__;
  wire __552__;
  wire __553__;
  wire __554__;
  wire __555__;
  wire __556__;
  wire __557__;
  wire __558__;
  wire __559__;
  wire __560__;
  wire __561__;
  wire __562__;
  wire __563__;
  wire __564__;
  wire __565__;
  wire __566__;
  wire __567__;
  wire __568__;
  wire __569__;
  wire __570__;
  wire __571__;
  wire __572__;
  wire __573__;
  wire __574__;
  wire __575__;
  wire __576__;
  wire __577__;
  wire __578__;
  wire __579__;
  wire __580__;
  wire __581__;
  wire __582__;
  wire __583__;
  wire __584__;
  wire __585__;
  wire __586__;
  wire __587__;
  wire __588__;
  wire __589__;
  wire __590__;
  wire __591__;
  wire __592__;
  wire __593__;
  wire __594__;
  wire __595__;
  wire __596__;
  wire __597__;
  wire __598__;
  wire __599__;
  wire __600__;
  wire __601__;
  wire __602__;
  wire __603__;
  wire __604__;
  wire __605__;
  wire __606__;
  wire __607__;
  wire __608__;
  wire __609__;
  wire __610__;
  wire __611__;
  wire __612__;
  wire __613__;
  wire __614__;
  wire __615__;
  wire __616__;
  wire __617__;
  wire __618__;
  wire __619__;
  wire __620__;
  wire __621__;
  wire __622__;
  wire __623__;
  wire __624__;
  wire __625__;
  wire __626__;
  wire __627__;
  wire __628__;
  wire __629__;
  wire __630__;
  wire __631__;
  wire __632__;
  wire __633__;
  wire __634__;
  wire __635__;
  wire __636__;
  wire __637__;
  wire __638__;
  wire __639__;
  wire __640__;
  wire __641__;
  wire __642__;
  wire __643__;
  wire __644__;
  wire __645__;
  wire __646__;
  wire __647__;
  wire __648__;
  wire __649__;
  wire __650__;
  wire __651__;
  wire __652__;
  wire __653__;
  wire __654__;
  wire __655__;
  wire __656__;
  wire __657__;
  wire __658__;
  wire __659__;
  wire __660__;
  wire __661__;
  wire __662__;
  wire __663__;
  wire __664__;
  wire __665__;
  wire __666__;
  wire __667__;
  wire __668__;
  wire __669__;
  wire __670__;
  wire __671__;
  wire __672__;
  wire __673__;
  wire __674__;
  wire __675__;
  wire __676__;
  wire __677__;
  wire __678__;
  wire __679__;
  wire __680__;
  wire __681__;
  wire __682__;
  wire __683__;
  wire __684__;
  wire __685__;
  wire __686__;
  wire __687__;
  wire __688__;
  wire __689__;
  wire __690__;
  wire __691__;
  wire __692__;
  wire __693__;
  wire __694__;
  wire __695__;
  wire __696__;
  wire __697__;
  wire __698__;
  wire __699__;
  wire __700__;
  wire __701__;
  wire __702__;
  wire __703__;
  wire __704__;
  wire __705__;
  wire __706__;
  wire __707__;
  wire __708__;
  wire __709__;
  wire __710__;
  wire __711__;
  wire __712__;
  wire __713__;
  wire __714__;
  wire __715__;
  wire __716__;
  wire __717__;
  wire __718__;
  wire __719__;
  wire __720__;
  wire __721__;
  wire __722__;
  wire __723__;
  wire __724__;
  wire __725__;
  wire __726__;
  wire __727__;
  wire __728__;
  wire __729__;
  wire __730__;
  wire __731__;
  wire __732__;
  wire __733__;
  wire __734__;
  wire __735__;
  wire __736__;
  wire __737__;
  wire __738__;
  wire __739__;
  wire __740__;
  wire __741__;
  wire __742__;
  wire __743__;
  wire __744__;
  wire __745__;
  wire __746__;
  wire __747__;
  wire __748__;
  wire __749__;
  wire __750__;
  wire __751__;
  wire __752__;
  wire __753__;
  wire __754__;
  wire __755__;
  wire __756__;
  wire __757__;
  wire __758__;
  wire __759__;
  wire __760__;
  wire __761__;
  wire __762__;
  wire __763__;
  wire __764__;
  wire __765__;
  wire __766__;
  wire __767__;
  wire __768__;
  wire __769__;
  wire __770__;
  wire __771__;
  wire __772__;
  wire __773__;
  wire __774__;
  wire __775__;
  wire __776__;
  wire __777__;
  wire __778__;
  wire __779__;
  wire __780__;
  wire __781__;
  wire __782__;
  wire __783__;
  wire __784__;
  wire __785__;
  wire __786__;
  wire __787__;
  wire __788__;
  wire __789__;
  wire __790__;
  wire __791__;
  wire __792__;
  wire __793__;
  wire __794__;
  wire __795__;
  wire __796__;
  wire __797__;
  wire __798__;
  wire __799__;
  wire __800__;
  wire __801__;
  wire __802__;
  wire __803__;
  wire __804__;
  wire __805__;
  wire __806__;
  wire __807__;
  wire __808__;
  wire __809__;
  wire __810__;
  wire __811__;
  wire __812__;
  wire __813__;
  wire __814__;
  wire __815__;
  wire __816__;
  wire __817__;
  wire __818__;
  wire __819__;
  wire __820__;
  wire __821__;
  wire __822__;
  wire __823__;
  wire __824__;
  wire __825__;
  wire __826__;
  wire __827__;
  wire __828__;
  wire __829__;
  wire __830__;
  wire __831__;
  wire __832__;
  wire __833__;
  wire __834__;
  wire __835__;
  wire __836__;
  wire __837__;
  wire __838__;
  wire __839__;
  wire __840__;
  wire __841__;
  wire __842__;
  wire __843__;
  wire __844__;
  wire __845__;
  wire __846__;
  wire __847__;
  wire __848__;
  wire __849__;
  wire __850__;
  wire __851__;
  wire __852__;
  wire __853__;
  wire __854__;
  wire __855__;
  wire __856__;
  wire __857__;
  wire __858__;
  wire __859__;
  wire __860__;
  wire __861__;
  wire __862__;
  wire __863__;
  wire __864__;
  wire __865__;
  wire __866__;
  wire __867__;
  wire __868__;
  wire __869__;
  wire __870__;
  wire __871__;
  wire __872__;
  wire __873__;
  wire __874__;
  wire __875__;
  wire __876__;
  wire __877__;
  wire __878__;
  wire __879__;
  wire __880__;
  wire __881__;
  wire __882__;
  wire __883__;
  wire __884__;
  wire __885__;
  wire __886__;
  wire __887__;
  wire __888__;
  wire __889__;
  wire __890__;
  wire __891__;
  wire __892__;
  wire __893__;
  wire __894__;
  wire __895__;
  wire __896__;
  wire __897__;
  wire __898__;
  wire __899__;
  wire __900__;
  wire __901__;
  wire __902__;
  wire __903__;
  wire __904__;
  wire __905__;
  wire __906__;
  wire __907__;
  wire __908__;
  wire __909__;
  wire __910__;
  wire __911__;
  wire __912__;
  wire __913__;
  wire __914__;
  wire __915__;
  wire __916__;
  wire __917__;
  wire __918__;
  wire __919__;
  wire __920__;
  wire __921__;
  wire __922__;
  wire __923__;
  wire __924__;
  wire __925__;
  wire __926__;
  wire __927__;
  wire __928__;
  wire __929__;
  wire __930__;
  wire __931__;
  wire __932__;
  wire __933__;
  wire __934__;
  wire __935__;
  wire __936__;
  wire __937__;
  wire __938__;
  wire __939__;
  wire __940__;
  wire __941__;
  wire __942__;
  wire __943__;
  wire __944__;
  wire __945__;
  wire __946__;
  wire __947__;
  wire __948__;
  wire __949__;
  wire __950__;
  wire __951__;
  wire __952__;
  wire __953__;
  wire __954__;
  wire __955__;
  wire __956__;
  wire __957__;
  wire __958__;
  wire __959__;
  wire __960__;
  wire __961__;
  wire __962__;
  wire __963__;
  wire __964__;
  wire __965__;
  wire __966__;
  wire __967__;
  wire __968__;
  wire __969__;
  wire __970__;
  wire __971__;
  wire __972__;
  wire __973__;
  wire __974__;
  wire __975__;
  wire __976__;
  wire __977__;
  wire __978__;
  wire __979__;
  wire __980__;
  wire __981__;
  wire __982__;
  wire __983__;
  wire __984__;
  wire __985__;
  wire __986__;
  wire __987__;
  wire __988__;
  wire __989__;
  wire __990__;
  wire __991__;
  wire __992__;
  wire __993__;
  wire __994__;
  wire __995__;
  wire __996__;
  wire __997__;
  wire __998__;
  wire __999__;
  wire __1000__;
  wire __1001__;
  wire __1002__;
  wire __1003__;
  wire __1004__;
  wire __1005__;
  wire __1006__;
  wire __1007__;
  wire __1008__;
  wire __1009__;
  wire __1010__;
  wire __1011__;
  wire __1012__;
  wire __1013__;
  wire __1014__;
  wire __1015__;
  wire __1016__;
  wire __1017__;
  wire __1018__;
  wire __1019__;
  wire __1020__;
  wire __1021__;
  wire __1022__;
  wire __1023__;
  wire __1024__;
  wire __1025__;
  wire __1026__;
  wire __1027__;
  wire __1028__;
  wire __1029__;
  wire __1030__;
  wire __1031__;
  wire __1032__;
  wire __1033__;
  wire __1034__;
  wire __1035__;
  wire __1036__;
  wire __1037__;
  wire __1038__;
  wire __1039__;
  wire __1040__;
  wire __1041__;
  wire __1042__;
  wire __1043__;
  wire __1044__;
  wire __1045__;
  wire __1046__;
  wire __1047__;
  wire __1048__;
  wire __1049__;
  wire __1050__;
  wire __1051__;
  wire __1052__;
  wire __1053__;
  wire __1054__;
  wire __1055__;
  wire __1056__;
  wire __1057__;
  wire __1058__;
  wire __1059__;
  wire __1060__;
  wire __1061__;
  wire __1062__;
  wire __1063__;
  wire __1064__;
  wire __1065__;
  wire __1066__;
  wire __1067__;
  wire __1068__;
  wire __1069__;
  wire __1070__;
  wire __1071__;
  wire __1072__;
  wire __1073__;
  wire __1074__;
  wire __1075__;
  wire __1076__;
  wire __1077__;
  wire __1078__;
  wire __1079__;
  wire __1080__;
  wire __1081__;
  wire __1082__;
  wire __1083__;
  wire __1084__;
  wire __1085__;
  wire __1086__;
  wire __1087__;
  wire __1088__;
  wire __1089__;
  wire __1090__;
  wire __1091__;
  wire __1092__;
  wire __1093__;
  wire __1094__;
  wire __1095__;
  wire __1096__;
  wire __1097__;
  wire __1098__;
  wire __1099__;
  wire __1100__;
  wire __1101__;
  wire __1102__;
  wire __1103__;
  wire __1104__;
  wire __1105__;
  wire __1106__;
  wire __1107__;
  wire __1108__;
  wire __1109__;
  wire __1110__;
  wire __1111__;
  wire __1112__;
  wire __1113__;
  wire __1114__;
  wire __1115__;
  wire __1116__;
  wire __1117__;
  wire __1118__;
  wire __1119__;
  wire __1120__;
  wire __1121__;
  wire __1122__;
  wire __1123__;
  wire __1124__;
  wire __1125__;
  wire __1126__;
  wire __1127__;
  wire __1128__;
  wire __1129__;
  wire __1130__;
  wire __1131__;
  wire __1132__;
  wire __1133__;
  wire __1134__;
  wire __1135__;
  wire __1136__;
  wire __1137__;
  wire __1138__;
  wire __1139__;
  wire __1140__;
  wire __1141__;
  wire __1142__;
  wire __1143__;
  wire __1144__;
  wire __1145__;
  wire __1146__;
  wire __1147__;
  wire __1148__;
  wire __1149__;
  wire __1150__;
  wire __1151__;
  wire __1152__;
  wire __1153__;
  wire __1154__;
  wire __1155__;
  wire __1156__;
  wire __1157__;
  wire __1158__;
  wire __1159__;
  wire __1160__;
  wire __1161__;
  wire __1162__;
  wire __1163__;
  wire __1164__;
  wire __1165__;
  wire __1166__;
  wire __1167__;
  wire __1168__;
  wire __1169__;
  wire __1170__;
  wire __1171__;
  wire __1172__;
  wire __1173__;
  wire __1174__;
  wire __1175__;
  wire __1176__;
  wire __1177__;
  wire __1178__;
  wire __1179__;
  wire __1180__;
  wire __1181__;
  wire __1182__;
  wire __1183__;
  wire __1184__;
  wire __1185__;
  wire __1186__;
  wire __1187__;
  wire __1188__;
  wire __1189__;
  wire __1190__;
  wire __1191__;
  wire __1192__;
  wire __1193__;
  wire __1194__;
  wire __1195__;
  wire __1196__;
  wire __1197__;
  wire __1198__;
  wire __1199__;
  wire __1200__;
  wire __1201__;
  wire __1202__;
  wire __1203__;
  wire __1204__;
  wire __1205__;
  wire __1206__;
  wire __1207__;
  wire __1208__;
  wire __1209__;
  wire __1210__;
  wire __1211__;
  wire __1212__;
  wire __1213__;
  wire __1214__;
  wire __1215__;
  wire __1216__;
  wire __1217__;
  wire __1218__;
  wire __1219__;
  wire __1220__;
  wire __1221__;
  wire __1222__;
  wire __1223__;
  wire __1224__;
  wire __1225__;
  wire __1226__;
  wire __1227__;
  wire __1228__;
  wire __1229__;
  wire __1230__;
  wire __1231__;
  wire __1232__;
  wire __1233__;
  wire __1234__;
  wire __1235__;
  wire __1236__;
  wire __1237__;
  wire __1238__;
  wire __1239__;
  wire __1240__;
  wire __1241__;
  wire __1242__;
  wire __1243__;
  wire __1244__;
  wire __1245__;
  wire __1246__;
  wire __1247__;
  wire __1248__;
  wire __1249__;
  wire __1250__;
  wire __1251__;
  wire __1252__;
  wire __1253__;
  wire __1254__;
  wire __1255__;
  wire __1256__;
  wire __1257__;
  wire __1258__;
  wire __1259__;
  wire __1260__;
  wire __1261__;
  wire __1262__;
  wire __1263__;
  wire __1264__;
  wire __1265__;
  wire __1266__;
  wire __1267__;
  wire __1268__;
  wire __1269__;
  wire __1270__;
  wire __1271__;
  wire __1272__;
  wire __1273__;
  wire __1274__;
  wire __1275__;
  wire __1276__;
  wire __1277__;
  wire __1278__;
  wire __1279__;
  wire __1280__;
  wire __1282__;
  wire __1283__;
  wire __1284__;
  wire __1285__;
  wire __1286__;
  wire __1287__;
  wire __1289__;
  wire __1290__;
  wire __1291__;
  wire __1292__;
  wire __1293__;
  wire __1294__;
  wire __1295__;
  wire __1296__;
  wire __1297__;
  wire __1298__;
  wire __1299__;
  wire __1300__;
  wire __1301__;
  wire __1302__;
  wire __1303__;
  wire __1304__;
  wire __1305__;
  wire __1306__;
  wire __1307__;
  wire __1308__;
  wire __1309__;
  wire __1310__;
  wire __1311__;
  wire __1312__;
  wire __1313__;
  wire __1314__;
  wire __1315__;
  wire __1316__;
  wire __1317__;
  wire __1318__;
  wire __1319__;
  wire __1320__;
  wire __1321__;
  wire __1322__;
  wire __1323__;
  wire __1324__;
  wire __1325__;
  wire __1326__;
  wire __1327__;
  wire __1328__;
  wire __1329__;
  wire __1330__;
  wire __1331__;
  wire __1332__;
  wire __1333__;
  wire __1334__;
  wire __1335__;
  wire __1336__;
  wire __1337__;
  wire __1338__;
  wire __1339__;
  wire __1340__;
  wire __1341__;
  wire __1342__;
  wire __1343__;
  wire __1344__;
  wire __1345__;
  wire __1346__;
  wire __1347__;
  wire __1348__;
  wire __1349__;
  wire __1350__;
  wire __1351__;
  wire __1352__;
  wire __1353__;
  wire __1354__;
  wire __1355__;
  wire __1356__;
  wire __1357__;
  wire __1358__;
  wire __1359__;
  wire __1360__;
  wire __1361__;
  wire __1362__;
  wire __1363__;
  wire __1364__;
  wire __1365__;
  wire __1366__;
  wire __1367__;
  wire __1368__;
  wire __1369__;
  wire __1370__;
  wire __1371__;
  wire __1372__;
  wire __1373__;
  wire __1374__;
  wire __1375__;
  wire __1376__;
  wire __1377__;
  wire __1378__;
  wire __1379__;
  wire __1380__;
  wire __1381__;
  wire __1382__;
  wire __1383__;
  wire __1384__;
  wire __1385__;
  wire __1386__;
  wire __1387__;
  wire __1388__;
  wire __1389__;
  wire __1390__;
  wire __1391__;
  wire __1392__;
  wire __1393__;
  wire __1394__;
  wire __1395__;
  wire __1396__;
  wire __1397__;
  wire __1398__;
  wire __1399__;
  wire __1400__;
  wire __1401__;
  wire __1402__;
  wire __1403__;
  wire __1404__;
  wire __1405__;
  wire __1406__;
  wire __1407__;
  wire __1408__;
  wire __1409__;
  wire __1410__;
  wire __1411__;
  wire __1412__;
  wire __1413__;
  wire __1414__;
  wire __1415__;
  wire __1416__;
  wire __1417__;
  wire __1418__;
  wire __1419__;
  wire __1420__;
  wire __1421__;
  wire __1422__;
  wire __1423__;
  wire __1424__;
  wire __1425__;
  wire __1426__;
  wire __1427__;
  wire __1428__;
  wire __1429__;
  wire __1430__;
  wire __1431__;
  wire __1432__;
  wire __1433__;
  wire __1434__;
  wire __1435__;
  wire __1436__;
  wire __1437__;
  wire __1438__;
  wire __1439__;
  wire __1440__;
  wire __1441__;
  wire __1442__;
  wire __1443__;
  wire __1444__;
  wire __1445__;
  wire __1446__;
  wire __1447__;
  wire __1448__;
  wire __1449__;
  wire __1450__;
  wire __1451__;
  wire __1452__;
  wire __1453__;
  wire __1454__;
  wire __1455__;
  wire __1456__;
  wire __1457__;
  wire __1458__;
  wire __1459__;
  wire __1460__;
  wire __1461__;
  wire __1462__;
  wire __1463__;
  wire __1464__;
  wire __1465__;
  wire __1466__;
  wire __1467__;
  wire __1468__;
  wire __1469__;
  wire __1470__;
  wire __1471__;
  wire __1472__;
  wire __1473__;
  wire __1474__;
  wire __1475__;
  wire __1476__;
  wire __1477__;
  wire __1478__;
  wire __1479__;
  wire __1480__;
  wire __1481__;
  wire __1482__;
  wire __1483__;
  wire __1484__;
  wire __1485__;
  wire __1486__;
  wire __1487__;
  wire __1488__;
  wire __1489__;
  wire __1490__;
  wire __1491__;
  wire __1492__;
  wire __1493__;
  wire __1494__;
  wire __1495__;
  wire __1496__;
  wire __1497__;
  wire __1498__;
  wire __1499__;
  wire __1500__;
  wire __1501__;
  wire __1502__;
  wire __1503__;
  wire __1504__;
  wire __1505__;
  wire __1506__;
  wire __1507__;
  wire __1508__;
  wire __1509__;
  wire __1510__;
  wire __1511__;
  wire __1512__;
  wire __1513__;
  wire __1514__;
  wire __1515__;
  wire __1516__;
  wire __1517__;
  wire __1518__;
  wire __1519__;
  wire __1520__;
  wire __1521__;
  wire __1522__;
  wire __1523__;
  wire __1524__;
  wire __1525__;
  wire __1526__;
  wire __1527__;
  wire __1528__;
  wire __1529__;
  wire __1530__;
  wire __1531__;
  wire __1532__;
  wire __1533__;
  wire __1534__;
  wire __1535__;
  wire __1536__;
  wire __1537__;
  wire __1538__;
  wire __1539__;
  wire __1540__;
  wire __1541__;
  wire __1542__;
  wire __1543__;
  wire __1544__;
  wire __1545__;
  wire __1546__;
  wire __1547__;
  wire __1548__;
  wire __1549__;
  wire __1550__;
  wire __1551__;
  wire __1552__;
  wire __1553__;
  wire __1554__;
  wire __1555__;
  wire __1556__;
  wire __1557__;
  wire __1558__;
  wire __1559__;
  wire __1560__;
  wire __1561__;
  wire __1562__;
  wire __1563__;
  wire __1564__;
  wire __1565__;
  wire __1566__;
  wire __1567__;
  wire __1568__;
  wire __1569__;
  wire __1570__;
  wire __1571__;
  wire __1572__;
  wire __1573__;
  wire __1574__;
  wire __1575__;
  wire __1576__;
  wire __1577__;
  wire __1578__;
  wire __1579__;
  wire __1580__;
  wire __1581__;
  wire __1582__;
  wire __1583__;
  wire __1584__;
  wire __1585__;
  wire __1586__;
  wire __1587__;
  wire __1588__;
  wire __1589__;
  wire __1590__;
  wire __1591__;
  wire __1592__;
  wire __1593__;
  wire __1594__;
  wire __1595__;
  wire __1596__;
  wire __1597__;
  wire __1598__;
  wire __1599__;
  wire __1600__;
  wire __1601__;
  wire __1602__;
  wire __1603__;
  wire __1604__;
  wire __1605__;
  wire __1606__;
  wire __1607__;
  wire __1608__;
  wire __1609__;
  wire __1610__;
  wire __1611__;
  wire __1612__;
  wire __1613__;
  wire __1614__;
  wire __1615__;
  wire __1616__;
  wire __1617__;
  wire __1618__;
  wire __1619__;
  wire __1620__;
  wire __1621__;
  wire __1622__;
  wire __1623__;
  wire __1624__;
  wire __1625__;
  wire __1626__;
  wire __1627__;
  wire __1628__;
  wire __1629__;
  wire __1630__;
  wire __1631__;
  wire __1632__;
  wire __1633__;
  wire __1634__;
  wire __1635__;
  wire __1636__;
  wire __1637__;
  wire __1638__;
  wire __1639__;
  wire __1640__;
  wire __1641__;
  wire __1642__;
  wire __1643__;
  wire __1644__;
  wire __1645__;
  wire __1646__;
  wire __1647__;
  wire __1648__;
  wire __1649__;
  wire __1650__;
  wire __1651__;
  wire __1652__;
  wire __1653__;
  wire __1654__;
  wire __1655__;
  wire __1656__;
  wire __1657__;
  wire __1658__;
  wire __1659__;
  wire __1660__;
  wire __1661__;
  wire __1662__;
  wire __1663__;
  wire __1664__;
  wire __1665__;
  wire __1666__;
  wire __1667__;
  wire __1668__;
  wire __1669__;
  wire __1670__;
  wire __1671__;
  wire __1672__;
  wire __1673__;
  wire __1674__;
  wire __1675__;
  wire __1676__;
  wire __1677__;
  wire __1678__;
  wire __1679__;
  wire __1680__;
  wire __1681__;
  wire __1682__;
  wire __1683__;
  wire __1684__;
  wire __1685__;
  wire __1686__;
  wire __1687__;
  wire __1688__;
  wire __1689__;
  wire __1690__;
  wire __1691__;
  wire __1692__;
  wire __1693__;
  wire __1694__;
  wire __1695__;
  wire __1696__;
  wire __1697__;
  wire __1698__;
  wire __1699__;
  wire __1700__;
  wire __1701__;
  wire __1702__;
  wire __1703__;
  wire __1704__;
  wire __1705__;
  wire __1706__;
  wire __1707__;
  wire __1708__;
  wire __1709__;
  wire __1710__;
  wire __1711__;
  wire __1712__;
  wire __1713__;
  wire __1714__;
  wire __1715__;
  wire __1716__;
  wire __1717__;
  wire __1718__;
  wire __1719__;
  wire __1720__;
  wire __1721__;
  wire __1722__;
  wire __1723__;
  wire __1724__;
  wire __1725__;
  wire __1726__;
  wire __1727__;
  wire __1728__;
  wire __1729__;
  wire __1730__;
  wire __1731__;
  wire __1732__;
  wire __1733__;
  wire __1734__;
  wire __1735__;
  wire __1736__;
  wire __1737__;
  wire __1738__;
  wire __1739__;
  wire __1740__;
  wire __1741__;
  wire __1742__;
  wire __1743__;
  wire __1744__;
  wire __1745__;
  wire __1746__;
  wire __1747__;
  wire __1748__;
  wire __1749__;
  wire __1750__;
  wire __1751__;
  wire __1752__;
  wire __1753__;
  wire __1754__;
  wire __1755__;
  wire __1756__;
  wire __1757__;
  wire __1758__;
  wire __1759__;
  wire __1760__;
  wire __1761__;
  wire __1762__;
  wire __1763__;
  wire __1764__;
  wire __1765__;
  wire __1766__;
  wire __1767__;
  wire __1768__;
  wire __1769__;
  wire __1770__;
  wire __1771__;
  wire __1772__;
  wire __1773__;
  wire __1774__;
  wire __1775__;
  wire __1776__;
  wire __1777__;
  wire __1778__;
  wire __1779__;
  wire __1780__;
  wire __1781__;
  wire __1782__;
  wire __1783__;
  wire __1784__;
  wire __1785__;
  wire __1786__;
  wire __1787__;
  wire __1788__;
  wire __1789__;
  wire __1790__;
  wire __1791__;
  wire __1792__;
  wire __1793__;
  wire __1794__;
  wire __1795__;
  wire __1796__;
  wire __1797__;
  wire __1798__;
  wire __1799__;
  wire __1800__;
  wire __1801__;
  wire __1802__;
  wire __1803__;
  wire __1804__;
  wire __1805__;
  wire __1806__;
  wire __1807__;
  wire __1808__;
  wire __1809__;
  wire __1810__;
  wire __1811__;
  wire __1812__;
  wire __1813__;
  wire __1814__;
  wire __1815__;
  wire __1816__;
  wire __1817__;
  wire __1818__;
  wire __1819__;
  wire __1820__;
  wire __1821__;
  wire __1822__;
  wire __1823__;
  wire __1824__;
  wire __1825__;
  wire __1826__;
  wire __1827__;
  wire __1828__;
  wire __1829__;
  wire __1830__;
  wire __1831__;
  wire __1832__;
  wire __1833__;
  wire __1834__;
  wire __1835__;
  wire __1836__;
  wire __1837__;
  wire __1838__;
  wire __1839__;
  wire __1840__;
  wire __1841__;
  wire __1842__;
  wire __1843__;
  wire __1844__;
  wire __1845__;
  wire __1846__;
  wire __1847__;
  wire __1848__;
  wire __1849__;
  wire __1850__;
  wire __1851__;
  wire __1852__;
  wire __1853__;
  wire __1854__;
  wire __1855__;
  wire __1856__;
  wire __1857__;
  wire __1858__;
  wire __1859__;
  wire __1860__;
  wire __1861__;
  wire __1862__;
  wire __1863__;
  wire __1864__;
  wire __1865__;
  wire __1866__;
  wire __1867__;
  wire __1868__;
  wire __1869__;
  wire __1870__;
  wire __1871__;
  wire __1872__;
  wire __1873__;
  wire __1874__;
  wire __1875__;
  wire __1876__;
  wire __1877__;
  wire __1878__;
  wire __1879__;
  wire __1880__;
  wire __1881__;
  wire __1882__;
  wire __1883__;
  wire __1884__;
  wire __1885__;
  wire __1886__;
  wire __1887__;
  wire __1888__;
  wire __1889__;
  wire __1890__;
  wire __1891__;
  wire __1892__;
  wire __1893__;
  wire __1894__;
  wire __1895__;
  wire __1896__;
  wire __1897__;
  wire __1898__;
  wire __1899__;
  wire __1900__;
  wire __1901__;
  wire __1902__;
  wire __1903__;
  wire __1904__;
  wire __1905__;
  wire __1906__;
  wire __1907__;
  wire __1908__;
  wire __1909__;
  wire __1910__;
  wire __1911__;
  wire __1912__;
  wire __1913__;
  wire __1914__;
  wire __1915__;
  wire __1916__;
  wire __1917__;
  wire __1918__;
  wire __1919__;
  wire __1920__;
  wire __1921__;
  wire __1922__;
  wire __1923__;
  wire __1924__;
  wire __1925__;
  wire __1926__;
  wire __1927__;
  wire __1928__;
  wire __1929__;
  wire __1930__;
  wire __1931__;
  wire __1932__;
  wire __1933__;
  wire __1934__;
  wire __1935__;
  wire __1936__;
  wire __1937__;
  wire __1938__;
  wire __1939__;
  wire __1940__;
  wire __1941__;
  wire __1942__;
  wire __1943__;
  wire __1944__;
  wire __1945__;
  wire __1946__;
  wire __1947__;
  wire __1948__;
  wire __1949__;
  wire __1950__;
  wire __1951__;
  wire __1952__;
  wire __1953__;
  wire __1954__;
  wire __1955__;
  wire __1956__;
  wire __1957__;
  wire __1958__;
  wire __1959__;
  wire __1960__;
  wire __1961__;
  wire __1962__;
  wire __1963__;
  wire __1964__;
  wire __1965__;
  wire __1966__;
  wire __1967__;
  wire __1968__;
  wire __1969__;
  wire __1970__;
  wire __1971__;
  wire __1972__;
  wire __1973__;
  wire __1974__;
  wire __1975__;
  wire __1976__;
  wire __1977__;
  wire __1978__;
  wire __1979__;
  wire __1980__;
  wire __1981__;
  wire __1982__;
  wire __1983__;
  wire __1984__;
  wire __1985__;
  wire __1986__;
  wire __1987__;
  wire __1988__;
  wire __1989__;
  wire __1990__;
  wire __1991__;
  wire __1992__;
  wire __1993__;
  wire __1994__;
  wire __1995__;
  wire __1996__;
  wire __1997__;
  wire __1998__;
  wire __1999__;
  wire __2000__;
  wire __2001__;
  wire __2002__;
  wire __2003__;
  wire __2004__;
  wire __2005__;
  wire __2006__;
  wire __2007__;
  wire __2008__;
  wire __2009__;
  wire __2010__;
  wire __2011__;
  wire __2012__;
  wire __2013__;
  wire __2014__;
  wire __2015__;
  wire __2016__;
  wire __2017__;
  wire __2018__;
  wire __2019__;
  wire __2020__;
  wire __2021__;
  wire __2022__;
  wire __2023__;
  wire __2024__;
  wire __2025__;
  wire __2026__;
  wire __2027__;
  wire __2028__;
  wire __2029__;
  wire __2030__;
  wire __2031__;
  wire __2032__;
  wire __2033__;
  wire __2034__;
  wire __2035__;
  wire __2036__;
  wire __2037__;
  wire __2038__;
  wire __2039__;
  wire __2040__;
  wire __2041__;
  wire __2042__;
  wire __2043__;
  wire __2044__;
  wire __2045__;
  wire __2046__;
  wire __2047__;
  wire __2048__;
  wire __2049__;
  wire __2050__;
  wire __2051__;
  wire __2052__;
  wire __2053__;
  wire __2054__;
  wire __2055__;
  wire __2056__;
  wire __2057__;
  wire __2058__;
  wire __2059__;
  wire __2060__;
  wire __2061__;
  wire __2062__;
  wire __2063__;
  wire __2064__;
  wire __2065__;
  wire __2066__;
  wire __2067__;
  wire __2068__;
  wire __2069__;
  wire __2070__;
  wire __2071__;
  wire __2072__;
  wire __2073__;
  wire __2074__;
  wire __2075__;
  wire __2076__;
  wire __2077__;
  wire __2078__;
  wire __2079__;
  wire __2080__;
  wire __2081__;
  wire __2082__;
  wire __2083__;
  wire __2084__;
  wire __2085__;
  wire __2086__;
  wire __2087__;
  wire __2088__;
  wire __2089__;
  wire __2090__;
  wire __2091__;
  wire __2092__;
  wire __2093__;
  wire __2094__;
  wire __2095__;
  wire __2096__;
  wire __2097__;
  wire __2098__;
  wire __2099__;
  wire __2100__;
  wire __2101__;
  wire __2102__;
  wire __2103__;
  wire __2104__;
  wire __2105__;
  wire __2106__;
  wire __2107__;
  wire __2108__;
  wire __2109__;
  wire __2110__;
  wire __2111__;
  wire __2112__;
  wire __2113__;
  wire __2114__;
  wire __2115__;
  wire __2116__;
  wire __2117__;
  wire __2118__;
  wire __2119__;
  wire __2120__;
  wire __2121__;
  wire __2122__;
  wire __2123__;
  wire __2124__;
  wire __2125__;
  wire __2126__;
  wire __2127__;
  wire __2128__;
  wire __2129__;
  wire __2130__;
  wire __2131__;
  wire __2132__;
  wire __2133__;
  wire __2134__;
  wire __2135__;
  wire __2136__;
  wire __2137__;
  wire __2138__;
  wire __2139__;
  wire __2140__;
  wire __2141__;
  wire __2142__;
  wire __2143__;
  wire __2144__;
  wire __2145__;
  wire __2146__;
  wire __2147__;
  wire __2148__;
  wire __2149__;
  wire __2150__;
  wire __2151__;
  wire __2152__;
  wire __2153__;
  wire __2154__;
  wire __2155__;
  wire __2156__;
  wire __2157__;
  wire __2158__;
  wire __2159__;
  wire __2160__;
  wire __2161__;
  wire __2162__;
  wire __2163__;
  wire __2164__;
  wire __2165__;
  wire __2166__;
  wire __2167__;
  wire __2168__;
  wire __2169__;
  wire __2170__;
  wire __2171__;
  wire __2172__;
  wire __2173__;
  wire __2174__;
  wire __2175__;
  wire __2176__;
  wire __2177__;
  wire __2178__;
  wire __2179__;
  wire __2180__;
  wire __2181__;
  wire __2182__;
  wire __2183__;
  wire __2184__;
  wire __2185__;
  wire __2186__;
  wire __2187__;
  wire __2188__;
  wire __2189__;
  wire __2190__;
  wire __2191__;
  wire __2192__;
  wire __2193__;
  wire __2194__;
  wire __2195__;
  wire __2196__;
  wire __2197__;
  wire __2198__;
  wire __2199__;
  wire __2200__;
  wire __2201__;
  wire __2202__;
  wire __2203__;
  wire __2204__;
  wire __2205__;
  wire __2206__;
  wire __2207__;
  wire __2208__;
  wire __2209__;
  wire __2210__;
  wire __2211__;
  wire __2212__;
  wire __2213__;
  wire __2214__;
  wire __2215__;
  wire __2216__;
  wire __2217__;
  wire __2218__;
  wire __2219__;
  wire __2220__;
  wire __2221__;
  wire __2222__;
  wire __2223__;
  wire __2224__;
  wire __2225__;
  wire __2226__;
  wire __2227__;
  wire __2228__;
  wire __2229__;
  wire __2230__;
  wire __2231__;
  wire __2232__;
  wire __2233__;
  wire __2234__;
  wire __2235__;
  wire __2236__;
  wire __2237__;
  wire __2238__;
  wire __2239__;
  wire __2240__;
  wire __2241__;
  wire __2242__;
  wire __2243__;
  wire __2244__;
  wire __2245__;
  wire __2246__;
  wire __2247__;
  wire __2248__;
  wire __2249__;
  wire __2250__;
  wire __2251__;
  wire __2252__;
  wire __2253__;
  wire __2254__;
  wire __2255__;
  wire __2256__;
  wire __2257__;
  wire __2258__;
  wire __2259__;
  wire __2260__;
  wire __2261__;
  wire __2262__;
  wire __2263__;
  wire __2264__;
  wire __2265__;
  wire __2266__;
  wire __2267__;
  wire __2268__;
  wire __2269__;
  wire __2270__;
  wire __2271__;
  wire __2272__;
  wire __2273__;
  wire __2274__;
  wire __2275__;
  wire __2276__;
  wire __2277__;
  wire __2278__;
  wire __2279__;
  wire __2280__;
  wire __2281__;
  wire __2282__;
  wire __2283__;
  wire __2284__;
  wire __2285__;
  wire __2286__;
  wire __2287__;
  wire __2288__;
  wire __2289__;
  wire __2290__;
  wire __2291__;
  wire __2292__;
  wire __2293__;
  wire __2294__;
  wire __2295__;
  wire __2296__;
  wire __2297__;
  wire __2298__;
  wire __2299__;
  wire __2300__;
  wire __2301__;
  wire __2302__;
  wire __2303__;
  wire __2304__;
  wire __2305__;
  wire __2306__;
  wire __2307__;
  wire __2308__;
  wire __2309__;
  wire __2310__;
  wire __2311__;
  wire __2312__;
  wire __2313__;
  wire __2314__;
  wire __2315__;
  wire __2316__;
  wire __2317__;
  wire __2318__;
  wire __2319__;
  wire __2320__;
  wire __2321__;
  wire __2322__;
  wire __2323__;
  wire __2324__;
  wire __2325__;
  wire __2326__;
  wire __2327__;
  wire __2328__;
  wire __2329__;
  wire __2330__;
  wire __2331__;
  wire __2332__;
  wire __2333__;
  wire __2334__;
  wire __2335__;
  wire __2336__;
  wire __2337__;
  wire __2338__;
  wire __2339__;
  wire __2340__;
  wire __2341__;
  wire __2342__;
  wire __2343__;
  wire __2344__;
  wire __2345__;
  wire __2346__;
  wire __2347__;
  wire __2348__;
  wire __2349__;
  wire __2350__;
  wire __2351__;
  wire __2352__;
  wire __2353__;
  wire __2354__;
  wire __2355__;
  wire __2356__;
  wire __2357__;
  wire __2358__;
  wire __2359__;
  wire __2360__;
  wire __2361__;
  wire __2362__;
  wire __2363__;
  wire __2364__;
  wire __2365__;
  wire __2366__;
  wire __2367__;
  wire __2368__;
  wire __2369__;
  wire __2370__;
  wire __2371__;
  wire __2372__;
  wire __2373__;
  wire __2374__;
  wire __2375__;
  wire __2376__;
  wire __2377__;
  wire __2378__;
  wire __2379__;
  wire __2380__;
  wire __2381__;
  wire __2382__;
  wire __2383__;
  wire __2384__;
  wire __2385__;
  wire __2386__;
  wire __2387__;
  wire __2388__;
  wire __2389__;
  wire __2390__;
  wire __2391__;
  wire __2392__;
  wire __2393__;
  wire __2394__;
  wire __2395__;
  wire __2396__;
  wire __2397__;
  wire __2398__;
  wire __2399__;
  wire __2400__;
  wire __2401__;
  wire __2402__;
  wire __2403__;
  wire __2404__;
  wire __2405__;
  wire __2406__;
  wire __2407__;
  wire __2408__;
  wire __2409__;
  wire __2410__;
  wire __2411__;
  wire __2412__;
  wire __2413__;
  wire __2414__;
  wire __2415__;
  wire __2416__;
  wire __2417__;
  wire __2418__;
  wire __2419__;
  wire __2420__;
  wire __2421__;
  wire __2422__;
  wire __2423__;
  wire __2424__;
  wire __2425__;
  wire __2426__;
  wire __2427__;
  wire __2428__;
  wire __2429__;
  wire __2430__;
  wire __2431__;
  wire __2432__;
  wire __2433__;
  wire __2434__;
  wire __2435__;
  wire __2436__;
  wire __2437__;
  wire __2438__;
  wire __2439__;
  wire __2440__;
  wire __2441__;
  wire __2442__;
  wire __2443__;
  wire __2444__;
  wire __2445__;
  wire __2446__;
  wire __2447__;
  wire __2448__;
  wire __2449__;
  wire __2450__;
  wire __2451__;
  wire __2452__;
  wire __2453__;
  wire __2454__;
  wire __2455__;
  wire __2456__;
  wire __2457__;
  wire __2458__;
  wire __2459__;
  wire __2460__;
  wire __2461__;
  wire __2462__;
  wire __2463__;
  wire __2464__;
  wire __2465__;
  wire __2466__;
  wire __2467__;
  wire __2468__;
  wire __2469__;
  wire __2470__;
  wire __2471__;
  wire __2472__;
  wire __2473__;
  wire __2474__;
  wire __2475__;
  wire __2476__;
  wire __2477__;
  wire __2478__;
  wire __2479__;
  wire __2480__;
  wire __2481__;
  wire __2482__;
  wire __2483__;
  wire __2484__;
  wire __2485__;
  wire __2486__;
  wire __2487__;
  wire __2488__;
  wire __2489__;
  wire __2490__;
  wire __2491__;
  wire __2492__;
  wire __2493__;
  wire __2494__;
  wire __2495__;
  wire __2496__;
  wire __2497__;
  wire __2498__;
  wire __2499__;
  wire __2500__;
  wire __2501__;
  wire __2502__;
  wire __2503__;
  wire __2504__;
  wire __2505__;
  wire __2506__;
  wire __2507__;
  wire __2508__;
  wire __2509__;
  wire __2510__;
  wire __2511__;
  wire __2512__;
  wire __2513__;
  wire __2514__;
  wire __2515__;
  wire __2516__;
  wire __2517__;
  wire __2518__;
  wire __2519__;
  wire __2520__;
  wire __2521__;
  wire __2522__;
  wire __2523__;
  wire __2524__;
  wire __2525__;
  wire __2526__;
  wire __2527__;
  wire __2528__;
  wire __2529__;
  wire __2530__;
  wire __2531__;
  wire __2532__;
  wire __2533__;
  wire __2534__;
  wire __2535__;
  wire __2536__;
  wire __2537__;
  wire __2538__;
  wire __2539__;
  wire __2540__;
  wire __2541__;
  wire __2542__;
  wire __2543__;
  wire __2544__;
  wire __2545__;
  wire __2546__;
  wire __2547__;
  wire __2548__;
  wire __2549__;
  wire __2550__;
  wire __2551__;
  wire __2552__;
  wire __2553__;
  wire __2554__;
  wire __2555__;
  wire __2556__;
  wire __2557__;
  wire __2558__;
  wire __2559__;
  wire __2560__;
  wire __2561__;
  wire __2562__;
  wire __2563__;
  wire __2564__;
  wire __2565__;
  wire __2566__;
  wire __2567__;
  wire __2568__;
  wire __2569__;
  wire __2570__;
  wire __2571__;
  wire __2572__;
  wire __2573__;
  wire __2574__;
  wire __2575__;
  wire __2576__;
  wire __2577__;
  wire __2578__;
  wire __2579__;
  wire __2580__;
  wire __2581__;
  wire __2582__;
  wire __2583__;
  wire __2584__;
  wire __2585__;
  wire __2586__;
  wire __2587__;
  wire __2588__;
  wire __2589__;
  wire __2590__;
  wire __2591__;
  wire __2592__;
  wire __2593__;
  wire __2594__;
  wire __2595__;
  wire __2596__;
  wire __2597__;
  wire __2598__;
  wire __2599__;
  wire __2600__;
  wire __2601__;
  wire __2602__;
  wire __2603__;
  wire __2604__;
  wire __2605__;
  wire __2606__;
  wire __2607__;
  wire __2608__;
  wire __2609__;
  wire __2610__;
  wire __2611__;
  wire __2612__;
  wire __2613__;
  wire __2614__;
  wire __2615__;
  wire __2616__;
  wire __2617__;
  wire __2618__;
  wire __2619__;
  wire __2620__;
  wire __2621__;
  wire __2622__;
  wire __2623__;
  wire __2624__;
  wire __2625__;
  wire __2626__;
  wire __2627__;
  wire __2628__;
  wire __2629__;
  wire __2630__;
  wire __2631__;
  wire __2632__;
  wire __2633__;
  wire __2634__;
  wire __2635__;
  wire __2636__;
  wire __2637__;
  wire __2638__;
  wire __2639__;
  wire __2640__;
  wire __2641__;
  wire __2642__;
  wire __2643__;
  wire __2644__;
  wire __2645__;
  wire __2646__;
  wire __2647__;
  wire __2648__;
  wire __2649__;
  wire __2650__;
  wire __2651__;
  wire __2652__;
  wire __2653__;
  wire __2654__;
  wire __2655__;
  wire __2656__;
  wire __2657__;
  wire __2658__;
  wire __2659__;
  wire __2660__;
  wire __2661__;
  wire __2662__;
  wire __2663__;
  wire __2664__;
  wire __2665__;
  wire __2666__;
  wire __2667__;
  wire __2668__;
  wire __2669__;
  wire __2670__;
  wire __2671__;
  wire __2672__;
  wire __2673__;
  wire __2674__;
  wire __2675__;
  wire __2676__;
  wire __2677__;
  wire __2678__;
  wire __2679__;
  wire __2680__;
  wire __2681__;
  wire __2682__;
  wire __2683__;
  wire __2684__;
  wire __2685__;
  wire __2686__;
  wire __2687__;
  wire __2688__;
  wire __2689__;
  wire __2690__;
  wire __2691__;
  wire __2692__;
  wire __2693__;
  wire __2694__;
  wire __2695__;
  wire __2696__;
  wire __2697__;
  wire __2698__;
  wire __2699__;
  wire __2700__;
  wire __2701__;
  wire __2702__;
  wire __2703__;
  wire __2704__;
  wire __2705__;
  wire __2706__;
  wire __2707__;
  wire __2708__;
  wire __2709__;
  wire __2710__;
  wire __2711__;
  wire __2712__;
  wire __2713__;
  wire __2714__;
  wire __2715__;
  wire __2716__;
  wire __2717__;
  wire __2718__;
  wire __2719__;
  wire __2720__;
  wire __2721__;
  wire __2722__;
  wire __2723__;
  wire __2724__;
  wire __2725__;
  wire __2726__;
  wire __2727__;
  wire __2728__;
  wire __2729__;
  wire __2730__;
  wire __2731__;
  wire __2732__;
  wire __2733__;
  wire __2734__;
  wire __2735__;
  wire __2736__;
  wire __2737__;
  wire __2738__;
  wire __2739__;
  wire __2740__;
  wire __2741__;
  wire __2742__;
  wire __2743__;
  wire __2744__;
  wire __2745__;
  wire __2746__;
  wire __2747__;
  wire __2748__;
  wire __2749__;
  wire __2750__;
  wire __2751__;
  wire __2752__;
  wire __2753__;
  wire __2754__;
  wire __2755__;
  wire __2756__;
  wire __2757__;
  wire __2758__;
  wire __2759__;
  wire __2760__;
  wire __2761__;
  wire __2762__;
  wire __2763__;
  wire __2764__;
  wire __2765__;
  wire __2766__;
  wire __2767__;
  wire __2768__;
  wire __2769__;
  wire __2770__;
  wire __2771__;
  wire __2772__;
  wire __2773__;
  wire __2774__;
  wire __2775__;
  wire __2776__;
  wire __2777__;
  wire __2778__;
  wire __2779__;
  wire __2780__;
  wire __2781__;
  wire __2782__;
  wire __2783__;
  wire __2784__;
  wire __2785__;
  wire __2786__;
  wire __2787__;
  wire __2788__;
  wire __2789__;
  wire __2790__;
  wire __2791__;
  wire __2792__;
  wire __2793__;
  wire __2794__;
  wire __2795__;
  wire __2796__;
  wire __2797__;
  wire __2798__;
  wire __2799__;
  wire __2800__;
  wire __2801__;
  wire __2802__;
  wire __2803__;
  wire __2804__;
  wire __2805__;
  wire __2806__;
  wire __2807__;
  wire __2808__;
  wire __2809__;
  wire __2810__;
  wire __2811__;
  wire __2812__;
  wire __2813__;
  wire __2814__;
  wire __2815__;
  wire __2816__;
  wire __2817__;
  wire __2818__;
  wire __2819__;
  wire __2820__;
  wire __2821__;
  wire __2822__;
  wire __2823__;
  wire __2824__;
  wire __2825__;
  wire __2826__;
  wire __2827__;
  wire __2828__;
  wire __2829__;
  wire __2830__;
  wire __2831__;
  wire __2832__;
  wire __2833__;
  wire __2834__;
  wire __2835__;
  wire __2836__;
  wire __2837__;
  wire __2838__;
  wire __2839__;
  wire __2840__;
  wire __2841__;
  wire __2842__;
  wire __2843__;
  wire __2844__;
  wire __2845__;
  wire __2846__;
  wire __2847__;
  wire __2848__;
  wire __2849__;
  wire __2850__;
  wire __2851__;
  wire __2852__;
  wire __2853__;
  wire __2854__;
  wire __2855__;
  wire __2856__;
  wire __2857__;
  wire __2858__;
  wire __2859__;
  wire __2860__;
  wire __2861__;
  wire __2862__;
  wire __2863__;
  wire __2864__;
  wire __2865__;
  wire __2866__;
  wire __2867__;
  wire __2868__;
  wire __2869__;
  wire __2870__;
  wire __2871__;
  wire __2872__;
  wire __2873__;
  wire __2874__;
  wire __2875__;
  wire __2876__;
  wire __2877__;
  wire __2878__;
  wire __2879__;
  wire __2880__;
  wire __2881__;
  wire __2882__;
  wire __2883__;
  wire __2884__;
  wire __2885__;
  wire __2886__;
  wire __2887__;
  wire __2888__;
  wire __2889__;
  wire __2890__;
  wire __2891__;
  wire __2892__;
  wire __2893__;
  wire __2894__;
  wire __2895__;
  wire __2896__;
  wire __2897__;
  wire __2898__;
  wire __2899__;
  wire __2900__;
  wire __2901__;
  wire __2902__;
  wire __2903__;
  wire __2904__;
  wire __2905__;
  wire __2906__;
  wire __2907__;
  wire __2908__;
  wire __2909__;
  wire __2910__;
  wire __2911__;
  wire __2912__;
  wire __2913__;
  wire __2914__;
  wire __2915__;
  wire __2916__;
  wire __2917__;
  wire __2918__;
  wire __2919__;
  wire __2920__;
  wire __2921__;
  wire __2922__;
  wire __2923__;
  wire __2924__;
  wire __2925__;
  wire __2926__;
  wire __2927__;
  wire __2928__;
  wire __2929__;
  wire __2930__;
  wire __2931__;
  wire __2932__;
  wire __2933__;
  wire __2934__;
  wire __2935__;
  wire __2936__;
  wire __2937__;
  wire __2938__;
  wire __2939__;
  wire __2940__;
  wire __2941__;
  wire __2942__;
  wire __2943__;
  wire __2944__;
  wire __2945__;
  wire __2946__;
  wire __2947__;
  wire __2948__;
  wire __2949__;
  wire __2950__;
  wire __2951__;
  wire __2952__;
  wire __2953__;
  wire __2954__;
  wire __2955__;
  wire __2956__;
  wire __2957__;
  wire __2958__;
  wire __2959__;
  wire __2960__;
  wire __2961__;
  wire __2962__;
  wire __2963__;
  wire __2964__;
  wire __2965__;
  wire __2966__;
  wire __2967__;
  wire __2968__;
  wire __2969__;
  wire __2970__;
  wire __2971__;
  wire __2972__;
  wire __2973__;
  wire __2974__;
  wire __2975__;
  wire __2976__;
  wire __2977__;
  wire __2978__;
  wire __2979__;
  wire __2980__;
  wire __2981__;
  wire __2982__;
  wire __2983__;
  wire __2984__;
  wire __2985__;
  wire __2986__;
  wire __2987__;
  wire __2988__;
  wire __2989__;
  wire __2990__;
  wire __2991__;
  wire __2992__;
  wire __2993__;
  wire __2994__;
  wire __2995__;
  wire __2996__;
  wire __2997__;
  wire __2998__;
  wire __2999__;
  wire __3000__;
  wire __3001__;
  wire __3002__;
  wire __3003__;
  wire __3004__;
  wire __3005__;
  wire __3006__;
  wire __3007__;
  wire __3008__;
  wire __3009__;
  wire __3010__;
  wire __3011__;
  wire __3012__;
  wire __3013__;
  wire __3014__;
  wire __3015__;
  wire __3016__;
  wire __3017__;
  wire __3018__;
  wire __3019__;
  wire __3020__;
  wire __3021__;
  wire __3022__;
  wire __3023__;
  wire __3024__;
  wire __3025__;
  wire __3026__;
  wire __3027__;
  wire __3028__;
  wire __3029__;
  wire __3030__;
  wire __3031__;
  wire __3032__;
  wire __3033__;
  wire __3034__;
  wire __3035__;
  wire __3036__;
  wire __3037__;
  wire __3038__;
  wire __3039__;
  wire __3040__;
  wire __3041__;
  wire __3042__;
  wire __3043__;
  wire __3044__;
  wire __3045__;
  wire __3046__;
  wire __3047__;
  wire __3048__;
  wire __3049__;
  wire __3050__;
  wire __3051__;
  wire __3052__;
  wire __3053__;
  wire __3054__;
  wire __3055__;
  wire __3056__;
  wire __3057__;
  wire __3058__;
  wire __3059__;
  wire __3060__;
  wire __3061__;
  wire __3062__;
  wire __3063__;
  wire __3064__;
  wire __3065__;
  wire __3066__;
  wire __3067__;
  wire __3068__;
  wire __3069__;
  wire __3070__;
  wire __3071__;
  wire __3072__;
  wire __3073__;
  wire __3074__;
  wire __3075__;
  wire __3076__;
  wire __3077__;
  wire __3078__;
  wire __3079__;
  wire __3080__;
  wire __3081__;
  wire __3082__;
  wire __3083__;
  wire __3084__;
  wire __3085__;
  wire __3086__;
  wire __3087__;
  wire __3088__;
  wire __3089__;
  wire __3090__;
  wire __3091__;
  wire __3092__;
  wire __3093__;
  wire __3094__;
  wire __3095__;
  wire __3096__;
  wire __3097__;
  wire __3098__;
  wire __3099__;
  wire __3100__;
  wire __3101__;
  wire __3102__;
  wire __3103__;
  wire __3104__;
  wire __3105__;
  wire __3106__;
  wire __3107__;
  wire __3108__;
  wire __3109__;
  wire __3110__;
  wire __3111__;
  wire __3112__;
  wire __3113__;
  wire __3114__;
  wire __3115__;
  wire __3116__;
  wire __3117__;
  wire __3118__;
  wire __3119__;
  wire __3120__;
  wire __3121__;
  wire __3122__;
  wire __3123__;
  wire __3124__;
  wire __3125__;
  wire __3126__;
  wire __3127__;
  wire __3128__;
  wire __3129__;
  wire __3130__;
  wire __3131__;
  wire __3132__;
  wire __3133__;
  wire __3134__;
  wire __3135__;
  wire __3136__;
  wire __3137__;
  wire __3138__;
  wire __3139__;
  wire __3140__;
  wire __3141__;
  wire __3142__;
  wire __3143__;
  wire __3144__;
  wire __3145__;
  wire __3146__;
  wire __3147__;
  wire __3148__;
  wire __3149__;
  wire __3150__;
  wire __3151__;
  wire __3152__;
  wire __3153__;
  wire __3154__;
  wire __3155__;
  wire __3156__;
  wire __3157__;
  wire __3158__;
  wire __3159__;
  wire __3160__;
  wire __3161__;
  wire __3162__;
  wire __3163__;
  wire __3164__;
  wire __3165__;
  wire __3166__;
  wire __3167__;
  wire __3168__;
  wire __3169__;
  wire __3170__;
  wire __3171__;
  wire __3172__;
  wire __3173__;
  wire __3174__;
  wire __3175__;
  wire __3176__;
  wire __3177__;
  wire __3178__;
  wire __3179__;
  wire __3180__;
  wire __3181__;
  wire __3182__;
  wire __3183__;
  wire __3184__;
  wire __3185__;
  wire __3186__;
  wire __3187__;
  wire __3188__;
  wire __3189__;
  wire __3190__;
  wire __3191__;
  wire __3192__;
  wire __3193__;
  wire __3194__;
  wire __3195__;
  wire __3196__;
  wire __3197__;
  wire __3198__;
  wire __3199__;
  wire __3200__;
  wire __3201__;
  wire __3202__;
  wire __3203__;
  wire __3204__;
  wire __3205__;
  wire __3206__;
  wire __3207__;
  wire __3208__;
  wire __3209__;
  wire __3210__;
  wire __3211__;
  wire __3212__;
  wire __3213__;
  wire __3214__;
  wire __3215__;
  wire __3216__;
  wire __3217__;
  wire __3218__;
  wire __3219__;
  wire __3220__;
  wire __3221__;
  wire __3222__;
  wire __3223__;
  wire __3224__;
  wire __3225__;
  wire __3226__;
  wire __3227__;
  wire __3228__;
  wire __3229__;
  wire __3230__;
  wire __3231__;
  wire __3232__;
  wire __3233__;
  wire __3234__;
  wire __3235__;
  wire __3236__;
  wire __3237__;
  wire __3238__;
  wire __3239__;
  wire __3240__;
  wire __3241__;
  wire __3242__;
  wire __3243__;
  wire __3244__;
  wire __3245__;
  wire __3246__;
  wire __3247__;
  wire __3248__;
  wire __3249__;
  wire __3250__;
  wire __3251__;
  wire __3252__;
  wire __3253__;
  wire __3254__;
  wire __3255__;
  wire __3256__;
  wire __3257__;
  wire __3258__;
  wire __3259__;
  wire __3260__;
  wire __3261__;
  wire __3262__;
  wire __3263__;
  wire __3264__;
  wire __3265__;
  wire __3266__;
  wire __3267__;
  wire __3268__;
  wire __3269__;
  wire __3270__;
  wire __3271__;
  wire __3272__;
  wire __3273__;
  wire __3274__;
  wire __3275__;
  wire __3276__;
  wire __3277__;
  wire __3278__;
  wire __3279__;
  wire __3280__;
  wire __3281__;
  wire __3282__;
  wire __3283__;
  wire __3284__;
  wire __3285__;
  wire __3286__;
  wire __3287__;
  wire __3288__;
  wire __3289__;
  wire __3290__;
  wire __3291__;
  wire __3292__;
  wire __3293__;
  wire __3294__;
  wire __3295__;
  wire __3296__;
  wire __3297__;
  wire __3298__;
  wire __3299__;
  wire __3300__;
  wire __3301__;
  wire __3302__;
  wire __3303__;
  wire __3304__;
  wire __3305__;
  wire __3306__;
  wire __3307__;
  wire __3308__;
  wire __3309__;
  wire __3310__;
  wire __3311__;
  wire __3312__;
  wire __3313__;
  wire __3314__;
  wire __3315__;
  wire __3316__;
  wire __3317__;
  wire __3318__;
  wire __3319__;
  wire __3320__;
  wire __3321__;
  wire __3322__;
  wire __3323__;
  wire __3324__;
  wire __3325__;
  wire __3326__;
  wire __3327__;
  wire __3328__;
  wire __3329__;
  wire __3330__;
  wire __3331__;
  wire __3332__;
  wire __3333__;
  wire __3334__;
  wire __3335__;
  wire __3336__;
  wire __3337__;
  wire __3338__;
  wire __3339__;
  wire __3340__;
  wire __3341__;
  wire __3342__;
  wire __3343__;
  wire __3344__;
  wire __3345__;
  wire __3346__;
  wire __3347__;
  wire __3348__;
  wire __3349__;
  wire __3350__;
  wire __3351__;
  wire __3352__;
  wire __3353__;
  wire __3354__;
  wire __3355__;
  wire __3356__;
  wire __3357__;
  wire __3358__;
  wire __3359__;
  wire __3360__;
  wire __3361__;
  wire __3362__;
  wire __3363__;
  wire __3364__;
  wire __3365__;
  wire __3366__;
  wire __3367__;
  wire __3368__;
  wire __3369__;
  wire __3370__;
  wire __3371__;
  wire __3372__;
  wire __3373__;
  wire __3374__;
  wire __3375__;
  wire __3376__;
  wire __3377__;
  wire __3378__;
  wire __3379__;
  INV __3380__ (
    .I(__1__),
    .O(__0__)
  );
  LUT4 #(
    .INIT(16'h4000)
  ) __3381__ (
    .I3(__1100__),
    .I2(__876__),
    .I1(__825__),
    .I0(__720__),
    .O(__1__)
  );
  INV __3382__ (
    .I(__868__),
    .O(__2__)
  );
  INV __3383__ (
    .I(__535__),
    .O(__3__)
  );
  INV __3384__ (
    .I(__221__),
    .O(__4__)
  );
  INV __3385__ (
    .I(g5),
    .O(__5__)
  );
  INV __3386__ (
    .I(__884__),
    .O(__6__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3387__ (
    .D(__3230__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__7__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3388__ (
    .D(__2731__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__8__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3389__ (
    .D(__2605__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__9__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3390__ (
    .D(__2692__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__10__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3391__ (
    .D(__3069__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__11__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3392__ (
    .D(__3330__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__12__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3393__ (
    .D(__1719__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__13__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3394__ (
    .D(__3178__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__14__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3395__ (
    .D(__3344__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__15__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3396__ (
    .D(__3265__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__16__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3397__ (
    .D(__2598__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__17__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3398__ (
    .D(__2578__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__18__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3399__ (
    .D(__1985__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__19__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3400__ (
    .D(__2165__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__20__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3401__ (
    .D(__1699__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__21__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3402__ (
    .D(__2655__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__22__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3403__ (
    .D(__2703__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__23__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3404__ (
    .D(__2262__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__24__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3405__ (
    .D(__2200__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__25__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3406__ (
    .D(__1829__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__26__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3407__ (
    .D(__3010__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__27__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3408__ (
    .D(__1834__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__28__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3409__ (
    .D(__2422__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__29__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3410__ (
    .D(__1276__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__30__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3411__ (
    .D(__3177__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__31__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3412__ (
    .D(__2669__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__32__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3413__ (
    .D(__2894__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__33__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3414__ (
    .D(__2249__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__34__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3415__ (
    .D(__2843__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__35__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3416__ (
    .D(__2038__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__36__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3417__ (
    .D(__1693__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__37__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3418__ (
    .D(__1505__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__38__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3419__ (
    .D(__2180__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__39__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3420__ (
    .D(__2914__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__40__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3421__ (
    .D(__1802__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__41__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3422__ (
    .D(__1940__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__42__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3423__ (
    .D(__2985__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__43__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3424__ (
    .D(__2003__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__44__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3425__ (
    .D(__502__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__45__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3426__ (
    .D(__2581__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__46__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3427__ (
    .D(__2998__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__47__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3428__ (
    .D(__994__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__48__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3429__ (
    .D(__521__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__49__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3430__ (
    .D(__2082__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__50__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3431__ (
    .D(__2988__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__51__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3432__ (
    .D(__1878__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__52__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3433__ (
    .D(__3257__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__53__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3434__ (
    .D(__2406__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__54__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3435__ (
    .D(__3083__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__55__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3436__ (
    .D(__635__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__56__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3437__ (
    .D(__2547__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__57__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3438__ (
    .D(__1787__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__58__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3439__ (
    .D(__1169__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__59__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3440__ (
    .D(__1675__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__60__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3441__ (
    .D(__2256__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__61__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3442__ (
    .D(__2971__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__62__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3443__ (
    .D(__2176__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__63__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3444__ (
    .D(__1982__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__64__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3445__ (
    .D(__3349__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__65__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3446__ (
    .D(__2958__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__66__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3447__ (
    .D(__2327__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__67__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3448__ (
    .D(__3352__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__68__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3449__ (
    .D(__2463__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__69__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3450__ (
    .D(__1601__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__70__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3451__ (
    .D(__945__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__71__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3452__ (
    .D(__887__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__72__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3453__ (
    .D(__3333__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__73__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3454__ (
    .D(__1879__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__74__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3455__ (
    .D(__1174__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__75__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3456__ (
    .D(__2380__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__76__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3457__ (
    .D(__2897__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__77__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3458__ (
    .D(__1641__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__78__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3459__ (
    .D(__3320__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__79__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3460__ (
    .D(__419__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__80__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3461__ (
    .D(__2170__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__81__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3462__ (
    .D(__2714__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__82__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3463__ (
    .D(__2590__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__83__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3464__ (
    .D(__1513__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__84__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3465__ (
    .D(__2167__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__85__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3466__ (
    .D(__3249__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__86__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3467__ (
    .D(__3308__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__87__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3468__ (
    .D(__2009__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__88__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3469__ (
    .D(__3074__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__89__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3470__ (
    .D(__42__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__90__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3471__ (
    .D(__2732__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__91__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3472__ (
    .D(__2764__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__92__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3473__ (
    .D(__401__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__93__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3474__ (
    .D(__1764__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__94__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3475__ (
    .D(__3209__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__95__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3476__ (
    .D(__1935__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__96__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3477__ (
    .D(__2926__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__97__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3478__ (
    .D(__398__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__98__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3479__ (
    .D(__3323__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__99__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3480__ (
    .D(__2942__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__100__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3481__ (
    .D(__1560__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__101__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3482__ (
    .D(__3263__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__102__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3483__ (
    .D(__1199__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__103__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3484__ (
    .D(__2723__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__104__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3485__ (
    .D(__991__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__105__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3486__ (
    .D(__1495__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__106__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3487__ (
    .D(__2369__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__107__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3488__ (
    .D(__2702__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__108__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3489__ (
    .D(__1966__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__109__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3490__ (
    .D(__3235__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__110__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3491__ (
    .D(__2973__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__111__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3492__ (
    .D(__1524__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__112__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3493__ (
    .D(__2927__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__113__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3494__ (
    .D(__2987__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__114__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3495__ (
    .D(__873__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__115__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3496__ (
    .D(__2676__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__116__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3497__ (
    .D(__1991__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__117__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3498__ (
    .D(__2139__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__118__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3499__ (
    .D(__2001__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__119__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3500__ (
    .D(__1726__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__120__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3501__ (
    .D(__2431__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__121__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3502__ (
    .D(__155__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__122__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3503__ (
    .D(__3003__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__123__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3504__ (
    .D(__2948__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__124__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3505__ (
    .D(__2696__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__125__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3506__ (
    .D(__2025__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__126__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3507__ (
    .D(__2332__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__127__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3508__ (
    .D(__1703__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__128__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3509__ (
    .D(__1607__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__129__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3510__ (
    .D(__2993__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__130__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3511__ (
    .D(__3141__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__131__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3512__ (
    .D(__1860__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__132__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3513__ (
    .D(__122__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__133__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3514__ (
    .D(__2366__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__134__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3515__ (
    .D(__2517__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__135__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3516__ (
    .D(__2452__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__136__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3517__ (
    .D(__3222__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__137__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3518__ (
    .D(__2573__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__138__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3519__ (
    .D(__2064__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__139__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3520__ (
    .D(__1851__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__140__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3521__ (
    .D(__1997__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__141__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3522__ (
    .D(__1467__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__142__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3523__ (
    .D(__1961__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__143__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3524__ (
    .D(__1705__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__144__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3525__ (
    .D(__3057__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__145__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3526__ (
    .D(__3150__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__146__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3527__ (
    .D(__1875__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__147__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3528__ (
    .D(__2747__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__148__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3529__ (
    .D(__2979__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__149__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3530__ (
    .D(__3281__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__150__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3531__ (
    .D(__2653__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__151__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3532__ (
    .D(__3085__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__152__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3533__ (
    .D(__3035__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__153__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3534__ (
    .D(__2242__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__154__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3535__ (
    .D(__759__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__155__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3536__ (
    .D(__2473__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__156__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3537__ (
    .D(__3369__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__157__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3538__ (
    .D(__1308__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__158__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3539__ (
    .D(__1767__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__159__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3540__ (
    .D(__45__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__160__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3541__ (
    .D(__2217__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__161__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3542__ (
    .D(__2362__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__162__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3543__ (
    .D(__2710__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__163__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3544__ (
    .D(__2925__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__164__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3545__ (
    .D(__2886__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__165__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3546__ (
    .D(__3219__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__166__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3547__ (
    .D(__2481__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__167__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3548__ (
    .D(__484__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__168__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3549__ (
    .D(__257__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__169__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3550__ (
    .D(__2045__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__170__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3551__ (
    .D(__2333__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__171__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3552__ (
    .D(__3239__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__172__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3553__ (
    .D(__2742__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__173__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3554__ (
    .D(__2684__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__174__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3555__ (
    .D(__2325__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__175__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3556__ (
    .D(__2390__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__176__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3557__ (
    .D(__2870__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__177__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3558__ (
    .D(__2893__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__178__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3559__ (
    .D(__2799__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__179__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3560__ (
    .D(__329__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__180__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3561__ (
    .D(__208__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__181__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3562__ (
    .D(__2393__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__182__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3563__ (
    .D(__3192__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__183__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3564__ (
    .D(__2370__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__184__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3565__ (
    .D(__3300__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__185__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3566__ (
    .D(__1985__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__186__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3567__ (
    .D(__103__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__187__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3568__ (
    .D(__1962__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__188__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3569__ (
    .D(__1635__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__189__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3570__ (
    .D(__1796__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__190__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3571__ (
    .D(__3268__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__191__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3572__ (
    .D(__481__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__192__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3573__ (
    .D(__2589__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__193__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3574__ (
    .D(__1867__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__194__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3575__ (
    .D(__3182__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__195__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3576__ (
    .D(__1490__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__196__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3577__ (
    .D(__1989__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__197__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3578__ (
    .D(__1865__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__198__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3579__ (
    .D(__1457__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__199__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3580__ (
    .D(__3054__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__200__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3581__ (
    .D(__3350__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__201__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3582__ (
    .D(__3071__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__202__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3583__ (
    .D(__2608__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__203__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3584__ (
    .D(__2472__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__204__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3585__ (
    .D(__2096__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__205__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3586__ (
    .D(__1419__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__206__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3587__ (
    .D(__1789__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__207__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3588__ (
    .D(__133__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__208__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3589__ (
    .D(__2778__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__209__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3590__ (
    .D(__2912__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__210__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3591__ (
    .D(__1666__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__211__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3592__ (
    .D(__3197__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__212__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3593__ (
    .D(__859__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__213__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3594__ (
    .D(__3363__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__214__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3595__ (
    .D(__433__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__215__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3596__ (
    .D(__3366__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__216__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3597__ (
    .D(__56__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__217__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3598__ (
    .D(__3040__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__218__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3599__ (
    .D(__3128__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__219__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3600__ (
    .D(__3294__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__220__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3601__ (
    .D(__3240__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__221__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3602__ (
    .D(__2345__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__222__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3603__ (
    .D(__1669__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__223__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3604__ (
    .D(__3236__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__224__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3605__ (
    .D(__1639__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__225__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3606__ (
    .D(__2442__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__226__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3607__ (
    .D(__2603__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__227__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3608__ (
    .D(__3125__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__228__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3609__ (
    .D(__2319__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__229__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3610__ (
    .D(__19__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__230__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3611__ (
    .D(__1582__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__231__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3612__ (
    .D(__3140__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__232__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3613__ (
    .D(__2644__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__233__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3614__ (
    .D(__1795__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__234__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3615__ (
    .D(__2004__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__235__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3616__ (
    .D(__2059__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__236__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3617__ (
    .D(__1510__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__237__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3618__ (
    .D(__2458__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__238__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3619__ (
    .D(__2204__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__239__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3620__ (
    .D(__1821__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__240__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3621__ (
    .D(__2048__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__241__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3622__ (
    .D(__3309__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__242__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3623__ (
    .D(__3278__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__243__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3624__ (
    .D(__1784__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__244__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3625__ (
    .D(__1695__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__245__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3626__ (
    .D(__3145__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__246__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3627__ (
    .D(__2818__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__247__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3628__ (
    .D(__2124__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__248__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3629__ (
    .D(__3046__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__249__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3630__ (
    .D(__3187__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__250__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3631__ (
    .D(__2042__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__251__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3632__ (
    .D(__3335__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__252__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3633__ (
    .D(__2878__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__253__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3634__ (
    .D(__1631__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__254__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3635__ (
    .D(__2267__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__255__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3636__ (
    .D(__1209__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__256__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3637__ (
    .D(__815__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__257__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3638__ (
    .D(__1848__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__258__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3639__ (
    .D(__661__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__259__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3640__ (
    .D(__1870__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__260__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3641__ (
    .D(__2041__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__261__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3642__ (
    .D(__966__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__262__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3643__ (
    .D(__684__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__263__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3644__ (
    .D(__2911__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__264__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3645__ (
    .D(__1882__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__265__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3646__ (
    .D(__2483__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__266__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3647__ (
    .D(__3058__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__267__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3648__ (
    .D(__2277__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__268__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3649__ (
    .D(__3188__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__269__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3650__ (
    .D(__2273__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__270__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3651__ (
    .D(__3062__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__271__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3652__ (
    .D(__2875__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__272__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3653__ (
    .D(__2990__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__273__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3654__ (
    .D(__3109__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__274__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3655__ (
    .D(__3139__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__275__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3656__ (
    .D(__328__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__276__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3657__ (
    .D(__2745__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__277__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3658__ (
    .D(__3365__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__278__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3659__ (
    .D(__973__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__279__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3660__ (
    .D(__3354__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__280__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3661__ (
    .D(__2807__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__281__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3662__ (
    .D(__2751__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__282__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3663__ (
    .D(__3207__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__283__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3664__ (
    .D(__2810__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__284__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3665__ (
    .D(__2805__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__285__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3666__ (
    .D(__3317__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__286__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3667__ (
    .D(__186__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__287__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3668__ (
    .D(__1877__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__288__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3669__ (
    .D(__3081__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__289__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3670__ (
    .D(__2238__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__290__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3671__ (
    .D(__2735__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__291__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3672__ (
    .D(__1797__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__292__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3673__ (
    .D(__1293__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__293__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3674__ (
    .D(__1624__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__294__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3675__ (
    .D(__3204__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__295__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3676__ (
    .D(__2957__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__296__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3677__ (
    .D(__2673__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__297__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3678__ (
    .D(__2741__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__298__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3679__ (
    .D(__2480__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__299__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3680__ (
    .D(__3302__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__300__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3681__ (
    .D(__1873__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__301__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3682__ (
    .D(__451__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__302__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3683__ (
    .D(__2008__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__303__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3684__ (
    .D(__2498__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__304__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3685__ (
    .D(__526__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__305__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3686__ (
    .D(__2478__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__306__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3687__ (
    .D(__2774__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__307__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3688__ (
    .D(__2769__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__308__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3689__ (
    .D(__3000__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__309__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3690__ (
    .D(__2316__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__310__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3691__ (
    .D(__2251__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__311__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3692__ (
    .D(__98__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__312__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3693__ (
    .D(__2921__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__313__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3694__ (
    .D(__3331__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__314__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3695__ (
    .D(__1653__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__315__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3696__ (
    .D(__3001__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__316__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3697__ (
    .D(__2479__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__317__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3698__ (
    .D(__2462__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__318__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3699__ (
    .D(__2030__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__319__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3700__ (
    .D(__239__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__320__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3701__ (
    .D(__3167__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__321__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3702__ (
    .D(__1804__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__322__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3703__ (
    .D(__2241__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__323__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3704__ (
    .D(__1792__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__324__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3705__ (
    .D(__2121__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__325__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3706__ (
    .D(__3132__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__326__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3707__ (
    .D(__3097__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__327__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3708__ (
    .D(__2443__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__328__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3709__ (
    .D(__486__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__329__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3710__ (
    .D(__371__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__330__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3711__ (
    .D(__3228__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__331__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3712__ (
    .D(__2652__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__332__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3713__ (
    .D(__1542__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__333__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3714__ (
    .D(__2756__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__334__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3715__ (
    .D(__3008__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__335__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3716__ (
    .D(__2036__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__336__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3717__ (
    .D(__2708__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__337__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3718__ (
    .D(__2275__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__338__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3719__ (
    .D(__3162__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__339__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3720__ (
    .D(__3237__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__340__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3721__ (
    .D(__2970__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__341__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3722__ (
    .D(__1753__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__342__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3723__ (
    .D(__2436__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__343__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3724__ (
    .D(__2657__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__344__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3725__ (
    .D(__2687__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__345__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3726__ (
    .D(__1097__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__346__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3727__ (
    .D(__2339__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__347__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3728__ (
    .D(__1390__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__348__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3729__ (
    .D(__979__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__349__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3730__ (
    .D(__1963__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__350__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3731__ (
    .D(__1040__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__351__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3732__ (
    .D(__2749__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__352__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3733__ (
    .D(__2456__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__353__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3734__ (
    .D(__3195__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__354__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3735__ (
    .D(__2407__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__355__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3736__ (
    .D(__2376__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__356__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3737__ (
    .D(__1671__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__357__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3738__ (
    .D(__2984__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__358__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3739__ (
    .D(__115__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__359__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3740__ (
    .D(__3180__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__360__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3741__ (
    .D(__1332__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__361__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3742__ (
    .D(__1676__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__362__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3743__ (
    .D(__2392__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__363__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3744__ (
    .D(__1702__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__364__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3745__ (
    .D(__3307__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__365__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3746__ (
    .D(__774__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__366__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3747__ (
    .D(__2032__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__367__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3748__ (
    .D(__1917__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__368__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3749__ (
    .D(__2740__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__369__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3750__ (
    .D(__2896__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__370__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3751__ (
    .D(__48__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__371__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3752__ (
    .D(__2722__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__372__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3753__ (
    .D(__2753__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__373__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3754__ (
    .D(__3297__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__374__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3755__ (
    .D(__3196__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__375__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3756__ (
    .D(__1765__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__376__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3757__ (
    .D(__2727__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__377__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3758__ (
    .D(__2931__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__378__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3759__ (
    .D(__3095__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__379__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3760__ (
    .D(__674__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__380__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3761__ (
    .D(__1580__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__381__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3762__ (
    .D(__3324__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__382__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3763__ (
    .D(__1714__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__383__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3764__ (
    .D(__3151__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__384__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3765__ (
    .D(__998__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__385__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3766__ (
    .D(__1304__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__386__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3767__ (
    .D(__1618__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__387__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3768__ (
    .D(__2699__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__388__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3769__ (
    .D(__2401__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__389__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3770__ (
    .D(__2693__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__390__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3771__ (
    .D(__3316__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__391__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3772__ (
    .D(__3030__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__392__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3773__ (
    .D(__3328__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__393__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3774__ (
    .D(__612__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__394__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3775__ (
    .D(__3111__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__395__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3776__ (
    .D(__2391__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__396__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3777__ (
    .D(__1453__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__397__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3778__ (
    .D(__1006__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__398__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3779__ (
    .D(__2244__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__399__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3780__ (
    .D(__3373__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__400__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3781__ (
    .D(__1691__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__401__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3782__ (
    .D(__2642__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__402__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3783__ (
    .D(__1550__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__403__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3784__ (
    .D(__2280__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__404__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3785__ (
    .D(__2607__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__405__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3786__ (
    .D(__3103__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__406__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3787__ (
    .D(__2396__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__407__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3788__ (
    .D(__3273__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__408__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3789__ (
    .D(__3199__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__409__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3790__ (
    .D(__2949__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__410__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3791__ (
    .D(__2024__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__411__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3792__ (
    .D(__2183__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__412__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3793__ (
    .D(__2871__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__413__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3794__ (
    .D(__2899__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__414__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3795__ (
    .D(__2618__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__415__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3796__ (
    .D(__312__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__416__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3797__ (
    .D(__2447__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__417__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3798__ (
    .D(__1968__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__418__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3799__ (
    .D(__3227__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__419__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3800__ (
    .D(__2648__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__420__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3801__ (
    .D(__1824__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__421__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3802__ (
    .D(__3348__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__422__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3803__ (
    .D(__3090__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__423__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3804__ (
    .D(__2937__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__424__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3805__ (
    .D(__2647__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__425__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3806__ (
    .D(__3021__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__426__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3807__ (
    .D(__3166__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__427__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3808__ (
    .D(__3127__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__428__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3809__ (
    .D(__2615__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__429__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3810__ (
    .D(__2953__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__430__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3811__ (
    .D(__2705__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__431__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3812__ (
    .D(__2960__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__432__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3813__ (
    .D(__259__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__433__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3814__ (
    .D(__3190__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__434__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3815__ (
    .D(__3272__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__435__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3816__ (
    .D(__3060__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__436__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3817__ (
    .D(__2348__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__437__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3818__ (
    .D(__2808__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__438__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3819__ (
    .D(__3117__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__439__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3820__ (
    .D(__2518__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__440__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3821__ (
    .D(__1629__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__441__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3822__ (
    .D(__160__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__442__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3823__ (
    .D(__2082__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__443__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3824__ (
    .D(__2748__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__444__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3825__ (
    .D(__2771__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__445__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3826__ (
    .D(__3244__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__446__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3827__ (
    .D(__2766__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__447__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3828__ (
    .D(__2207__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__448__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3829__ (
    .D(__3376__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__449__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3830__ (
    .D(__573__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__450__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3831__ (
    .D(__2864__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__451__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3832__ (
    .D(__3318__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__452__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3833__ (
    .D(__2679__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__453__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3834__ (
    .D(__2809__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__454__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3835__ (
    .D(__3255__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__455__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3836__ (
    .D(__3339__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__456__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3837__ (
    .D(__1296__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__457__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3838__ (
    .D(__2733__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__458__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3839__ (
    .D(__2454__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__459__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3840__ (
    .D(__3047__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__460__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3841__ (
    .D(__1587__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__461__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3842__ (
    .D(__1461__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__462__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3843__ (
    .D(__3108__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__463__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3844__ (
    .D(__193__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__464__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3845__ (
    .D(__2672__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__465__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3846__ (
    .D(__294__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__466__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3847__ (
    .D(__1952__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__467__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3848__ (
    .D(__1836__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__468__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3849__ (
    .D(__1447__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__469__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3850__ (
    .D(__1811__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__470__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3851__ (
    .D(__3134__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__471__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3852__ (
    .D(__2109__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__472__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3853__ (
    .D(__701__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__473__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3854__ (
    .D(__379__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__474__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3855__ (
    .D(__3229__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__475__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3856__ (
    .D(__2956__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__476__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3857__ (
    .D(__2995__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__477__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3858__ (
    .D(__2720__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__478__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3859__ (
    .D(__1758__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__479__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3860__ (
    .D(__2432__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__480__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3861__ (
    .D(__2403__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__481__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3862__ (
    .D(__2491__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__482__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3863__ (
    .D(__2488__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__483__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3864__ (
    .D(__2359__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__484__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3865__ (
    .D(__1103__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__485__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3866__ (
    .D(__2822__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__486__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3867__ (
    .D(__2364__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__487__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3868__ (
    .D(__2999__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__488__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3869__ (
    .D(__1603__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__489__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3870__ (
    .D(__1645__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__490__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3871__ (
    .D(__1938__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__491__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3872__ (
    .D(__3223__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__492__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3873__ (
    .D(__2640__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__493__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3874__ (
    .D(__3245__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__494__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3875__ (
    .D(__3377__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__495__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3876__ (
    .D(__2405__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__496__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3877__ (
    .D(__1809__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__497__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3878__ (
    .D(__3231__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__498__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3879__ (
    .D(__1578__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__499__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3880__ (
    .D(__3215__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__500__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3881__ (
    .D(__3191__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__501__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3882__ (
    .D(__1657__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__502__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3883__ (
    .D(__2021__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__503__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3884__ (
    .D(__3260__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__504__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3885__ (
    .D(__2154__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__505__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3886__ (
    .D(__1799__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__506__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3887__ (
    .D(__3293__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__507__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3888__ (
    .D(__3362__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__508__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3889__ (
    .D(__1458__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__509__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3890__ (
    .D(__3292__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__510__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3891__ (
    .D(__2759__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__511__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3892__ (
    .D(__2492__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__512__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3893__ (
    .D(__2549__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__513__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3894__ (
    .D(__2168__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__514__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3895__ (
    .D(__1292__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__515__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3896__ (
    .D(__1655__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__516__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3897__ (
    .D(__3048__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__517__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3898__ (
    .D(__901__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__518__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3899__ (
    .D(__3183__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__519__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3900__ (
    .D(__450__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__520__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3901__ (
    .D(__1157__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__521__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3902__ (
    .D(__2913__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__522__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3903__ (
    .D(__3189__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__523__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3904__ (
    .D(__3213__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__524__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3905__ (
    .D(__3271__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__525__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3906__ (
    .D(__1112__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__526__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3907__ (
    .D(__3113__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__527__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3908__ (
    .D(__330__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__528__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3909__ (
    .D(__2374__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__529__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3910__ (
    .D(__771__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__530__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3911__ (
    .D(__3198__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__531__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3912__ (
    .D(__3007__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__532__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3913__ (
    .D(__2545__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__533__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3914__ (
    .D(__2707__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__534__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3915__ (
    .D(__2213__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__535__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3916__ (
    .D(__654__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__536__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3917__ (
    .D(__1593__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__537__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3918__ (
    .D(__528__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__538__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3919__ (
    .D(__3079__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__539__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3920__ (
    .D(__3289__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__540__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3921__ (
    .D(__2951__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__541__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3922__ (
    .D(__3279__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__542__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3923__ (
    .D(__2923__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__543__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3924__ (
    .D(__709__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__544__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3925__ (
    .D(__2847__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__545__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3926__ (
    .D(__3275__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__546__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3927__ (
    .D(__2160__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__547__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3928__ (
    .D(__1683__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__548__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3929__ (
    .D(__2821__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__549__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3930__ (
    .D(__3208__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__550__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3931__ (
    .D(__3206__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__551__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3932__ (
    .D(__1565__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__552__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3933__ (
    .D(__2596__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__553__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3934__ (
    .D(__2433__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__554__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3935__ (
    .D(__1833__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__555__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3936__ (
    .D(__1634__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__556__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3937__ (
    .D(__2205__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__557__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3938__ (
    .D(__3036__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__558__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3939__ (
    .D(__2580__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__559__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3940__ (
    .D(__2011__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__560__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3941__ (
    .D(__1895__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__561__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3942__ (
    .D(__3112__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__562__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3943__ (
    .D(__1305__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__563__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3944__ (
    .D(__2588__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__564__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3945__ (
    .D(__2961__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__565__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3946__ (
    .D(__2043__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__566__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3947__ (
    .D(__2888__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__567__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3948__ (
    .D(__2681__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__568__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3949__ (
    .D(__3290__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__569__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3950__ (
    .D(__2379__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__570__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3951__ (
    .D(__1585__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__571__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3952__ (
    .D(__3165__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__572__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3953__ (
    .D(__217__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__573__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3954__ (
    .D(__1395__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__574__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3955__ (
    .D(__2845__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__575__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3956__ (
    .D(__3210__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__576__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3957__ (
    .D(__2247__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__577__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3958__ (
    .D(__2713__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__578__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3959__ (
    .D(__2583__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__579__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3960__ (
    .D(__1085__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__580__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3961__ (
    .D(__2476__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__581__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3962__ (
    .D(__1433__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__582__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3963__ (
    .D(__1884__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__583__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3964__ (
    .D(__3133__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__584__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3965__ (
    .D(__2505__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__585__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3966__ (
    .D(__128__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__586__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3967__ (
    .D(__2804__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__587__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3968__ (
    .D(__3218__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__588__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3969__ (
    .D(__2726__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__589__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3970__ (
    .D(__2803__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__590__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3971__ (
    .D(__1464__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__591__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3972__ (
    .D(__3120__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__592__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3973__ (
    .D(__1762__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__593__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3974__ (
    .D(__2617__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__594__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3975__ (
    .D(__2658__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__595__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3976__ (
    .D(__2674__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__596__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3977__ (
    .D(__2276__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__597__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3978__ (
    .D(__3107__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__598__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3979__ (
    .D(__1588__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__599__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3980__ (
    .D(__1202__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__600__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3981__ (
    .D(__2383__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__601__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3982__ (
    .D(__2757__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__602__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3983__ (
    .D(__1297__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__603__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3984__ (
    .D(__2494__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__604__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3985__ (
    .D(__2214__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__605__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3986__ (
    .D(__2039__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__606__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3987__ (
    .D(__3194__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__607__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3988__ (
    .D(__3225__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__608__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3989__ (
    .D(__2798__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__609__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3990__ (
    .D(__3020__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__610__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3991__ (
    .D(__2381__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__611__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3992__ (
    .D(__1335__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__612__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3993__ (
    .D(__1741__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__613__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3994__ (
    .D(__2342__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__614__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3995__ (
    .D(__1622__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__615__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3996__ (
    .D(__2352__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__616__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3997__ (
    .D(__2904__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__617__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3998__ (
    .D(__3186__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__618__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __3999__ (
    .D(__2974__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__619__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4000__ (
    .D(__2819__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__620__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4001__ (
    .D(__3024__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__621__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4002__ (
    .D(__1654__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__622__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4003__ (
    .D(__3142__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__623__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4004__ (
    .D(__2677__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__624__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4005__ (
    .D(__2539__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__625__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4006__ (
    .D(__1935__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__626__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4007__ (
    .D(__3163__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__627__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4008__ (
    .D(__2649__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__628__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4009__ (
    .D(__2007__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__629__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4010__ (
    .D(__2666__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__630__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4011__ (
    .D(__580__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__631__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4012__ (
    .D(__2712__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__632__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4013__ (
    .D(__3157__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__633__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4014__ (
    .D(__1626__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__634__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4015__ (
    .D(__30__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__635__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4016__ (
    .D(__1448__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__636__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4017__ (
    .D(__3371__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__637__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4018__ (
    .D(__2721__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__638__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4019__ (
    .D(__2519__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__639__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4020__ (
    .D(__3104__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__640__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4021__ (
    .D(__2457__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__641__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4022__ (
    .D(__1941__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__642__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4023__ (
    .D(__2509__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__643__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4024__ (
    .D(__723__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__644__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4025__ (
    .D(__2754__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__645__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4026__ (
    .D(__802__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__646__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4027__ (
    .D(__3149__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__647__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4028__ (
    .D(__2412__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__648__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4029__ (
    .D(__3326__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__649__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4030__ (
    .D(__85__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__650__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4031__ (
    .D(__3101__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__651__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4032__ (
    .D(__1855__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__652__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4033__ (
    .D(__1955__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__653__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4034__ (
    .D(__1135__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__654__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4035__ (
    .D(__2312__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__655__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4036__ (
    .D(__2638__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__656__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4037__ (
    .D(__3357__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__657__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4038__ (
    .D(__2752__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__658__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4039__ (
    .D(__2916__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__659__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4040__ (
    .D(__2619__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__660__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4041__ (
    .D(__442__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__661__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4042__ (
    .D(__3093__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__662__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4043__ (
    .D(__2919__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__663__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4044__ (
    .D(__3248__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__664__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4045__ (
    .D(__2167__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__665__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4046__ (
    .D(__2520__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__666__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4047__ (
    .D(__1333__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__667__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4048__ (
    .D(__1557__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__668__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4049__ (
    .D(__1606__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__669__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4050__ (
    .D(__3016__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__670__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4051__ (
    .D(__2326__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__671__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4052__ (
    .D(__2171__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__672__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4053__ (
    .D(__1748__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__673__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4054__ (
    .D(__1893__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__674__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4055__ (
    .D(__1350__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__675__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4056__ (
    .D(__2743__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__676__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4057__ (
    .D(__3247__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__677__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4058__ (
    .D(__3370__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__678__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4059__ (
    .D(__2885__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__679__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4060__ (
    .D(__1370__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__680__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4061__ (
    .D(__105__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__681__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4062__ (
    .D(__1435__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__682__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4063__ (
    .D(__867__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__683__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4064__ (
    .D(__1063__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__684__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4065__ (
    .D(__967__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__685__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4066__ (
    .D(__1729__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__686__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4067__ (
    .D(__2609__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__687__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4068__ (
    .D(__3274__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__688__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4069__ (
    .D(__2929__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__689__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4070__ (
    .D(__2315__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__690__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4071__ (
    .D(__3061__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__691__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4072__ (
    .D(__3184__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__692__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4073__ (
    .D(__1820__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__693__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4074__ (
    .D(__2924__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__694__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4075__ (
    .D(__3129__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__695__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4076__ (
    .D(__1339__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__696__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4077__ (
    .D(__3315__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__697__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4078__ (
    .D(__3076__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__698__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4079__ (
    .D(__3098__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__699__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4080__ (
    .D(__2334__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__700__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4081__ (
    .D(__2892__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__701__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4082__ (
    .D(__3168__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__702__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4083__ (
    .D(__2010__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__703__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4084__ (
    .D(__2814__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__704__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4085__ (
    .D(__2917__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__705__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4086__ (
    .D(__2413__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__706__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4087__ (
    .D(__117__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__707__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4088__ (
    .D(__2323__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__708__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4089__ (
    .D(__321__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__709__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4090__ (
    .D(__2261__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__710__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4091__ (
    .D(__2689__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__711__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4092__ (
    .D(__3052__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__712__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4093__ (
    .D(__2174__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__713__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4094__ (
    .D(__2306__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__714__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4095__ (
    .D(__2161__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__715__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4096__ (
    .D(__2813__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__716__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4097__ (
    .D(__2986__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__717__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4098__ (
    .D(__2898__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__718__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4099__ (
    .D(__3311__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__719__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4100__ (
    .D(__2124__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__720__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4101__ (
    .D(__2014__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__721__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4102__ (
    .D(__3075__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__722__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4103__ (
    .D(__518__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__723__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4104__ (
    .D(__474__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__724__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4105__ (
    .D(__3226__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__725__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4106__ (
    .D(__2928__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__726__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4107__ (
    .D(__2972__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__727__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4108__ (
    .D(__1984__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__728__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4109__ (
    .D(__2994__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__729__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4110__ (
    .D(__2360__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__730__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4111__ (
    .D(__3148__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__731__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4112__ (
    .D(__2933__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__732__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4113__ (
    .D(__3252__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__733__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4114__ (
    .D(__2750__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__734__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4115__ (
    .D(__2164__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__735__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4116__ (
    .D(__1177__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__736__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4117__ (
    .D(__3015__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__737__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4118__ (
    .D(__2408__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__738__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4119__ (
    .D(__214__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__739__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4120__ (
    .D(__2177__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__740__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4121__ (
    .D(__3009__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__741__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4122__ (
    .D(__2991__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__742__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4123__ (
    .D(__2576__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__743__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4124__ (
    .D(__3087__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__744__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4125__ (
    .D(__1644__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__745__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4126__ (
    .D(__2602__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__746__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4127__ (
    .D(__3146__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__747__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4128__ (
    .D(__2430__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__748__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4129__ (
    .D(__2508__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__749__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4130__ (
    .D(__3059__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__750__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4131__ (
    .D(__350__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__751__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4132__ (
    .D(__665__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__752__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4133__ (
    .D(__2330__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__753__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4134__ (
    .D(__1868__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__754__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4135__ (
    .D(__1482__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__755__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4136__ (
    .D(__1771__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__756__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4137__ (
    .D(__2670__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__757__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4138__ (
    .D(__3254__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__758__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4139__ (
    .D(__724__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__759__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4140__ (
    .D(__1711__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__760__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4141__ (
    .D(__1815__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__761__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4142__ (
    .D(__547__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__762__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4143__ (
    .D(__3217__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__763__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4144__ (
    .D(__2219__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__764__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4145__ (
    .D(__2654__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__765__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4146__ (
    .D(__2801__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__766__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4147__ (
    .D(__3038__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__767__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4148__ (
    .D(__1147__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__768__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4149__ (
    .D(__2440__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__769__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4150__ (
    .D(__2823__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__770__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4151__ (
    .D(__1225__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__771__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4152__ (
    .D(__14__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__772__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4153__ (
    .D(__1496__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__773__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4154__ (
    .D(__1038__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__774__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4155__ (
    .D(__2772__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__775__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4156__ (
    .D(__1945__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__776__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4157__ (
    .D(__2066__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__777__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4158__ (
    .D(__2426__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__778__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4159__ (
    .D(__2002__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__779__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4160__ (
    .D(__2968__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__780__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4161__ (
    .D(__3116__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__781__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4162__ (
    .D(__1418__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__782__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4163__ (
    .D(__2610__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__783__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4164__ (
    .D(__1583__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__784__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4165__ (
    .D(__1138__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__785__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4166__ (
    .D(__3283__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__786__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4167__ (
    .D(__1845__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__787__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4168__ (
    .D(__1858__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__788__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4169__ (
    .D(__2063__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__789__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4170__ (
    .D(__2572__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__790__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4171__ (
    .D(__2272__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__791__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4172__ (
    .D(__3170__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__792__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4173__ (
    .D(__3155__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__793__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4174__ (
    .D(__2613__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__794__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4175__ (
    .D(__2802__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__795__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4176__ (
    .D(__1745__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__796__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4177__ (
    .D(__2691__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__797__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4178__ (
    .D(__3152__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__798__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4179__ (
    .D(__2887__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__799__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4180__ (
    .D(__2513__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__800__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4181__ (
    .D(__3374__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__801__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4182__ (
    .D(__364__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__802__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4183__ (
    .D(__1736__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__803__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4184__ (
    .D(__2934__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__804__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4185__ (
    .D(__1613__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__805__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4186__ (
    .D(__2166__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__806__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4187__ (
    .D(__2639__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__807__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4188__ (
    .D(__2418__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__808__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4189__ (
    .D(__3102__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__809__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4190__ (
    .D(__3233__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__810__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4191__ (
    .D(__1216__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__811__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4192__ (
    .D(__2497__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__812__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4193__ (
    .D(__305__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__813__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4194__ (
    .D(__3032__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__814__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4195__ (
    .D(__49__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__815__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4196__ (
    .D(__3123__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__816__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4197__ (
    .D(__2872__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__817__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4198__ (
    .D(__2511__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__818__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4199__ (
    .D(__1287__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__819__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4200__ (
    .D(__2920__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__820__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4201__ (
    .D(__2571__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__821__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4202__ (
    .D(__2349__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__822__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4203__ (
    .D(__2595__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__823__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4204__ (
    .D(__2982__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__824__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4205__ (
    .D(__2109__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__825__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4206__ (
    .D(__3176__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__826__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4207__ (
    .D(__2185__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__827__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4208__ (
    .D(__1475__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__828__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4209__ (
    .D(__2253__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__829__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4210__ (
    .D(__2698__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__830__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4211__ (
    .D(__1526__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__831__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4212__ (
    .D(__1774__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__832__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4213__ (
    .D(__187__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__833__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4214__ (
    .D(__2341__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__834__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4215__ (
    .D(__2486__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__835__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4216__ (
    .D(__3306__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__836__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4217__ (
    .D(__3092__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__837__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4218__ (
    .D(__3205__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__838__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4219__ (
    .D(__1735__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__839__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4220__ (
    .D(__2013__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__840__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4221__ (
    .D(__3158__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__841__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4222__ (
    .D(__1614__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__842__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4223__ (
    .D(__2389__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__843__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4224__ (
    .D(__2612__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__844__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4225__ (
    .D(__3314__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__845__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4226__ (
    .D(__1971__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__846__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4227__ (
    .D(__1595__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__847__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4228__ (
    .D(__624__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__848__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4229__ (
    .D(__1713__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__849__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4230__ (
    .D(__1706__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__850__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4231__ (
    .D(__2313__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__851__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4232__ (
    .D(__3234__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__852__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4233__ (
    .D(__1947__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__853__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4234__ (
    .D(__2882__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__854__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4235__ (
    .D(__1850__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__855__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4236__ (
    .D(__1716__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__856__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4237__ (
    .D(__1184__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__857__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4238__ (
    .D(__2375__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__858__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4239__ (
    .D(__2900__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__859__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4240__ (
    .D(__2515__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__860__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4241__ (
    .D(__2936__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__861__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4242__ (
    .D(__3267__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__862__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4243__ (
    .D(__2962__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__863__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4244__ (
    .D(__1752__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__864__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4245__ (
    .D(__2667__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__865__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4246__ (
    .D(__1291__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__866__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4247__ (
    .D(__2510__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__867__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4248__ (
    .D(__2947__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__868__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4249__ (
    .D(__751__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__869__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4250__ (
    .D(__3185__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__870__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4251__ (
    .D(__3321__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__871__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4252__ (
    .D(__2976__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__872__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4253__ (
    .D(__394__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__873__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4254__ (
    .D(__1967__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__874__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4255__ (
    .D(__1515__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__875__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4256__ (
    .D(__2121__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__876__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4257__ (
    .D(__1846__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__877__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4258__ (
    .D(__1009__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__878__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4259__ (
    .D(__2265__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__879__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4260__ (
    .D(__1749__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__880__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4261__ (
    .D(__1402__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__881__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4262__ (
    .D(__1341__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__882__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4263__ (
    .D(__2767__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__883__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4264__ (
    .D(__2775__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__884__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4265__ (
    .D(__181__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__885__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4266__ (
    .D(__1352__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__886__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4267__ (
    .D(__263__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__887__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4268__ (
    .D(__3159__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__888__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4269__ (
    .D(__2827__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__889__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4270__ (
    .D(__2815__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__890__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4271__ (
    .D(__3028__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__891__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4272__ (
    .D(__2700__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__892__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4273__ (
    .D(__2980__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__893__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4274__ (
    .D(__2824__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__894__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4275__ (
    .D(__2964__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__895__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4276__ (
    .D(__1977__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__896__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4277__ (
    .D(__2846__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__897__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4278__ (
    .D(__2724__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__898__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4279__ (
    .D(__1529__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__899__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4280__ (
    .D(__2709__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__900__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4281__ (
    .D(__68__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__901__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4282__ (
    .D(__2569__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__902__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4283__ (
    .D(__3341__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__903__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4284__ (
    .D(__3089__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__904__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4285__ (
    .D(__2950__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__905__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4286__ (
    .D(__2593__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__906__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4287__ (
    .D(__3338__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__907__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4288__ (
    .D(__1783__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__908__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4289__ (
    .D(__2668__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__909__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4290__ (
    .D(__2151__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__910__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4291__ (
    .D(__1744__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__911__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4292__ (
    .D(__66__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__912__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4293__ (
    .D(__1978__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__913__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4294__ (
    .D(__2050__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__914__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4295__ (
    .D(__2761__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__915__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4296__ (
    .D(__3286__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__916__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4297__ (
    .D(__1992__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__917__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4298__ (
    .D(__2344__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__918__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4299__ (
    .D(__2378__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__919__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4300__ (
    .D(__72__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__920__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4301__ (
    .D(__3073__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__921__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4302__ (
    .D(__2660__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__922__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4303__ (
    .D(__1889__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__923__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4304__ (
    .D(__2881__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__924__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4305__ (
    .D(__1301__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__925__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4306__ (
    .D(__2579__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__926__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4307__ (
    .D(__2321__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__927__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4308__ (
    .D(__2386__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__928__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4309__ (
    .D(__1970__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__929__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4310__ (
    .D(__2417__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__930__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4311__ (
    .D(__1826__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__931__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4312__ (
    .D(__2437__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__932__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4313__ (
    .D(__3287__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__933__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4314__ (
    .D(__2811__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__934__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4315__ (
    .D(__302__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__935__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4316__ (
    .D(__2400__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__936__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4317__ (
    .D(__2047__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__937__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4318__ (
    .D(__1822__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__938__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4319__ (
    .D(__3154__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__939__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4320__ (
    .D(__924__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__940__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4321__ (
    .D(__1986__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__941__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4322__ (
    .D(__3310__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__942__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4323__ (
    .D(__1760__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__943__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4324__ (
    .D(__2880__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__944__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4325__ (
    .D(__1272__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__945__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4326__ (
    .D(__3284__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__946__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4327__ (
    .D(__1831__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__947__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4328__ (
    .D(__2159__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__948__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4329__ (
    .D(__2656__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__949__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4330__ (
    .D(__2279__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__950__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4331__ (
    .D(__2240__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__951__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4332__ (
    .D(__3137__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__952__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4333__ (
    .D(__2028__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__953__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4334__ (
    .D(__2651__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__954__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4335__ (
    .D(__2493__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__955__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4336__ (
    .D(__712__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__956__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4337__ (
    .D(__2354__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__957__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4338__ (
    .D(__2600__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__958__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4339__ (
    .D(__3012__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__959__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4340__ (
    .D(__2538__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__960__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4341__ (
    .D(__2883__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__961__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4342__ (
    .D(__3269__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__962__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4343__ (
    .D(__2719__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__963__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4344__ (
    .D(__2939__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__964__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4345__ (
    .D(__2932__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__965__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4346__ (
    .D(__3261__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__966__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4347__ (
    .D(__2996__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__967__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4348__ (
    .D(__2333__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__968__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4349__ (
    .D(__2597__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__969__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4350__ (
    .D(__2467__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__970__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4351__ (
    .D(__3295__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__971__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4352__ (
    .D(__1825__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__972__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4353__ (
    .D(__28__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__973__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4354__ (
    .D(__2860__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__974__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4355__ (
    .D(__2336__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__975__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4356__ (
    .D(__3343__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__976__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4357__ (
    .D(__2449__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__977__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4358__ (
    .D(__2646__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__978__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4359__ (
    .D(__359__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__979__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4360__ (
    .D(__1951__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__980__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4361__ (
    .D(__2394__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__981__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4362__ (
    .D(__2977__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__982__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4363__ (
    .D(__2694__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__983__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4364__ (
    .D(__2946__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__984__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4365__ (
    .D(__3301__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__985__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4366__ (
    .D(__2902__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__986__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4367__ (
    .D(__1937__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__987__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4368__ (
    .D(__3126__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__988__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4369__ (
    .D(__1387__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__989__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4370__ (
    .D(__287__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__990__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4371__ (
    .D(__349__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__991__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4372__ (
    .D(__2425__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__992__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4373__ (
    .D(__3319__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__993__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4374__ (
    .D(__80__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__994__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4375__ (
    .D(__1518__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__995__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4376__ (
    .D(__1856__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__996__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4377__ (
    .D(__1664__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__997__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4378__ (
    .D(__380__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__998__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4379__ (
    .D(__2817__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__999__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4380__ (
    .D(__2259__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1000__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4381__ (
    .D(__2018__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1001__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4382__ (
    .D(__2424__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1002__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4383__ (
    .D(__3375__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1003__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4384__ (
    .D(__2816__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1004__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4385__ (
    .D(__230__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1005__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4386__ (
    .D(__644__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1006__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4387__ (
    .D(__1559__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1007__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4388__ (
    .D(__2963__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1008__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4389__ (
    .D(__168__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1009__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4390__ (
    .D(__3266__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1010__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4391__ (
    .D(__2918__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1011__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4392__ (
    .D(__1340__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1012__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4393__ (
    .D(__1478__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1013__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4394__ (
    .D(__2216__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1014__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4395__ (
    .D(__2760__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1015__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4396__ (
    .D(__1384__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1016__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4397__ (
    .D(__1628__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1017__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4398__ (
    .D(__3065__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1018__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4399__ (
    .D(__1731__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1019__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4400__ (
    .D(__2675__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1020__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4401__ (
    .D(__1888__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1021__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4402__ (
    .D(__1544__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1022__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4403__ (
    .D(__2250__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1023__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4404__ (
    .D(__2734__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1024__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4405__ (
    .D(__1509__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1025__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4406__ (
    .D(__1739__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1026__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4407__ (
    .D(__2490__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1027__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4408__ (
    .D(__3212__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1028__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4409__ (
    .D(__2895__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1029__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4410__ (
    .D(__3175__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1030__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4411__ (
    .D(__2404__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1031__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4412__ (
    .D(__3298__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1032__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4413__ (
    .D(__1195__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1033__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4414__ (
    .D(__2274__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1034__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4415__ (
    .D(__3136__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1035__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4416__ (
    .D(__1814__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1036__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4417__ (
    .D(__3329__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1037__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4418__ (
    .D(__1217__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1038__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4419__ (
    .D(__2015__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1039__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4420__ (
    .D(__3304__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1040__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4421__ (
    .D(__3027__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1041__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4422__ (
    .D(__3280__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1042__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4423__ (
    .D(__3325__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1043__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4424__ (
    .D(__3131__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1044__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4425__ (
    .D(__3078__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1045__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4426__ (
    .D(__3296__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1046__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4427__ (
    .D(__3088__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1047__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4428__ (
    .D(__2665__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1048__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4429__ (
    .D(__2218__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1049__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4430__ (
    .D(__3161__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1050__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4431__ (
    .D(__2876__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1051__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4432__ (
    .D(__2862__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1052__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4433__ (
    .D(__2577__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1053__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4434__ (
    .D(__1998__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1054__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4435__ (
    .D(__990__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1055__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4436__ (
    .D(__2865__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1056__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4437__ (
    .D(__1434__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1057__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4438__ (
    .D(__1959__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1058__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4439__ (
    .D(__2905__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1059__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4440__ (
    .D(__1579__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1060__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4441__ (
    .D(__1740__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1061__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4442__ (
    .D(__2162__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1062__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4443__ (
    .D(__1123__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1063__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4444__ (
    .D(__2685__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1064__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4445__ (
    .D(__1617__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1065__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4446__ (
    .D(__1685__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1066__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4447__ (
    .D(__2192__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1067__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4448__ (
    .D(__2506__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1068__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4449__ (
    .D(__1005__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1069__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4450__ (
    .D(__3172__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1070__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4451__ (
    .D(__1543__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1071__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4452__ (
    .D(__1862__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1072__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4453__ (
    .D(__1392__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1073__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4454__ (
    .D(__351__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1074__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4455__ (
    .D(__2540__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1075__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4456__ (
    .D(__3238__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1076__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4457__ (
    .D(__2959__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1077__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4458__ (
    .D(__3118__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1078__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4459__ (
    .D(__3063__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1079__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4460__ (
    .D(__2586__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1080__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4461__ (
    .D(__3220__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1081__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4462__ (
    .D(__3121__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1082__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4463__ (
    .D(__2879__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1083__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4464__ (
    .D(__1944__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1084__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4465__ (
    .D(__3130__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1085__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4466__ (
    .D(__1863__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1086__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4467__ (
    .D(__256__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1087__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4468__ (
    .D(__2186__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1088__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4469__ (
    .D(__3179__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1089__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4470__ (
    .D(__2943__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1090__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4471__ (
    .D(__3379__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1091__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4472__ (
    .D(__1492__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1092__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4473__ (
    .D(__2466__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1093__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4474__ (
    .D(__1431__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1094__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4475__ (
    .D(__1772__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1095__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4476__ (
    .D(__2840__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1096__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4477__ (
    .D(__215__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1097__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4478__ (
    .D(__1623__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1098__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4479__ (
    .D(__3291__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1099__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4480__ (
    .D(__2096__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1100__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4481__ (
    .D(__1999__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1101__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4482__ (
    .D(__813__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1102__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4483__ (
    .D(__1755__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1103__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4484__ (
    .D(__2338__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1104__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4485__ (
    .D(__3106__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1105__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4486__ (
    .D(__559__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1106__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4487__ (
    .D(__2151__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1107__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4488__ (
    .D(__2455__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1108__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4489__ (
    .D(__1994__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1109__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4490__ (
    .D(__2701__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1110__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4491__ (
    .D(__2278__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1111__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4492__ (
    .D(__2429__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1112__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4493__ (
    .D(__2271__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1113__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4494__ (
    .D(__2269__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1114__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4495__ (
    .D(__1976__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1115__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4496__ (
    .D(__2203__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1116__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4497__ (
    .D(__2768__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1117__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4498__ (
    .D(__2776__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1118__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4499__ (
    .D(__2901__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1119__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4500__ (
    .D(__2544__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1120__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4501__ (
    .D(__1737__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1121__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4502__ (
    .D(__2388__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1122__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4503__ (
    .D(__1074__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1123__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4504__ (
    .D(__3364__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1124__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4505__ (
    .D(__2730__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1125__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4506__ (
    .D(__2303__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1126__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4507__ (
    .D(__2438__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1127__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4508__ (
    .D(__3361__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1128__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4509__ (
    .D(__2915__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1129__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4510__ (
    .D(__2903__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1130__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4511__ (
    .D(__2460__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1131__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4512__ (
    .D(__3246__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1132__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4513__ (
    .D(__1686__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1133__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4514__ (
    .D(__1972__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1134__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4515__ (
    .D(__811__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1135__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4516__ (
    .D(__3084__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1136__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4517__ (
    .D(__3005__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1137__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4518__ (
    .D(__1690__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1138__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4519__ (
    .D(__2337__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1139__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4520__ (
    .D(__3358__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1140__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4521__ (
    .D(__3353__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1141__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4522__ (
    .D(__2245__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1142__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4523__ (
    .D(__2997__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1143__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4524__ (
    .D(__2464__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1144__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4525__ (
    .D(__2941__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1145__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4526__ (
    .D(__1500__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1146__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4527__ (
    .D(__1511__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1147__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4528__ (
    .D(__2206__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1148__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4529__ (
    .D(__2485__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1149__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4530__ (
    .D(__2989__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1150__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4531__ (
    .D(__2062__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1151__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4532__ (
    .D(__1769__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1152__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4533__ (
    .D(__2828__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1153__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4534__ (
    .D(__2444__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1154__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4535__ (
    .D(__3033__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1155__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4536__ (
    .D(__3110__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1156__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4537__ (
    .D(__554__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1157__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4538__ (
    .D(__2575__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1158__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4539__ (
    .D(__3327__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1159__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4540__ (
    .D(__2874__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1160__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4541__ (
    .D(__2507__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1161__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4542__ (
    .D(__935__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1162__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4543__ (
    .D(__1838__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1163__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4544__ (
    .D(__3224__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1164__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4545__ (
    .D(__2645__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1165__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4546__ (
    .D(__3135__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1166__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4547__ (
    .D(__2671__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1167__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4548__ (
    .D(__3056__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1168__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4549__ (
    .D(__520__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1169__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4550__ (
    .D(__3193__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1170__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4551__ (
    .D(__3004__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1171__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4552__ (
    .D(__1222__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1172__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4553__ (
    .D(__2169__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1173__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4554__ (
    .D(__1939__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1174__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4555__ (
    .D(__3066__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1175__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4556__ (
    .D(__2305__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1176__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4557__ (
    .D(__170__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1177__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4558__ (
    .D(__3045__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1178__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4559__ (
    .D(__1610__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1179__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4560__ (
    .D(__1439__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1180__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4561__ (
    .D(__1768__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1181__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4562__ (
    .D(__1527__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1182__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4563__ (
    .D(__3181__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1183__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4564__ (
    .D(__3022__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1184__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4565__ (
    .D(__1661__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1185__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4566__ (
    .D(__2328__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1186__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4567__ (
    .D(__1886__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1187__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4568__ (
    .D(__2139__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1188__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4569__ (
    .D(__2397__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1189__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4570__ (
    .D(__3119__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1190__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4571__ (
    .D(__2049__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1191__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4572__ (
    .D(__1442__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1192__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4573__ (
    .D(__2869__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1193__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4574__ (
    .D(__2680__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1194__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4575__ (
    .D(__3006__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1195__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4576__ (
    .D(__3153__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1196__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4577__ (
    .D(__2471__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1197__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4578__ (
    .D(__1659__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1198__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4579__ (
    .D(__823__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1199__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4580__ (
    .D(__2181__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1200__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4581__ (
    .D(__1668__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1201__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4582__ (
    .D(__169__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1202__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4583__ (
    .D(__2981__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1203__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4584__ (
    .D(__2812__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1204__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4585__ (
    .D(__1682__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1205__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4586__ (
    .D(__2975__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1206__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4587__ (
    .D(__1547__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1207__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4588__ (
    .D(__2542__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1208__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4589__ (
    .D(__1987__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1209__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4590__ (
    .D(__1916__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1210__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4591__ (
    .D(__1679__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1211__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4592__ (
    .D(__1507__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1212__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4593__ (
    .D(__2248__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1213__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4594__ (
    .D(__3051__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1214__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4595__ (
    .D(__2468__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1215__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4596__ (
    .D(__833__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1216__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4597__ (
    .D(__1162__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1217__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4598__ (
    .D(__3288__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1218__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4599__ (
    .D(__1494__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1219__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4600__ (
    .D(__2201__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1220__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4601__ (
    .D(__3334__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1221__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4602__ (
    .D(__366__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1222__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4603__ (
    .D(__3342__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1223__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4604__ (
    .D(__2682__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1224__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4605__ (
    .D(__2514__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1225__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4606__ (
    .D(__3256__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1226__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4607__ (
    .D(__3144__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1227__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4608__ (
    .D(__2355__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1228__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4609__ (
    .D(__1881__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1229__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4610__ (
    .D(__1990__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1230__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4611__ (
    .D(__2992__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1231__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4612__ (
    .D(__3086__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1232__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4613__ (
    .D(__2022__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1233__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4614__ (
    .D(__2300__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1234__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4615__ (
    .D(__3262__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1235__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4616__ (
    .D(__2446__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1236__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4617__ (
    .D(__1709__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1237__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4618__ (
    .D(__2410__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1238__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4619__ (
    .D(__2844__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1239__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4620__ (
    .D(__1777__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1240__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4621__ (
    .D(__2322__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1241__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4622__ (
    .D(__3070__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1242__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4623__ (
    .D(__3356__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1243__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4624__ (
    .D(__1861__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1244__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4625__ (
    .D(__3096__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1245__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4626__ (
    .D(__1854__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1246__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4627__ (
    .D(__3156__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1247__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4628__ (
    .D(__71__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1248__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4629__ (
    .D(__2157__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1249__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4630__ (
    .D(__2384__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1250__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4631__ (
    .D(__3250__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1251__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4632__ (
    .D(__3368__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1252__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4633__ (
    .D(__2969__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1253__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4634__ (
    .D(__106__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1254__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4635__ (
    .D(__2944__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1255__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4636__ (
    .D(__2777__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1256__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4637__ (
    .D(__3160__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1257__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4638__ (
    .D(__3211__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1258__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4639__ (
    .D(__1806__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1259__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4640__ (
    .D(__2978__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1260__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4641__ (
    .D(__1307__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1261__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4642__ (
    .D(__3372__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1262__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4643__ (
    .D(__1604__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1263__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4644__ (
    .D(__1658__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1264__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4645__ (
    .D(__2825__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1265__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4646__ (
    .D(__2482__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1266__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4647__ (
    .D(__3340__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1267__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4648__ (
    .D(__3251__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1268__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4649__ (
    .D(__3067__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1269__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4650__ (
    .D(__2239__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1270__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4651__ (
    .D(__2243__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1271__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4652__ (
    .D(__1102__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1272__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4653__ (
    .D(__2606__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1273__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4654__ (
    .D(__1957__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1274__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4655__ (
    .D(__3050__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1275__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4656__ (
    .D(__1502__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1276__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4657__ (
    .D(__2966__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1277__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4658__ (
    .D(__3232__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1278__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4659__ (
    .D(__2016__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1279__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4660__ (
    .D(__2855__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1280__)
  );
  LUT5 #(
    .INIT(32'h82000082)
  ) __4662__ (
    .I4(g72),
    .I3(__591__),
    .I2(g73),
    .I1(__851__),
    .I0(__353__),
    .O(__1282__)
  );
  LUT3 #(
    .INIT(8'h07)
  ) __4663__ (
    .I2(g134),
    .I1(__884__),
    .I0(g99),
    .O(__1283__)
  );
  LUT6 #(
    .INIT(64'h0000000000000008)
  ) __4664__ (
    .I5(__917__),
    .I4(__972__),
    .I3(g113),
    .I2(__1283__),
    .I1(__749__),
    .I0(__1282__),
    .O(__1284__)
  );
  LUT4 #(
    .INIT(16'h0004)
  ) __4665__ (
    .I3(__917__),
    .I2(__353__),
    .I1(__1227__),
    .I0(__972__),
    .O(__1285__)
  );
  LUT6 #(
    .INIT(64'h000000000000fff4)
  ) __4666__ (
    .I5(__795__),
    .I4(__718__),
    .I3(__465__),
    .I2(__842__),
    .I1(__1285__),
    .I0(__1000__),
    .O(__1286__)
  );
  LUT5 #(
    .INIT(32'hffa0cfc0)
  ) __4667__ (
    .I4(__1286__),
    .I3(__769__),
    .I2(g35),
    .I1(__819__),
    .I0(__1284__),
    .O(__1287__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __4669__ (
    .I1(__1027__),
    .I0(__296__),
    .O(__1289__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __4670__ (
    .I1(__819__),
    .I0(__982__),
    .O(__1290__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __4671__ (
    .I5(g35),
    .I4(__1286__),
    .I3(__1290__),
    .I2(__866__),
    .I1(__923__),
    .I0(__1289__),
    .O(__1291__)
  );
  LUT6 #(
    .INIT(64'hff00ccccf0f0aaaa)
  ) __4672__ (
    .I5(__282__),
    .I4(__132__),
    .I3(__125__),
    .I2(__409__),
    .I1(__374__),
    .I0(__1179__),
    .O(__1292__)
  );
  LUT5 #(
    .INIT(32'hccaaf0f0)
  ) __4673__ (
    .I4(g35),
    .I3(__364__),
    .I2(__1018__),
    .I1(__1263__),
    .I0(__293__),
    .O(__1293__)
  );
  LUT6 #(
    .INIT(64'h8000080020000200)
  ) __4674__ (
    .I5(g72),
    .I4(g73),
    .I3(__757__),
    .I2(__664__),
    .I1(__629__),
    .I0(__605__),
    .O(__1294__)
  );
  LUT5 #(
    .INIT(32'h00000008)
  ) __4675__ (
    .I4(g113),
    .I3(__1283__),
    .I2(__810__),
    .I1(__236__),
    .I0(__1294__),
    .O(__1295__)
  );
  LUT5 #(
    .INIT(32'h10ff0000)
  ) __4676__ (
    .I4(__636__),
    .I3(g35),
    .I2(__688__),
    .I1(__457__),
    .I0(__1295__),
    .O(__1296__)
  );
  LUT6 #(
    .INIT(64'hefefff00ff00ff00)
  ) __4677__ (
    .I5(g35),
    .I4(__341__),
    .I3(__393__),
    .I2(g73),
    .I1(g72),
    .I0(__1280__),
    .O(__1297__)
  );
  LUT6 #(
    .INIT(64'h8000080020000200)
  ) __4678__ (
    .I5(g72),
    .I4(g73),
    .I3(__917__),
    .I2(__851__),
    .I1(__591__),
    .I0(__353__),
    .O(__1298__)
  );
  LUT6 #(
    .INIT(64'h00000000fff40000)
  ) __4679__ (
    .I5(__718__),
    .I4(__795__),
    .I3(__465__),
    .I2(__842__),
    .I1(__1285__),
    .I0(__864__),
    .O(__1299__)
  );
  LUT5 #(
    .INIT(32'h00000008)
  ) __4680__ (
    .I4(__972__),
    .I3(g113),
    .I2(__1283__),
    .I1(__1299__),
    .I0(__1298__),
    .O(__1300__)
  );
  LUT6 #(
    .INIT(64'hf30caaaaf0f0f0f0)
  ) __4681__ (
    .I5(g35),
    .I4(__1300__),
    .I3(__749__),
    .I2(__760__),
    .I1(__541__),
    .I0(__925__),
    .O(__1301__)
  );
  LUT6 #(
    .INIT(64'h0000000082000082)
  ) __4682__ (
    .I5(__757__),
    .I4(g72),
    .I3(__629__),
    .I2(g73),
    .I1(__664__),
    .I0(__605__),
    .O(__1302__)
  );
  LUT5 #(
    .INIT(32'h0000f800)
  ) __4683__ (
    .I4(g113),
    .I3(__236__),
    .I2(g134),
    .I1(__884__),
    .I0(g99),
    .O(__1303__)
  );
  LUT6 #(
    .INIT(64'h00dfdf00ffff0000)
  ) __4684__ (
    .I5(g35),
    .I4(__798__),
    .I3(__386__),
    .I2(__1303__),
    .I1(__810__),
    .I0(__1302__),
    .O(__1304__)
  );
  LUT6 #(
    .INIT(64'ha0aaf0ffcccccccc)
  ) __4685__ (
    .I5(g35),
    .I4(__1249__),
    .I3(__973__),
    .I2(__279__),
    .I1(__1127__),
    .I0(__563__),
    .O(__1305__)
  );
  LUT4 #(
    .INIT(16'h8000)
  ) __4686__ (
    .I3(__187__),
    .I2(__103__),
    .I1(__823__),
    .I0(__1199__),
    .O(__1306__)
  );
  LUT4 #(
    .INIT(16'h7f00)
  ) __4687__ (
    .I3(__1044__),
    .I2(g35),
    .I1(__62__),
    .I0(__1306__),
    .O(__1307__)
  );
  LUT5 #(
    .INIT(32'h00cef0f0)
  ) __4688__ (
    .I4(g35),
    .I3(__43__),
    .I2(__683__),
    .I1(__158__),
    .I0(__867__),
    .O(__1308__)
  );
  LUT3 #(
    .INIT(8'h04)
  ) __4689__ (
    .I2(__288__),
    .I1(__788__),
    .I0(__721__),
    .O(__1309__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __4690__ (
    .I2(__926__),
    .I1(__995__),
    .I0(__1192__),
    .O(__1310__)
  );
  LUT6 #(
    .INIT(64'h7fffffff00000000)
  ) __4691__ (
    .I5(__151__),
    .I4(__1310__),
    .I3(__69__),
    .I2(__1077__),
    .I1(__1309__),
    .I0(__780__),
    .O(__1311__)
  );
  LUT5 #(
    .INIT(32'h80000000)
  ) __4692__ (
    .I4(__1311__),
    .I3(__557__),
    .I2(__696__),
    .I1(__897__),
    .I0(__661__),
    .O(__1312__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __4693__ (
    .I1(__557__),
    .I0(__696__),
    .O(__1313__)
  );
  LUT6 #(
    .INIT(64'h0fffffffffff7777)
  ) __4694__ (
    .I5(__557__),
    .I4(__696__),
    .I3(__160__),
    .I2(__24__),
    .I1(__442__),
    .I0(__1185__),
    .O(__1314__)
  );
  LUT6 #(
    .INIT(64'h7f00000000007f00)
  ) __4695__ (
    .I5(__897__),
    .I4(__502__),
    .I3(__1314__),
    .I2(__1313__),
    .I1(__45__),
    .I0(__1015__),
    .O(__1315__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __4696__ (
    .I1(__696__),
    .I0(__557__),
    .O(__1316__)
  );
  LUT6 #(
    .INIT(64'hffff0fffffff7777)
  ) __4697__ (
    .I5(__557__),
    .I4(__696__),
    .I3(__442__),
    .I2(__714__),
    .I1(__670__),
    .I0(__45__),
    .O(__1317__)
  );
  LUT6 #(
    .INIT(64'h00007f007f000000)
  ) __4698__ (
    .I5(__897__),
    .I4(__502__),
    .I3(__1317__),
    .I2(__1316__),
    .I1(__911__),
    .I0(__160__),
    .O(__1318__)
  );
  LUT4 #(
    .INIT(16'h8000)
  ) __4699__ (
    .I3(__557__),
    .I2(__696__),
    .I1(__897__),
    .I0(__661__),
    .O(__1319__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __4700__ (
    .I1(__557__),
    .I0(__696__),
    .O(__1320__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __4701__ (
    .I1(__517__),
    .I0(__215__),
    .O(__1321__)
  );
  LUT6 #(
    .INIT(64'h007f7f7f00000000)
  ) __4702__ (
    .I5(__897__),
    .I4(__1313__),
    .I3(__1321__),
    .I2(__1097__),
    .I1(__1320__),
    .I0(__615__),
    .O(__1322__)
  );
  LUT6 #(
    .INIT(64'h000000f800000088)
  ) __4703__ (
    .I5(__238__),
    .I4(__557__),
    .I3(__696__),
    .I2(__346__),
    .I1(__259__),
    .I0(__317__),
    .O(__1323__)
  );
  LUT6 #(
    .INIT(64'h000007770000ffff)
  ) __4704__ (
    .I5(__1316__),
    .I4(__1323__),
    .I3(__1214__),
    .I2(__502__),
    .I1(__272__),
    .I0(__433__),
    .O(__1324__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __4705__ (
    .I1(__557__),
    .I0(__696__),
    .O(__1325__)
  );
  LUT6 #(
    .INIT(64'h0000f88800000000)
  ) __4706__ (
    .I5(__557__),
    .I4(__696__),
    .I3(__1137__),
    .I2(__346__),
    .I1(__259__),
    .I0(__119__),
    .O(__1326__)
  );
  LUT6 #(
    .INIT(64'h0000f88800000000)
  ) __4707__ (
    .I5(__696__),
    .I4(__557__),
    .I3(__475__),
    .I2(__1097__),
    .I1(__458__),
    .I0(__661__),
    .O(__1327__)
  );
  LUT6 #(
    .INIT(64'h000007770000ffff)
  ) __4708__ (
    .I5(__1320__),
    .I4(__1327__),
    .I3(__487__),
    .I2(__433__),
    .I1(__421__),
    .I0(__502__),
    .O(__1328__)
  );
  LUT6 #(
    .INIT(64'h0000007f00000000)
  ) __4709__ (
    .I5(__1328__),
    .I4(__897__),
    .I3(__1326__),
    .I2(__1042__),
    .I1(__1325__),
    .I0(__215__),
    .O(__1329__)
  );
  LUT3 #(
    .INIT(8'h07)
  ) __4710__ (
    .I2(__1329__),
    .I1(__1324__),
    .I0(__1322__),
    .O(__1330__)
  );
  LUT6 #(
    .INIT(64'hfffff11100000000)
  ) __4711__ (
    .I5(__1311__),
    .I4(__1330__),
    .I3(__1319__),
    .I2(__831__),
    .I1(__1318__),
    .I0(__1315__),
    .O(__1331__)
  );
  LUT5 #(
    .INIT(32'hcf30aaaa)
  ) __4712__ (
    .I4(g35),
    .I3(__1331__),
    .I2(__361__),
    .I1(__1312__),
    .I0(__754__),
    .O(__1332__)
  );
  LUT5 #(
    .INIT(32'hf3ff8ccc)
  ) __4713__ (
    .I4(__1019__),
    .I3(__1085__),
    .I2(__214__),
    .I1(g35),
    .I0(__896__),
    .O(__1333__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __4714__ (
    .I1(__359__),
    .I0(__979__),
    .O(__1334__)
  );
  LUT6 #(
    .INIT(64'h0a03000000000000)
  ) __4715__ (
    .I5(g35),
    .I4(__1334__),
    .I3(__394__),
    .I2(__115__),
    .I1(__873__),
    .I0(__612__),
    .O(__1335__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __4716__ (
    .I1(__1052__),
    .I0(__1236__),
    .O(__1336__)
  );
  LUT6 #(
    .INIT(64'h8000080020000200)
  ) __4717__ (
    .I5(g72),
    .I4(g73),
    .I3(__1240__),
    .I2(__738__),
    .I1(__976__),
    .I0(__1336__),
    .O(__1337__)
  );
  LUT5 #(
    .INIT(32'h0000f800)
  ) __4718__ (
    .I4(g113),
    .I3(__499__),
    .I2(g134),
    .I1(__884__),
    .I0(g99),
    .O(__1338__)
  );
  LUT6 #(
    .INIT(64'h0077ff00f0f0f0f0)
  ) __4719__ (
    .I5(g35),
    .I4(__1311__),
    .I3(__696__),
    .I2(__18__),
    .I1(__1338__),
    .I0(__1337__),
    .O(__1339__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __4720__ (
    .I2(g35),
    .I1(__1012__),
    .I0(__1121__),
    .O(__1340__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __4721__ (
    .I2(g35),
    .I1(g6748),
    .I0(__530__),
    .O(__1341__)
  );
  LUT6 #(
    .INIT(64'h00000000cfdfffff)
  ) __4722__ (
    .I5(g134),
    .I4(__1115__),
    .I3(__35__),
    .I2(__1249__),
    .I1(__304__),
    .I0(__437__),
    .O(__1342__)
  );
  LUT6 #(
    .INIT(64'h0000f3ff00005155)
  ) __4723__ (
    .I5(__1118__),
    .I4(__1342__),
    .I3(__65__),
    .I2(__493__),
    .I1(__895__),
    .I0(__710__),
    .O(__1343__)
  );
  LUT6 #(
    .INIT(64'h88d8888888d888d8)
  ) __4724__ (
    .I5(__710__),
    .I4(__1118__),
    .I3(__1342__),
    .I2(__1248__),
    .I1(__739__),
    .I0(__1343__),
    .O(__1344__)
  );
  LUT6 #(
    .INIT(64'h0000000000000008)
  ) __4725__ (
    .I5(__992__),
    .I4(__952__),
    .I3(__206__),
    .I2(__423__),
    .I1(__1019__),
    .I0(__631__),
    .O(__1345__)
  );
  LUT4 #(
    .INIT(16'hbf00)
  ) __4726__ (
    .I3(__168__),
    .I2(__1345__),
    .I1(__881__),
    .I0(__660__),
    .O(__1346__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __4727__ (
    .I1(__710__),
    .I0(__1118__),
    .O(__1347__)
  );
  LUT6 #(
    .INIT(64'h00000000000000f7)
  ) __4728__ (
    .I5(__1347__),
    .I4(__1346__),
    .I3(__1342__),
    .I2(__493__),
    .I1(__65__),
    .I0(__895__),
    .O(__1348__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __4729__ (
    .I1(__728__),
    .I0(__1348__),
    .O(__1349__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __4730__ (
    .I5(g35),
    .I4(__801__),
    .I3(__1349__),
    .I2(__675__),
    .I1(__78__),
    .I0(__1344__),
    .O(__1350__)
  );
  LUT3 #(
    .INIT(8'hd0)
  ) __4731__ (
    .I2(__218__),
    .I1(__751__),
    .I0(__350__),
    .O(__1351__)
  );
  LUT6 #(
    .INIT(64'h23af8c00ff00ff00)
  ) __4732__ (
    .I5(g35),
    .I4(__886__),
    .I3(__185__),
    .I2(__751__),
    .I1(__1351__),
    .I0(__869__),
    .O(__1352__)
  );
  LUT5 #(
    .INIT(32'h00000080)
  ) __4733__ (
    .I4(__96__),
    .I3(__720__),
    .I2(__1100__),
    .I1(__876__),
    .I0(__825__),
    .O(__1353__)
  );
  LUT4 #(
    .INIT(16'h0080)
  ) __4734__ (
    .I3(__1107__),
    .I2(__50__),
    .I1(__118__),
    .I0(__1353__),
    .O(__1354__)
  );
  LUT5 #(
    .INIT(32'h00000008)
  ) __4735__ (
    .I4(__1100__),
    .I3(__876__),
    .I2(__825__),
    .I1(__96__),
    .I0(__720__),
    .O(__1355__)
  );
  LUT4 #(
    .INIT(16'h0008)
  ) __4736__ (
    .I3(__50__),
    .I2(__1107__),
    .I1(__118__),
    .I0(__1355__),
    .O(__1356__)
  );
  LUT5 #(
    .INIT(32'h00000004)
  ) __4737__ (
    .I4(__1100__),
    .I3(__876__),
    .I2(__720__),
    .I1(__96__),
    .I0(__825__),
    .O(__1357__)
  );
  LUT5 #(
    .INIT(32'h00000080)
  ) __4738__ (
    .I4(__50__),
    .I3(__1107__),
    .I2(__118__),
    .I1(__1357__),
    .I0(__1057__),
    .O(__1358__)
  );
  LUT5 #(
    .INIT(32'h00008000)
  ) __4739__ (
    .I4(__720__),
    .I3(__96__),
    .I2(__1100__),
    .I1(__876__),
    .I0(__825__),
    .O(__1359__)
  );
  LUT4 #(
    .INIT(16'h0080)
  ) __4740__ (
    .I3(__118__),
    .I2(__50__),
    .I1(__1107__),
    .I0(__1359__),
    .O(__1360__)
  );
  LUT6 #(
    .INIT(64'h0000000000000777)
  ) __4741__ (
    .I5(__1360__),
    .I4(__1358__),
    .I3(g100),
    .I2(__1356__),
    .I1(__505__),
    .I0(__1354__),
    .O(__1361__)
  );
  LUT5 #(
    .INIT(32'h00000004)
  ) __4742__ (
    .I4(__96__),
    .I3(__1100__),
    .I2(__876__),
    .I1(__720__),
    .I0(__825__),
    .O(__1362__)
  );
  LUT3 #(
    .INIT(8'hd0)
  ) __4743__ (
    .I2(__1362__),
    .I1(__185__),
    .I0(g35),
    .O(__1363__)
  );
  LUT5 #(
    .INIT(32'h00000001)
  ) __4744__ (
    .I4(__96__),
    .I3(__1100__),
    .I2(__876__),
    .I1(__720__),
    .I0(__825__),
    .O(__1364__)
  );
  LUT6 #(
    .INIT(64'h000d000000000000)
  ) __4745__ (
    .I5(__1364__),
    .I4(__1107__),
    .I3(__50__),
    .I2(__118__),
    .I1(__33__),
    .I0(g35),
    .O(__1365__)
  );
  LUT3 #(
    .INIT(8'hd0)
  ) __4746__ (
    .I2(__1357__),
    .I1(__459__),
    .I0(g35),
    .O(__1366__)
  );
  LUT3 #(
    .INIT(8'h01)
  ) __4747__ (
    .I2(__50__),
    .I1(__1107__),
    .I0(__118__),
    .O(__1367__)
  );
  LUT6 #(
    .INIT(64'h07007777ffffffff)
  ) __4748__ (
    .I5(__1367__),
    .I4(__1355__),
    .I3(g35),
    .I2(__497__),
    .I1(__1364__),
    .I0(__113__),
    .O(__1368__)
  );
  LUT3 #(
    .INIT(8'h04)
  ) __4749__ (
    .I2(__50__),
    .I1(__1107__),
    .I0(__118__),
    .O(__1369__)
  );
  LUT5 #(
    .INIT(32'h00000004)
  ) __4750__ (
    .I4(g56),
    .I3(g57),
    .I2(g53),
    .I1(g54),
    .I0(__968__),
    .O(__1370__)
  );
  LUT5 #(
    .INIT(32'hf0ba0000)
  ) __4751__ (
    .I4(__1370__),
    .I3(__96__),
    .I2(__1367__),
    .I1(__720__),
    .I0(__1369__),
    .O(__1371__)
  );
  LUT5 #(
    .INIT(32'hfeff0000)
  ) __4752__ (
    .I4(__1371__),
    .I3(__1368__),
    .I2(__1366__),
    .I1(__1365__),
    .I0(__1363__),
    .O(__1372__)
  );
  LUT5 #(
    .INIT(32'h00000080)
  ) __4753__ (
    .I4(__50__),
    .I3(__118__),
    .I2(__1107__),
    .I1(__1370__),
    .I0(__1357__),
    .O(__1373__)
  );
  LUT5 #(
    .INIT(32'h00000080)
  ) __4754__ (
    .I4(__50__),
    .I3(__1107__),
    .I2(__1364__),
    .I1(__118__),
    .I0(__1370__),
    .O(__1374__)
  );
  LUT6 #(
    .INIT(64'h0000000080000000)
  ) __4755__ (
    .I5(__118__),
    .I4(__1186__),
    .I3(__50__),
    .I2(__1107__),
    .I1(__1370__),
    .I0(__1362__),
    .O(__1375__)
  );
  LUT6 #(
    .INIT(64'h0000000080000000)
  ) __4756__ (
    .I5(__118__),
    .I4(__50__),
    .I3(__1107__),
    .I2(__1370__),
    .I1(__1357__),
    .I0(__938__),
    .O(__1376__)
  );
  LUT6 #(
    .INIT(64'h0000000000000777)
  ) __4757__ (
    .I5(__1376__),
    .I4(__1375__),
    .I3(__216__),
    .I2(__1374__),
    .I1(__1373__),
    .I0(__1182__),
    .O(__1377__)
  );
  LUT5 #(
    .INIT(32'h33333233)
  ) __4758__ (
    .I4(g56),
    .I3(g54),
    .I2(g57),
    .I1(g53),
    .I0(__968__),
    .O(__1378__)
  );
  LUT5 #(
    .INIT(32'h00000080)
  ) __4759__ (
    .I4(__1107__),
    .I3(__118__),
    .I2(__1364__),
    .I1(__50__),
    .I0(__1370__),
    .O(__1379__)
  );
  LUT5 #(
    .INIT(32'h00008000)
  ) __4760__ (
    .I4(__118__),
    .I3(__1364__),
    .I2(__50__),
    .I1(__1107__),
    .I0(__1370__),
    .O(__1380__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __4761__ (
    .I5(__65__),
    .I4(__1380__),
    .I3(__54__),
    .I2(__1379__),
    .I1(__248__),
    .I0(__1378__),
    .O(__1381__)
  );
  LUT6 #(
    .INIT(64'hdfffffffcfffffff)
  ) __4762__ (
    .I5(__1370__),
    .I4(__680__),
    .I3(__1381__),
    .I2(__1377__),
    .I1(__1372__),
    .I0(__1361__),
    .O(__1382__)
  );
  LUT6 #(
    .INIT(64'hfff4000000000000)
  ) __4763__ (
    .I5(__795__),
    .I4(__718__),
    .I3(__465__),
    .I2(__842__),
    .I1(__1285__),
    .I0(__101__),
    .O(__1383__)
  );
  LUT6 #(
    .INIT(64'h5adaaa2affff0000)
  ) __4764__ (
    .I5(g35),
    .I4(__1178__),
    .I3(__964__),
    .I2(__1383__),
    .I1(__1114__),
    .I0(__1016__),
    .O(__1384__)
  );
  LUT5 #(
    .INIT(32'h00009009)
  ) __4765__ (
    .I4(__605__),
    .I3(g72),
    .I2(__629__),
    .I1(g73),
    .I0(__664__),
    .O(__1385__)
  );
  LUT6 #(
    .INIT(64'h0000000000000008)
  ) __4766__ (
    .I5(g113),
    .I4(__1283__),
    .I3(__757__),
    .I2(__810__),
    .I1(__1385__),
    .I0(__236__),
    .O(__1386__)
  );
  LUT5 #(
    .INIT(32'h10ff0000)
  ) __4767__ (
    .I4(__1173__),
    .I3(g35),
    .I2(__418__),
    .I1(__989__),
    .I0(__1386__),
    .O(__1387__)
  );
  LUT4 #(
    .INIT(16'h7cfc)
  ) __4768__ (
    .I3(__1227__),
    .I2(__917__),
    .I1(__353__),
    .I0(__972__),
    .O(__1388__)
  );
  LUT4 #(
    .INIT(16'hef00)
  ) __4769__ (
    .I3(g35),
    .I2(__972__),
    .I1(__917__),
    .I0(__353__),
    .O(__1389__)
  );
  LUT6 #(
    .INIT(64'hffff44f400f000f0)
  ) __4770__ (
    .I5(__1389__),
    .I4(__348__),
    .I3(g35),
    .I2(__930__),
    .I1(__1388__),
    .I0(__866__),
    .O(__1390__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __4771__ (
    .I1(__1248__),
    .I0(__1245__),
    .O(__1391__)
  );
  LUT6 #(
    .INIT(64'h2aaad55500000000)
  ) __4772__ (
    .I5(g35),
    .I4(__1391__),
    .I3(__509__),
    .I2(__306__),
    .I1(__705__),
    .I0(__1073__),
    .O(__1392__)
  );
  LUT3 #(
    .INIT(8'h01)
  ) __4773__ (
    .I2(__1145__),
    .I1(__798__),
    .I0(__386__),
    .O(__1393__)
  );
  LUT2 #(
    .INIT(4'h2)
  ) __4774__ (
    .I1(__1034__),
    .I0(__962__),
    .O(__1394__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __4775__ (
    .I5(g35),
    .I4(__1394__),
    .I3(__1393__),
    .I2(__574__),
    .I1(__1054__),
    .I0(__1391__),
    .O(__1395__)
  );
  LUT5 #(
    .INIT(32'h00009009)
  ) __4776__ (
    .I4(__1240__),
    .I3(g72),
    .I2(__976__),
    .I1(g73),
    .I0(__738__),
    .O(__1396__)
  );
  LUT3 #(
    .INIT(8'hd0)
  ) __4777__ (
    .I2(__862__),
    .I1(__1168__),
    .I0(__1396__),
    .O(__1397__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __4778__ (
    .I1(__631__),
    .I0(__299__),
    .O(__1398__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __4779__ (
    .I1(__35__),
    .I0(__437__),
    .O(__1399__)
  );
  LUT3 #(
    .INIT(8'h08)
  ) __4780__ (
    .I2(__717__),
    .I1(__204__),
    .I0(__299__),
    .O(__1400__)
  );
  LUT6 #(
    .INIT(64'h4000ffff00000000)
  ) __4781__ (
    .I5(__1400__),
    .I4(__1399__),
    .I3(__289__),
    .I2(__555__),
    .I1(__713__),
    .I0(__1398__),
    .O(__1401__)
  );
  LUT6 #(
    .INIT(64'h3fc0bfc8f0f0f0f0)
  ) __4782__ (
    .I5(g35),
    .I4(__1115__),
    .I3(__881__),
    .I2(__660__),
    .I1(__170__),
    .I0(__1401__),
    .O(__1402__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __4783__ (
    .I1(__1111__),
    .I0(__908__),
    .O(__1403__)
  );
  LUT6 #(
    .INIT(64'h0000000082000082)
  ) __4784__ (
    .I5(__639__),
    .I4(__1030__),
    .I3(g72),
    .I2(g73),
    .I1(__456__),
    .I0(__845__),
    .O(__1404__)
  );
  LUT6 #(
    .INIT(64'h0000000041000041)
  ) __4785__ (
    .I5(__845__),
    .I4(__1030__),
    .I3(g72),
    .I2(g73),
    .I1(__456__),
    .I0(__639__),
    .O(__1405__)
  );
  LUT6 #(
    .INIT(64'h77770777ffffffff)
  ) __4786__ (
    .I5(__779__),
    .I4(__179__),
    .I3(__1405__),
    .I2(__728__),
    .I1(__1404__),
    .I0(__1403__),
    .O(__1406__)
  );
  LUT2 #(
    .INIT(4'h2)
  ) __4787__ (
    .I1(__1027__),
    .I0(__944__),
    .O(__1407__)
  );
  LUT6 #(
    .INIT(64'hffffffff2a3f3f3f)
  ) __4788__ (
    .I5(__779__),
    .I4(__1405__),
    .I3(__645__),
    .I2(__1404__),
    .I1(__1407__),
    .I0(__1014__),
    .O(__1408__)
  );
  LUT6 #(
    .INIT(64'h0000000082000082)
  ) __4789__ (
    .I5(__845__),
    .I4(__1030__),
    .I3(g72),
    .I2(g73),
    .I1(__456__),
    .I0(__639__),
    .O(__1409__)
  );
  LUT6 #(
    .INIT(64'hcfffcfffffff55ff)
  ) __4790__ (
    .I5(__779__),
    .I4(__617__),
    .I3(__1409__),
    .I2(__595__),
    .I1(__540__),
    .I0(__318__),
    .O(__1410__)
  );
  LUT6 #(
    .INIT(64'h8000080020000200)
  ) __4791__ (
    .I5(__1030__),
    .I4(g73),
    .I3(__845__),
    .I2(__456__),
    .I1(g72),
    .I0(__639__),
    .O(__1411__)
  );
  LUT6 #(
    .INIT(64'hcfffcfffffff55ff)
  ) __4792__ (
    .I5(__779__),
    .I4(__352__),
    .I3(__1411__),
    .I2(__196__),
    .I1(__190__),
    .I0(__746__),
    .O(__1412__)
  );
  LUT4 #(
    .INIT(16'hf800)
  ) __4793__ (
    .I3(g113),
    .I2(g134),
    .I1(__884__),
    .I0(g99),
    .O(__1413__)
  );
  LUT4 #(
    .INIT(16'h9009)
  ) __4794__ (
    .I3(__1030__),
    .I2(g72),
    .I1(g73),
    .I0(__456__),
    .O(__1414__)
  );
  LUT6 #(
    .INIT(64'h7fffffffffffffff)
  ) __4795__ (
    .I5(__1414__),
    .I4(__1413__),
    .I3(__1412__),
    .I2(__1410__),
    .I1(__1408__),
    .I0(__1406__),
    .O(__1415__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __4796__ (
    .I1(__900__),
    .I0(__817__),
    .O(__1416__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __4797__ (
    .I1(__566__),
    .I0(__548__),
    .O(__1417__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __4798__ (
    .I5(g35),
    .I4(__1417__),
    .I3(__1416__),
    .I2(__782__),
    .I1(__1086__),
    .I0(__1391__),
    .O(__1418__)
  );
  LUT3 #(
    .INIT(8'h78)
  ) __4799__ (
    .I2(__878__),
    .I1(g35),
    .I0(__206__),
    .O(__1419__)
  );
  LUT6 #(
    .INIT(64'h000000000000001f)
  ) __4800__ (
    .I5(__300__),
    .I4(__1008__),
    .I3(__918__),
    .I2(g35),
    .I1(__1099__),
    .I0(__1255__),
    .O(__1420__)
  );
  LUT3 #(
    .INIT(8'he0)
  ) __4801__ (
    .I2(g35),
    .I1(__1099__),
    .I0(__1255__),
    .O(__1421__)
  );
  LUT4 #(
    .INIT(16'h01ff)
  ) __4802__ (
    .I3(g35),
    .I2(__20__),
    .I1(__750__),
    .I0(__1265__),
    .O(__1422__)
  );
  LUT6 #(
    .INIT(64'h00000001ffffffff)
  ) __4803__ (
    .I5(g35),
    .I4(__300__),
    .I3(__1081__),
    .I2(__1008__),
    .I1(__298__),
    .I0(__918__),
    .O(__1423__)
  );
  LUT5 #(
    .INIT(32'hcfff4f5f)
  ) __4804__ (
    .I4(__1081__),
    .I3(__1423__),
    .I2(__1422__),
    .I1(__1421__),
    .I0(__1420__),
    .O(__1424__)
  );
  LUT6 #(
    .INIT(64'h0001001403033c3c)
  ) __4805__ (
    .I5(g35),
    .I4(__300__),
    .I3(__1099__),
    .I2(__1008__),
    .I1(__918__),
    .I0(__1255__),
    .O(__1425__)
  );
  LUT5 #(
    .INIT(32'h0000ca00)
  ) __4806__ (
    .I4(__298__),
    .I3(__1422__),
    .I2(__1081__),
    .I1(__1420__),
    .I0(__1425__),
    .O(__1426__)
  );
  LUT5 #(
    .INIT(32'h01160000)
  ) __4807__ (
    .I4(__1423__),
    .I3(__20__),
    .I2(__750__),
    .I1(__1265__),
    .I0(__1421__),
    .O(__1427__)
  );
  LUT3 #(
    .INIT(8'hfd)
  ) __4808__ (
    .I2(__1427__),
    .I1(__1426__),
    .I0(__1424__),
    .O(__1428__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __4809__ (
    .I1(__23__),
    .I0(__243__),
    .O(__1429__)
  );
  LUT6 #(
    .INIT(64'h00000000fff40000)
  ) __4810__ (
    .I5(__718__),
    .I4(__795__),
    .I3(__465__),
    .I2(__842__),
    .I1(__1285__),
    .I0(__821__),
    .O(__1430__)
  );
  LUT6 #(
    .INIT(64'h3caaaaaaf0f0f0f0)
  ) __4811__ (
    .I5(g35),
    .I4(__1430__),
    .I3(__1429__),
    .I2(__373__),
    .I1(__829__),
    .I0(__1094__),
    .O(__1431__)
  );
  LUT6 #(
    .INIT(64'h1115111511151111)
  ) __4812__ (
    .I5(g113),
    .I4(__1283__),
    .I3(g72),
    .I2(g73),
    .I1(__473__),
    .I0(__10__),
    .O(__1432__)
  );
  LUT6 #(
    .INIT(64'h7fd55555aa000000)
  ) __4813__ (
    .I5(__1268__),
    .I4(__1432__),
    .I3(__582__),
    .I2(__482__),
    .I1(__794__),
    .I0(g35),
    .O(__1433__)
  );
  LUT4 #(
    .INIT(16'hbbf0)
  ) __4814__ (
    .I3(g35),
    .I2(__399__),
    .I1(g44),
    .I0(__1057__),
    .O(__1434__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __4815__ (
    .I2(g35),
    .I1(g6750),
    .I0(__140__),
    .O(__1435__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __4816__ (
    .I1(__1236__),
    .I0(__1052__),
    .O(__1436__)
  );
  LUT6 #(
    .INIT(64'h8000080020000200)
  ) __4817__ (
    .I5(g72),
    .I4(g73),
    .I3(__1240__),
    .I2(__738__),
    .I1(__976__),
    .I0(__1436__),
    .O(__1437__)
  );
  LUT6 #(
    .INIT(64'hbfffffff00000000)
  ) __4818__ (
    .I5(__678__),
    .I4(__1310__),
    .I3(__69__),
    .I2(__727__),
    .I1(__1309__),
    .I0(__1077__),
    .O(__1438__)
  );
  LUT6 #(
    .INIT(64'h0077ff00f0f0f0f0)
  ) __4819__ (
    .I5(g35),
    .I4(__1438__),
    .I3(__1180__),
    .I2(__514__),
    .I1(__1338__),
    .I0(__1437__),
    .O(__1439__)
  );
  LUT5 #(
    .INIT(32'h82000082)
  ) __4820__ (
    .I4(g72),
    .I3(__976__),
    .I2(g73),
    .I1(__738__),
    .I0(__1240__),
    .O(__1440__)
  );
  LUT6 #(
    .INIT(64'h00000000aa800000)
  ) __4821__ (
    .I5(g113),
    .I4(__1440__),
    .I3(g134),
    .I2(__884__),
    .I1(g99),
    .I0(__15__),
    .O(__1441__)
  );
  LUT4 #(
    .INIT(16'h3740)
  ) __4822__ (
    .I3(__151__),
    .I2(__1192__),
    .I1(g35),
    .I0(__1441__),
    .O(__1442__)
  );
  LUT4 #(
    .INIT(16'h9009)
  ) __4823__ (
    .I3(g72),
    .I2(__591__),
    .I1(g73),
    .I0(__851__),
    .O(__1443__)
  );
  LUT5 #(
    .INIT(32'h0000f800)
  ) __4824__ (
    .I4(g113),
    .I3(__749__),
    .I2(g134),
    .I1(__884__),
    .I0(g99),
    .O(__1444__)
  );
  LUT5 #(
    .INIT(32'h00008000)
  ) __4825__ (
    .I4(__917__),
    .I3(__353__),
    .I2(__972__),
    .I1(__1444__),
    .I0(__1443__),
    .O(__1445__)
  );
  LUT6 #(
    .INIT(64'h00000000fff40000)
  ) __4826__ (
    .I5(__795__),
    .I4(__718__),
    .I3(__465__),
    .I2(__842__),
    .I1(__1285__),
    .I0(__503__),
    .O(__1446__)
  );
  LUT5 #(
    .INIT(32'hffa0cfc0)
  ) __4827__ (
    .I4(__1446__),
    .I3(__462__),
    .I2(g35),
    .I1(__469__),
    .I0(__1445__),
    .O(__1447__)
  );
  LUT6 #(
    .INIT(64'h00dfdf00ffff0000)
  ) __4828__ (
    .I5(g35),
    .I4(__688__),
    .I3(__636__),
    .I2(__1303__),
    .I1(__810__),
    .I0(__1294__),
    .O(__1448__)
  );
  LUT6 #(
    .INIT(64'h1001000000000000)
  ) __4829__ (
    .I5(__560__),
    .I4(__1124__),
    .I3(__1228__),
    .I2(__579__),
    .I1(__939__),
    .I0(__1013__),
    .O(__1449__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __4830__ (
    .I2(__1449__),
    .I1(__584__),
    .I0(__77__),
    .O(__1450__)
  );
  LUT4 #(
    .INIT(16'h8000)
  ) __4831__ (
    .I3(__1043__),
    .I2(__1110__),
    .I1(__762__),
    .I0(__1251__),
    .O(__1451__)
  );
  LUT6 #(
    .INIT(64'h0000000000008000)
  ) __4832__ (
    .I5(__779__),
    .I4(__845__),
    .I3(__1030__),
    .I2(__456__),
    .I1(__1451__),
    .I0(__53__),
    .O(__1452__)
  );
  LUT6 #(
    .INIT(64'h1a001a00ffff0000)
  ) __4833__ (
    .I5(g35),
    .I4(__599__),
    .I3(__758__),
    .I2(__1452__),
    .I1(__1450__),
    .I0(__397__),
    .O(__1453__)
  );
  LUT6 #(
    .INIT(64'h880a000000000000)
  ) __4834__ (
    .I5(__185__),
    .I4(__218__),
    .I3(__751__),
    .I2(__350__),
    .I1(__869__),
    .I0(__886__),
    .O(__1454__)
  );
  LUT6 #(
    .INIT(64'h8000000000000000)
  ) __4835__ (
    .I5(__764__),
    .I4(__880__),
    .I3(__207__),
    .I2(__854__),
    .I1(__1113__),
    .I0(__1454__),
    .O(__1455__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __4836__ (
    .I2(__981__),
    .I1(__33__),
    .I0(__1455__),
    .O(__1456__)
  );
  LUT6 #(
    .INIT(64'h6c206c6cf0f0f0f0)
  ) __4837__ (
    .I5(g35),
    .I4(__751__),
    .I3(__869__),
    .I2(__744__),
    .I1(__199__),
    .I0(__1456__),
    .O(__1457__)
  );
  LUT6 #(
    .INIT(64'h06666666aaaaaaaa)
  ) __4838__ (
    .I5(g35),
    .I4(__1303__),
    .I3(__810__),
    .I2(__1294__),
    .I1(__509__),
    .I0(__306__),
    .O(__1458__)
  );
  LUT6 #(
    .INIT(64'h0000000082000082)
  ) __4839__ (
    .I5(__917__),
    .I4(g72),
    .I3(__591__),
    .I2(g73),
    .I1(__851__),
    .I0(__353__),
    .O(__1459__)
  );
  LUT6 #(
    .INIT(64'h3f3f002affff00aa)
  ) __4840__ (
    .I5(__972__),
    .I4(__784__),
    .I3(__462__),
    .I2(__1444__),
    .I1(__1459__),
    .I0(__469__),
    .O(__1460__)
  );
  LUT5 #(
    .INIT(32'h33aaf0f0)
  ) __4841__ (
    .I4(g35),
    .I3(__1446__),
    .I2(__1116__),
    .I1(__1460__),
    .I0(__462__),
    .O(__1461__)
  );
  LUT4 #(
    .INIT(16'h8000)
  ) __4842__ (
    .I3(__795__),
    .I2(__718__),
    .I1(__465__),
    .I0(__842__),
    .O(__1462__)
  );
  LUT4 #(
    .INIT(16'h8000)
  ) __4843__ (
    .I3(__1227__),
    .I2(__917__),
    .I1(__972__),
    .I0(__1462__),
    .O(__1463__)
  );
  LUT5 #(
    .INIT(32'h78ccffcc)
  ) __4844__ (
    .I4(__650__),
    .I3(g35),
    .I2(__591__),
    .I1(__353__),
    .I0(__1463__),
    .O(__1464__)
  );
  LUT6 #(
    .INIT(64'h0000000082000082)
  ) __4845__ (
    .I5(__353__),
    .I4(g72),
    .I3(__591__),
    .I2(g73),
    .I1(__851__),
    .I0(__917__),
    .O(__1465__)
  );
  LUT5 #(
    .INIT(32'h00000008)
  ) __4846__ (
    .I4(__972__),
    .I3(g113),
    .I2(__1283__),
    .I1(__749__),
    .I0(__1465__),
    .O(__1466__)
  );
  LUT6 #(
    .INIT(64'heeeef0f0ff00ff00)
  ) __4847__ (
    .I5(g35),
    .I4(__1430__),
    .I3(__957__),
    .I2(__142__),
    .I1(__23__),
    .I0(__1466__),
    .O(__1467__)
  );
  LUT3 #(
    .INIT(8'hfd)
  ) __4848__ (
    .I2(__99__),
    .I1(__1018__),
    .I0(g35),
    .O(__1468__)
  );
  LUT6 #(
    .INIT(64'h0000fff300005551)
  ) __4849__ (
    .I5(__1118__),
    .I4(__1342__),
    .I3(__493__),
    .I2(__65__),
    .I1(__895__),
    .I0(__500__),
    .O(__1469__)
  );
  LUT6 #(
    .INIT(64'h0a0a5f0a0a0a1b0a)
  ) __4850__ (
    .I5(__1118__),
    .I4(__1342__),
    .I3(__1248__),
    .I2(__739__),
    .I1(__500__),
    .I0(__1469__),
    .O(__1470__)
  );
  LUT4 #(
    .INIT(16'hbf00)
  ) __4851__ (
    .I3(__484__),
    .I2(__1345__),
    .I1(__660__),
    .I0(__881__),
    .O(__1471__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __4852__ (
    .I1(__500__),
    .I0(__1118__),
    .O(__1472__)
  );
  LUT6 #(
    .INIT(64'h00000000000000fd)
  ) __4853__ (
    .I5(__1342__),
    .I4(__1472__),
    .I3(__1471__),
    .I2(__493__),
    .I1(__65__),
    .I0(__895__),
    .O(__1473__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __4854__ (
    .I1(__645__),
    .I0(__1473__),
    .O(__1474__)
  );
  LUT6 #(
    .INIT(64'hf055f0f0cccccccc)
  ) __4855__ (
    .I5(g35),
    .I4(__1474__),
    .I3(__1014__),
    .I2(__828__),
    .I1(__63__),
    .I0(__1470__),
    .O(__1475__)
  );
  LUT6 #(
    .INIT(64'hffffff00efefefef)
  ) __4856__ (
    .I5(__1249__),
    .I4(__639__),
    .I3(__53__),
    .I2(__237__),
    .I1(__996__),
    .I0(__1183__),
    .O(__1476__)
  );
  LUT5 #(
    .INIT(32'h00000080)
  ) __4857__ (
    .I4(__1043__),
    .I3(__1476__),
    .I2(__1110__),
    .I1(__762__),
    .I0(__1251__),
    .O(__1477__)
  );
  LUT5 #(
    .INIT(32'hccaaf0f0)
  ) __4858__ (
    .I4(g35),
    .I3(__1477__),
    .I2(__1124__),
    .I1(__560__),
    .I0(__1013__),
    .O(__1478__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __4859__ (
    .I1(__1202__),
    .I0(__1157__),
    .O(__1479__)
  );
  LUT6 #(
    .INIT(64'h0000000000000004)
  ) __4860__ (
    .I5(__554__),
    .I4(__169__),
    .I3(__257__),
    .I2(__49__),
    .I1(__1479__),
    .I0(__521__),
    .O(__1480__)
  );
  LUT3 #(
    .INIT(8'h35)
  ) __4861__ (
    .I2(__1204__),
    .I1(__406__),
    .I0(__1108__),
    .O(__1481__)
  );
  LUT5 #(
    .INIT(32'hf0343cf8)
  ) __4862__ (
    .I4(__1481__),
    .I3(__815__),
    .I2(__600__),
    .I1(g35),
    .I0(__1480__),
    .O(__1482__)
  );
  LUT5 #(
    .INIT(32'h82000082)
  ) __4863__ (
    .I4(__1030__),
    .I3(g72),
    .I2(g73),
    .I1(__456__),
    .I0(__845__),
    .O(__1483__)
  );
  LUT6 #(
    .INIT(64'h0000000000008000)
  ) __4864__ (
    .I5(g113),
    .I4(__1283__),
    .I3(__1060__),
    .I2(__779__),
    .I1(__639__),
    .I0(__1483__),
    .O(__1484__)
  );
  LUT6 #(
    .INIT(64'h00000000cfdfffff)
  ) __4865__ (
    .I5(g134),
    .I4(__1249__),
    .I3(__1207__),
    .I2(__1041__),
    .I1(__304__),
    .I0(__936__),
    .O(__1485__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __4866__ (
    .I1(__245__),
    .I0(__441__),
    .O(__1486__)
  );
  LUT6 #(
    .INIT(64'h0000000000000008)
  ) __4867__ (
    .I5(__1181__),
    .I4(__770__),
    .I3(__1072__),
    .I2(__1233__),
    .I1(__544__),
    .I0(__269__),
    .O(__1487__)
  );
  LUT4 #(
    .INIT(16'h7f00)
  ) __4868__ (
    .I3(__998__),
    .I2(__1487__),
    .I1(__507__),
    .I0(__1032__),
    .O(__1488__)
  );
  LUT6 #(
    .INIT(64'h00000000000000f7)
  ) __4869__ (
    .I5(__1488__),
    .I4(__1486__),
    .I3(__1485__),
    .I2(__1186__),
    .I1(__1143__),
    .I0(__961__),
    .O(__1489__)
  );
  LUT5 #(
    .INIT(32'haaf030f0)
  ) __4870__ (
    .I4(__1489__),
    .I3(g35),
    .I2(__190__),
    .I1(__1484__),
    .I0(__196__),
    .O(__1490__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __4871__ (
    .I1(__1276__),
    .I0(__30__),
    .O(__1491__)
  );
  LUT6 #(
    .INIT(64'h007f00ffffff0000)
  ) __4872__ (
    .I5(g35),
    .I4(__395__),
    .I3(__514__),
    .I2(__56__),
    .I1(__635__),
    .I0(__1491__),
    .O(__1492__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __4873__ (
    .I2(__457__),
    .I1(__874__),
    .I0(__1264__),
    .O(__1493__)
  );
  LUT6 #(
    .INIT(64'hee22eeeef0f0f0f0)
  ) __4874__ (
    .I5(g35),
    .I4(__1248__),
    .I3(__1245__),
    .I2(__1056__),
    .I1(__1493__),
    .I0(__1219__),
    .O(__1494__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __4875__ (
    .I1(g35),
    .I0(__253__),
    .O(__1495__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __4876__ (
    .I2(g35),
    .I1(__773__),
    .I0(__505__),
    .O(__1496__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __4877__ (
    .I1(__152__),
    .I0(__365__),
    .O(__1497__)
  );
  LUT5 #(
    .INIT(32'habff5400)
  ) __4878__ (
    .I4(__1022__),
    .I3(__1115__),
    .I2(__35__),
    .I1(__437__),
    .I0(__667__),
    .O(__1498__)
  );
  LUT3 #(
    .INIT(8'h04)
  ) __4879__ (
    .I2(__881__),
    .I1(__580__),
    .I0(__660__),
    .O(__1499__)
  );
  LUT6 #(
    .INIT(64'hfa00f0f0cccccccc)
  ) __4880__ (
    .I5(g35),
    .I4(__1499__),
    .I3(__1498__),
    .I2(__1146__),
    .I1(__943__),
    .I0(__1497__),
    .O(__1500__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __4881__ (
    .I1(g35),
    .I0(__573__),
    .O(__1501__)
  );
  LUT6 #(
    .INIT(64'h000c000500000000)
  ) __4882__ (
    .I5(__1501__),
    .I4(__30__),
    .I3(__217__),
    .I2(__56__),
    .I1(__1276__),
    .I0(__635__),
    .O(__1502__)
  );
  LUT4 #(
    .INIT(16'h00f8)
  ) __4883__ (
    .I3(g113),
    .I2(g134),
    .I1(__884__),
    .I0(g99),
    .O(__1503__)
  );
  LUT6 #(
    .INIT(64'h8000000000000000)
  ) __4884__ (
    .I5(__465__),
    .I4(__842__),
    .I3(__1227__),
    .I2(__917__),
    .I1(__353__),
    .I0(__972__),
    .O(__1504__)
  );
  LUT6 #(
    .INIT(64'h0c3fff00aaaaff00)
  ) __4885__ (
    .I5(__1504__),
    .I4(g35),
    .I3(__993__),
    .I2(__1098__),
    .I1(__1503__),
    .I0(__38__),
    .O(__1505__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __4886__ (
    .I2(__962__),
    .I1(__1145__),
    .I0(__1034__),
    .O(__1506__)
  );
  LUT6 #(
    .INIT(64'hee22eeeef0f0f0f0)
  ) __4887__ (
    .I5(g35),
    .I4(__1248__),
    .I3(__1245__),
    .I2(__797__),
    .I1(__1506__),
    .I0(__1212__),
    .O(__1507__)
  );
  LUT6 #(
    .INIT(64'h0000000000000001)
  ) __4888__ (
    .I5(__757__),
    .I4(__605__),
    .I3(__810__),
    .I2(__445__),
    .I1(__519__),
    .I0(__1224__),
    .O(__1508__)
  );
  LUT6 #(
    .INIT(64'hccccccacaaaaaaaa)
  ) __4889__ (
    .I5(g35),
    .I4(__1190__),
    .I3(__614__),
    .I2(__1508__),
    .I1(__1025__),
    .I0(__1108__),
    .O(__1509__)
  );
  LUT4 #(
    .INIT(16'hca00)
  ) __4890__ (
    .I3(g35),
    .I2(__1451__),
    .I1(__1046__),
    .I0(__237__),
    .O(__1510__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __4891__ (
    .I2(g35),
    .I1(__367__),
    .I0(__1072__),
    .O(__1511__)
  );
  LUT6 #(
    .INIT(64'h00000000a8a8a8aa)
  ) __4892__ (
    .I5(__180__),
    .I4(__1283__),
    .I3(__1257__),
    .I2(g72),
    .I1(g73),
    .I0(__329__),
    .O(__1512__)
  );
  LUT6 #(
    .INIT(64'hffffbf00ff00ff00)
  ) __4893__ (
    .I5(g35),
    .I4(__1512__),
    .I3(__913__),
    .I2(__10__),
    .I1(__84__),
    .I0(__486__),
    .O(__1513__)
  );
  LUT4 #(
    .INIT(16'h0777)
  ) __4894__ (
    .I3(__671__),
    .I2(__177__),
    .I1(__695__),
    .I0(__414__),
    .O(__1514__)
  );
  LUT6 #(
    .INIT(64'hccfff0f0a000f0f0)
  ) __4895__ (
    .I5(__875__),
    .I4(g35),
    .I3(__1451__),
    .I2(__758__),
    .I1(__1514__),
    .I0(__671__),
    .O(__1515__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __4896__ (
    .I1(__151__),
    .I0(__1192__),
    .O(__1516__)
  );
  LUT5 #(
    .INIT(32'h00007fff)
  ) __4897__ (
    .I4(__1441__),
    .I3(__151__),
    .I2(__926__),
    .I1(__995__),
    .I0(__1192__),
    .O(__1517__)
  );
  LUT6 #(
    .INIT(64'hf8fff00000ff0000)
  ) __4898__ (
    .I5(__1517__),
    .I4(__241__),
    .I3(g35),
    .I2(__995__),
    .I1(__926__),
    .I0(__1516__),
    .O(__1518__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __4899__ (
    .I1(__943__),
    .I0(__1118__),
    .O(__1519__)
  );
  LUT4 #(
    .INIT(16'h7f00)
  ) __4900__ (
    .I3(__1009__),
    .I2(__1345__),
    .I1(__881__),
    .I0(__660__),
    .O(__1520__)
  );
  LUT6 #(
    .INIT(64'h00000000000000f7)
  ) __4901__ (
    .I5(__1342__),
    .I4(__1520__),
    .I3(__1519__),
    .I2(__65__),
    .I1(__493__),
    .I0(__895__),
    .O(__1521__)
  );
  LUT5 #(
    .INIT(32'h00009009)
  ) __4902__ (
    .I4(__845__),
    .I3(__1030__),
    .I2(g72),
    .I1(g73),
    .I0(__456__),
    .O(__1522__)
  );
  LUT6 #(
    .INIT(64'h0000000000008000)
  ) __4903__ (
    .I5(g113),
    .I4(__1283__),
    .I3(__1060__),
    .I2(__779__),
    .I1(__1522__),
    .I0(__639__),
    .O(__1523__)
  );
  LUT6 #(
    .INIT(64'hc0c0c0cd00000000)
  ) __4904__ (
    .I5(g35),
    .I4(__595__),
    .I3(__1523__),
    .I2(__1521__),
    .I1(__112__),
    .I0(__540__),
    .O(__1524__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __4905__ (
    .I2(__509__),
    .I1(__306__),
    .I0(__705__),
    .O(__1525__)
  );
  LUT6 #(
    .INIT(64'hee22eeeef0f0f0f0)
  ) __4906__ (
    .I5(g35),
    .I4(__1248__),
    .I3(__1245__),
    .I2(__714__),
    .I1(__1525__),
    .I0(__831__),
    .O(__1526__)
  );
  LUT6 #(
    .INIT(64'habffabffffff0000)
  ) __4907__ (
    .I5(g35),
    .I4(__432__),
    .I3(__1115__),
    .I2(__35__),
    .I1(__437__),
    .I0(__1182__),
    .O(__1527__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __4908__ (
    .I2(__157__),
    .I1(__561__),
    .I0(__863__),
    .O(__1528__)
  );
  LUT6 #(
    .INIT(64'hee22eeeef0f0f0f0)
  ) __4909__ (
    .I5(g35),
    .I4(__1248__),
    .I3(__1245__),
    .I2(__420__),
    .I1(__1528__),
    .I0(__899__),
    .O(__1529__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __4910__ (
    .I1(__786__),
    .I0(__693__),
    .O(__1530__)
  );
  LUT4 #(
    .INIT(16'h0080)
  ) __4911__ (
    .I3(__1043__),
    .I2(__1110__),
    .I1(__762__),
    .I0(__1251__),
    .O(__1531__)
  );
  LUT6 #(
    .INIT(64'h0000000000000004)
  ) __4912__ (
    .I5(__1030__),
    .I4(__456__),
    .I3(__845__),
    .I2(__639__),
    .I1(__1531__),
    .I0(__53__),
    .O(__1532__)
  );
  LUT6 #(
    .INIT(64'hff81ffff00000000)
  ) __4913__ (
    .I5(__1249__),
    .I4(__1532__),
    .I3(__1530__),
    .I2(__584__),
    .I1(__244__),
    .I0(__77__),
    .O(__1533__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __4914__ (
    .I1(__198__),
    .I0(__410__),
    .O(__1534__)
  );
  LUT6 #(
    .INIT(64'h0000000000004000)
  ) __4915__ (
    .I5(__501__),
    .I4(__439__),
    .I3(__22__),
    .I2(__149__),
    .I1(__1534__),
    .I0(__34__),
    .O(__1535__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __4916__ (
    .I1(__83__),
    .I0(__1535__),
    .O(__1536__)
  );
  LUT3 #(
    .INIT(8'h01)
  ) __4917__ (
    .I2(__198__),
    .I1(__410__),
    .I0(__22__),
    .O(__1537__)
  );
  LUT6 #(
    .INIT(64'h00000000bfffffff)
  ) __4918__ (
    .I5(__83__),
    .I4(__1537__),
    .I3(__501__),
    .I2(__439__),
    .I1(__34__),
    .I0(__149__),
    .O(__1538__)
  );
  LUT6 #(
    .INIT(64'h0000000000008000)
  ) __4919__ (
    .I5(__1538__),
    .I4(__1536__),
    .I3(__182__),
    .I2(__129__),
    .I1(__387__),
    .I0(__1533__),
    .O(__1539__)
  );
  LUT6 #(
    .INIT(64'h007e7e7e00000000)
  ) __4920__ (
    .I5(__1532__),
    .I4(__786__),
    .I3(__693__),
    .I2(__584__),
    .I1(__244__),
    .I0(__77__),
    .O(__1540__)
  );
  LUT5 #(
    .INIT(32'h000000d0)
  ) __4921__ (
    .I4(__1540__),
    .I3(__1538__),
    .I2(__1249__),
    .I1(__1535__),
    .I0(__83__),
    .O(__1541__)
  );
  LUT5 #(
    .INIT(32'h73bbc000)
  ) __4922__ (
    .I4(__210__),
    .I3(__333__),
    .I2(__1541__),
    .I1(g35),
    .I0(__1539__),
    .O(__1542__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __4923__ (
    .I2(g35),
    .I1(__1071__),
    .I0(__508__),
    .O(__1543__)
  );
  LUT6 #(
    .INIT(64'hdfff7555aaaa0000)
  ) __4924__ (
    .I5(__1146__),
    .I4(__1022__),
    .I3(__152__),
    .I2(__1499__),
    .I1(__985__),
    .I0(g35),
    .O(__1544__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __4925__ (
    .I1(__775__),
    .I0(__766__),
    .O(__1545__)
  );
  LUT6 #(
    .INIT(64'h331100001f3f0000)
  ) __4926__ (
    .I5(__544__),
    .I4(__1207__),
    .I3(__396__),
    .I2(__646__),
    .I1(__1545__),
    .I0(__594__),
    .O(__1546__)
  );
  LUT6 #(
    .INIT(64'hafaaeaaaff00ff00)
  ) __4927__ (
    .I5(g35),
    .I4(__544__),
    .I3(__936__),
    .I2(__396__),
    .I1(__646__),
    .I0(__1546__),
    .O(__1547__)
  );
  LUT5 #(
    .INIT(32'h80000000)
  ) __4928__ (
    .I4(__1043__),
    .I3(__1110__),
    .I2(__762__),
    .I1(__1251__),
    .I0(__265__),
    .O(__1548__)
  );
  LUT4 #(
    .INIT(16'h4f00)
  ) __4929__ (
    .I3(g35),
    .I2(__671__),
    .I1(__875__),
    .I0(__177__),
    .O(__1549__)
  );
  LUT5 #(
    .INIT(32'h7df05500)
  ) __4930__ (
    .I4(__1549__),
    .I3(__695__),
    .I2(__403__),
    .I1(__1548__),
    .I0(g35),
    .O(__1550__)
  );
  LUT6 #(
    .INIT(64'h00003fff00001555)
  ) __4931__ (
    .I5(__441__),
    .I4(__1485__),
    .I3(__1143__),
    .I2(__1186__),
    .I1(__961__),
    .I0(__1189__),
    .O(__1551__)
  );
  LUT6 #(
    .INIT(64'h88d8888888d888d8)
  ) __4932__ (
    .I5(__1189__),
    .I4(__441__),
    .I3(__1485__),
    .I2(__1248__),
    .I1(__768__),
    .I0(__1551__),
    .O(__1552__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __4933__ (
    .I1(__1189__),
    .I0(__441__),
    .O(__1553__)
  );
  LUT4 #(
    .INIT(16'hef00)
  ) __4934__ (
    .I3(__385__),
    .I2(__1487__),
    .I1(__507__),
    .I0(__1032__),
    .O(__1554__)
  );
  LUT6 #(
    .INIT(64'h000000000000007f)
  ) __4935__ (
    .I5(__1485__),
    .I4(__1554__),
    .I3(__1553__),
    .I2(__1143__),
    .I1(__1186__),
    .I0(__961__),
    .O(__1555__)
  );
  LUT3 #(
    .INIT(8'h01)
  ) __4936__ (
    .I2(__746__),
    .I1(__793__),
    .I0(__1555__),
    .O(__1556__)
  );
  LUT5 #(
    .INIT(32'h33aaf0f0)
  ) __4937__ (
    .I4(g35),
    .I3(__1556__),
    .I2(__332__),
    .I1(__1552__),
    .I0(__668__),
    .O(__1557__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __4938__ (
    .I1(__386__),
    .I0(__798__),
    .O(__1558__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __4939__ (
    .I5(g35),
    .I4(__1394__),
    .I3(__1558__),
    .I2(__1007__),
    .I1(__1163__),
    .I0(__1391__),
    .O(__1559__)
  );
  LUT6 #(
    .INIT(64'h0c3fff00aaaaff00)
  ) __4940__ (
    .I5(__1504__),
    .I4(g35),
    .I3(__81__),
    .I2(__999__),
    .I1(__1503__),
    .I0(__101__),
    .O(__1560__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __4941__ (
    .I1(__819__),
    .I0(__1109__),
    .O(__1561__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __4942__ (
    .I1(__70__),
    .I0(__819__),
    .O(__1562__)
  );
  LUT6 #(
    .INIT(64'hffccff00f0f0fafa)
  ) __4943__ (
    .I5(__769__),
    .I4(__982__),
    .I3(__1562__),
    .I2(__1561__),
    .I1(__987__),
    .I0(__923__),
    .O(__1563__)
  );
  LUT5 #(
    .INIT(32'h0f05030f)
  ) __4944__ (
    .I4(__819__),
    .I3(__982__),
    .I2(__1563__),
    .I1(__927__),
    .I0(__1021__),
    .O(__1564__)
  );
  LUT5 #(
    .INIT(32'h33aaf0f0)
  ) __4945__ (
    .I4(g35),
    .I3(__1286__),
    .I2(__982__),
    .I1(__1564__),
    .I0(__552__),
    .O(__1565__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __4946__ (
    .I1(__870__),
    .I0(__648__),
    .O(__1566__)
  );
  LUT4 #(
    .INIT(16'h9009)
  ) __4947__ (
    .I3(g72),
    .I2(__976__),
    .I1(g73),
    .I0(__738__),
    .O(__1567__)
  );
  LUT4 #(
    .INIT(16'h0004)
  ) __4948__ (
    .I3(__1240__),
    .I2(__1052__),
    .I1(__1567__),
    .I0(__1236__),
    .O(__1568__)
  );
  LUT4 #(
    .INIT(16'h0008)
  ) __4949__ (
    .I3(__1052__),
    .I2(__1236__),
    .I1(__1240__),
    .I0(__1567__),
    .O(__1569__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __4950__ (
    .I1(__527__),
    .I0(__254__),
    .O(__1570__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __4951__ (
    .I1(__1211__),
    .I0(__46__),
    .O(__1571__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __4952__ (
    .I1(__1154__),
    .I0(__1126__),
    .O(__1572__)
  );
  LUT6 #(
    .INIT(64'hf5f3ffffffffffff)
  ) __4953__ (
    .I5(__1567__),
    .I4(__1052__),
    .I3(__1240__),
    .I2(__1236__),
    .I1(__1572__),
    .I0(__1571__),
    .O(__1573__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __4954__ (
    .I1(__511__),
    .I0(__820__),
    .O(__1574__)
  );
  LUT6 #(
    .INIT(64'h77ff0fffffffffff)
  ) __4955__ (
    .I5(__1396__),
    .I4(__1052__),
    .I3(__1236__),
    .I2(__1574__),
    .I1(__726__),
    .I0(__830__),
    .O(__1575__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __4956__ (
    .I1(__1180__),
    .I0(__691__),
    .O(__1576__)
  );
  LUT6 #(
    .INIT(64'h002a2a2aaaaaaaaa)
  ) __4957__ (
    .I5(__1440__),
    .I4(__1576__),
    .I3(__1436__),
    .I2(__1336__),
    .I1(__1320__),
    .I0(__1575__),
    .O(__1577__)
  );
  LUT6 #(
    .INIT(64'hf888ffffffffffff)
  ) __4958__ (
    .I5(__1577__),
    .I4(__1573__),
    .I3(__1570__),
    .I2(__1569__),
    .I1(__1568__),
    .I0(__1566__),
    .O(__1578__)
  );
  LUT4 #(
    .INIT(16'h7fff)
  ) __4959__ (
    .I3(__1412__),
    .I2(__1410__),
    .I1(__1408__),
    .I0(__1406__),
    .O(__1579__)
  );
  LUT6 #(
    .INIT(64'h7f33b3b3cc000000)
  ) __4960__ (
    .I5(__333__),
    .I4(__381__),
    .I3(__1541__),
    .I2(__1539__),
    .I1(g35),
    .I0(__210__),
    .O(__1580__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __4961__ (
    .I1(__541__),
    .I0(__1197__),
    .O(__1581__)
  );
  LUT6 #(
    .INIT(64'hc3aaaaaaf0f0f0f0)
  ) __4962__ (
    .I5(g35),
    .I4(__1299__),
    .I3(__1581__),
    .I2(__893__),
    .I1(__850__),
    .I0(__231__),
    .O(__1582__)
  );
  LUT6 #(
    .INIT(64'heeeef0f0ff00ff00)
  ) __4963__ (
    .I5(g35),
    .I4(__1446__),
    .I3(__1201__),
    .I2(__784__),
    .I1(__469__),
    .I0(__1445__),
    .O(__1583__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __4964__ (
    .I2(__468__),
    .I1(__704__),
    .I0(__898__),
    .O(__1584__)
  );
  LUT5 #(
    .INIT(32'hc3aaf0f0)
  ) __4965__ (
    .I4(g35),
    .I3(__1584__),
    .I2(__490__),
    .I1(__271__),
    .I0(__571__),
    .O(__1585__)
  );
  LUT3 #(
    .INIT(8'h08)
  ) __4966__ (
    .I2(__1110__),
    .I1(__762__),
    .I0(__1251__),
    .O(__1586__)
  );
  LUT6 #(
    .INIT(64'hfff07f70ffff0000)
  ) __4967__ (
    .I5(g35),
    .I4(__1249__),
    .I3(__461__),
    .I2(__1586__),
    .I1(__758__),
    .I0(__1450__),
    .O(__1587__)
  );
  LUT6 #(
    .INIT(64'hccccacccaaaaaaaa)
  ) __4968__ (
    .I5(g35),
    .I4(__1110__),
    .I3(__762__),
    .I2(__1251__),
    .I1(__599__),
    .I0(__461__),
    .O(__1588__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __4969__ (
    .I1(__23__),
    .I0(__837__),
    .O(__1589__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __4970__ (
    .I1(__608__),
    .I0(__23__),
    .O(__1590__)
  );
  LUT6 #(
    .INIT(64'hffccff00f0f0fafa)
  ) __4971__ (
    .I5(__243__),
    .I4(__142__),
    .I3(__1590__),
    .I2(__1589__),
    .I1(__1051__),
    .I0(__8__),
    .O(__1591__)
  );
  LUT5 #(
    .INIT(32'h0f05030f)
  ) __4972__ (
    .I4(__142__),
    .I3(__23__),
    .I2(__1591__),
    .I1(__26__),
    .I0(__1277__),
    .O(__1592__)
  );
  LUT5 #(
    .INIT(32'h33aaf0f0)
  ) __4973__ (
    .I4(g35),
    .I3(__1430__),
    .I2(__142__),
    .I1(__1592__),
    .I0(__537__),
    .O(__1593__)
  );
  LUT4 #(
    .INIT(16'h8000)
  ) __4974__ (
    .I3(__379__),
    .I2(__759__),
    .I1(__474__),
    .I0(__724__),
    .O(__1594__)
  );
  LUT4 #(
    .INIT(16'h3caa)
  ) __4975__ (
    .I3(g35),
    .I2(__847__),
    .I1(__1594__),
    .I0(__885__),
    .O(__1595__)
  );
  LUT6 #(
    .INIT(64'h0000fff300005551)
  ) __4976__ (
    .I5(__441__),
    .I4(__1485__),
    .I3(__1143__),
    .I2(__1186__),
    .I1(__961__),
    .I0(__334__),
    .O(__1596__)
  );
  LUT6 #(
    .INIT(64'h0a0a5f0a0a0a1b0a)
  ) __4977__ (
    .I5(__441__),
    .I4(__1485__),
    .I3(__1248__),
    .I2(__768__),
    .I1(__334__),
    .I0(__1596__),
    .O(__1597__)
  );
  LUT4 #(
    .INIT(16'hbf00)
  ) __4978__ (
    .I3(__674__),
    .I2(__1487__),
    .I1(__1032__),
    .I0(__507__),
    .O(__1598__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __4979__ (
    .I1(__334__),
    .I0(__441__),
    .O(__1599__)
  );
  LUT6 #(
    .INIT(64'h00000000000000fd)
  ) __4980__ (
    .I5(__1485__),
    .I4(__1599__),
    .I3(__1598__),
    .I2(__1143__),
    .I1(__1186__),
    .I0(__961__),
    .O(__1600__)
  );
  LUT6 #(
    .INIT(64'hf055f0f0cccccccc)
  ) __4981__ (
    .I5(g35),
    .I4(__1289__),
    .I3(__1600__),
    .I2(__70__),
    .I1(__1021__),
    .I0(__1597__),
    .O(__1601__)
  );
  LUT3 #(
    .INIT(8'h04)
  ) __4982__ (
    .I2(__507__),
    .I1(__709__),
    .I0(__1032__),
    .O(__1602__)
  );
  LUT5 #(
    .INIT(32'h7f300000)
  ) __4983__ (
    .I4(g35),
    .I3(__489__),
    .I2(__1602__),
    .I1(__88__),
    .I0(__835__),
    .O(__1603__)
  );
  LUT5 #(
    .INIT(32'hccaaf0f0)
  ) __4984__ (
    .I4(g35),
    .I3(__364__),
    .I2(__507__),
    .I1(__396__),
    .I0(__1263__),
    .O(__1604__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __4985__ (
    .I1(__746__),
    .I0(__1555__),
    .O(__1605__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __4986__ (
    .I5(g35),
    .I4(__793__),
    .I3(__1605__),
    .I2(__669__),
    .I1(__402__),
    .I0(__1552__),
    .O(__1606__)
  );
  LUT5 #(
    .INIT(32'h7d55a000)
  ) __4987__ (
    .I4(__387__),
    .I3(__1541__),
    .I2(__129__),
    .I1(__182__),
    .I0(g35),
    .O(__1607__)
  );
  LUT5 #(
    .INIT(32'h00008000)
  ) __4988__ (
    .I4(__452__),
    .I3(__282__),
    .I2(__132__),
    .I1(__32__),
    .I0(__347__),
    .O(__1608__)
  );
  LUT5 #(
    .INIT(32'h000000f8)
  ) __4989__ (
    .I4(__19__),
    .I3(__1069__),
    .I2(g134),
    .I1(__884__),
    .I0(g99),
    .O(__1609__)
  );
  LUT6 #(
    .INIT(64'hccccf0aaf0f0f0f0)
  ) __4990__ (
    .I5(g35),
    .I4(__1609__),
    .I3(__1608__),
    .I2(__577__),
    .I1(__515__),
    .I0(__1179__),
    .O(__1610__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __4991__ (
    .I1(__253__),
    .I0(__689__),
    .O(__1611__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __4992__ (
    .I1(__357__),
    .I0(__613__),
    .O(__1612__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __4993__ (
    .I5(g35),
    .I4(__1612__),
    .I3(__1611__),
    .I2(__805__),
    .I1(__430__),
    .I0(__1391__),
    .O(__1613__)
  );
  LUT6 #(
    .INIT(64'h7dddddddf0f0f0f0)
  ) __4994__ (
    .I5(g35),
    .I4(__795__),
    .I3(__718__),
    .I2(__465__),
    .I1(__842__),
    .I0(__650__),
    .O(__1614__)
  );
  LUT3 #(
    .INIT(8'h01)
  ) __4995__ (
    .I2(__757__),
    .I1(__605__),
    .I0(__810__),
    .O(__1615__)
  );
  LUT6 #(
    .INIT(64'h0000000000000008)
  ) __4996__ (
    .I5(__445__),
    .I4(__519__),
    .I3(__1224__),
    .I2(__614__),
    .I1(__1190__),
    .I0(__1615__),
    .O(__1616__)
  );
  LUT5 #(
    .INIT(32'hccaaf0f0)
  ) __4997__ (
    .I4(g35),
    .I3(__1616__),
    .I2(__94__),
    .I1(__1108__),
    .I0(__1065__),
    .O(__1617__)
  );
  LUT4 #(
    .INIT(16'h7580)
  ) __4998__ (
    .I3(__182__),
    .I2(__1541__),
    .I1(__387__),
    .I0(g35),
    .O(__1618__)
  );
  LUT5 #(
    .INIT(32'hdddddfff)
  ) __4999__ (
    .I4(g134),
    .I3(__884__),
    .I2(g99),
    .I1(__701__),
    .I0(__1257__),
    .O(__1619__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __5000__ (
    .I1(__509__),
    .I0(__705__),
    .O(__1620__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5001__ (
    .I1(__463__),
    .I0(__120__),
    .O(__1621__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5002__ (
    .I5(g35),
    .I4(__1621__),
    .I3(__1620__),
    .I2(__615__),
    .I1(__517__),
    .I0(__1391__),
    .O(__1622__)
  );
  LUT6 #(
    .INIT(64'h00ff33330f0f5555)
  ) __5003__ (
    .I5(__465__),
    .I4(__842__),
    .I3(__38__),
    .I2(__864__),
    .I1(__503__),
    .I0(__1000__),
    .O(__1623__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5004__ (
    .I5(g35),
    .I4(__712__),
    .I3(__956__),
    .I2(__294__),
    .I1(__280__),
    .I0(__466__),
    .O(__1624__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __5005__ (
    .I1(__962__),
    .I0(__1034__),
    .O(__1625__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5006__ (
    .I5(g35),
    .I4(__1145__),
    .I3(__1625__),
    .I2(__634__),
    .I1(__852__),
    .I0(__1391__),
    .O(__1626__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5007__ (
    .I1(__351__),
    .I0(__1040__),
    .O(__1627__)
  );
  LUT6 #(
    .INIT(64'h007f00ffffff0000)
  ) __5008__ (
    .I5(g35),
    .I4(__376__),
    .I3(__729__),
    .I2(__1123__),
    .I1(__1074__),
    .I0(__1627__),
    .O(__1628__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5009__ (
    .I1(g35),
    .I0(__441__),
    .O(__1629__)
  );
  LUT6 #(
    .INIT(64'hefffffff00000000)
  ) __5010__ (
    .I5(__747__),
    .I4(__1310__),
    .I3(__1309__),
    .I2(__39__),
    .I1(__69__),
    .I0(__1077__),
    .O(__1630__)
  );
  LUT6 #(
    .INIT(64'h0077ff00f0f0f0f0)
  ) __5011__ (
    .I5(g35),
    .I4(__1630__),
    .I3(__254__),
    .I2(__729__),
    .I1(__1338__),
    .I0(__1569__),
    .O(__1631__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __5012__ (
    .I1(__468__),
    .I0(__704__),
    .O(__1632__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5013__ (
    .I1(__832__),
    .I0(__791__),
    .O(__1633__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5014__ (
    .I5(g35),
    .I4(__1633__),
    .I3(__1632__),
    .I2(__556__),
    .I1(__909__),
    .I0(__1391__),
    .O(__1634__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __5015__ (
    .I2(g35),
    .I1(__816__),
    .I0(__619__),
    .O(__1635__)
  );
  LUT4 #(
    .INIT(16'hef00)
  ) __5016__ (
    .I3(__878__),
    .I2(__1345__),
    .I1(__881__),
    .I0(__660__),
    .O(__1636__)
  );
  LUT2 #(
    .INIT(4'h2)
  ) __5017__ (
    .I1(__1118__),
    .I0(__1022__),
    .O(__1637__)
  );
  LUT6 #(
    .INIT(64'h000000000000007f)
  ) __5018__ (
    .I5(__1342__),
    .I4(__1637__),
    .I3(__1636__),
    .I2(__493__),
    .I1(__65__),
    .I0(__895__),
    .O(__1638__)
  );
  LUT6 #(
    .INIT(64'haaaaaaaccccccccc)
  ) __5019__ (
    .I5(g35),
    .I4(__1269__),
    .I3(__1638__),
    .I2(__318__),
    .I1(__1238__),
    .I0(__225__),
    .O(__1639__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5020__ (
    .I1(__179__),
    .I0(__801__),
    .O(__1640__)
  );
  LUT6 #(
    .INIT(64'hf055f0f0cccccccc)
  ) __5021__ (
    .I5(g35),
    .I4(__1640__),
    .I3(__1348__),
    .I2(__78__),
    .I1(__1023__),
    .I0(__1344__),
    .O(__1641__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5022__ (
    .I1(__1208__),
    .I0(__958__),
    .O(__1642__)
  );
  LUT6 #(
    .INIT(64'h000000000000fff4)
  ) __5023__ (
    .I5(__795__),
    .I4(__718__),
    .I3(__465__),
    .I2(__842__),
    .I1(__1285__),
    .I0(__9__),
    .O(__1643__)
  );
  LUT6 #(
    .INIT(64'h3caaaaaaf0f0f0f0)
  ) __5024__ (
    .I5(g35),
    .I4(__1643__),
    .I3(__1642__),
    .I2(__1152__),
    .I1(__1139__),
    .I0(__745__),
    .O(__1644__)
  );
  LUT6 #(
    .INIT(64'heaaa2aaaffff0000)
  ) __5025__ (
    .I5(g35),
    .I4(__271__),
    .I3(__468__),
    .I2(__704__),
    .I1(__898__),
    .I0(__490__),
    .O(__1645__)
  );
  LUT3 #(
    .INIT(8'h35)
  ) __5026__ (
    .I2(__949__),
    .I1(__843__),
    .I0(__446__),
    .O(__1646__)
  );
  LUT6 #(
    .INIT(64'h0300000305000005)
  ) __5027__ (
    .I5(__949__),
    .I4(__942__),
    .I3(__1646__),
    .I2(__1249__),
    .I1(__495__),
    .I0(__1183__),
    .O(__1647__)
  );
  LUT5 #(
    .INIT(32'h330f0f55)
  ) __5028__ (
    .I4(__700__),
    .I3(__949__),
    .I2(__159__),
    .I1(__184__),
    .I0(__996__),
    .O(__1648__)
  );
  LUT4 #(
    .INIT(16'h0080)
  ) __5029__ (
    .I3(__1251__),
    .I2(__1043__),
    .I1(__1110__),
    .I0(__547__),
    .O(__1649__)
  );
  LUT4 #(
    .INIT(16'h3e00)
  ) __5030__ (
    .I3(__1649__),
    .I2(__237__),
    .I1(__1648__),
    .I0(__1647__),
    .O(__1650__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __5031__ (
    .I2(__1110__),
    .I1(__1251__),
    .I0(__547__),
    .O(__1651__)
  );
  LUT6 #(
    .INIT(64'h0000f4ff00ff00ff)
  ) __5032__ (
    .I5(__188__),
    .I4(__315__),
    .I3(__891__),
    .I2(__1651__),
    .I1(__1650__),
    .I0(__758__),
    .O(__1652__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __5033__ (
    .I2(g35),
    .I1(__1652__),
    .I0(__1046__),
    .O(__1653__)
  );
  LUT5 #(
    .INIT(32'hbf80aaaa)
  ) __5034__ (
    .I4(g35),
    .I3(__622__),
    .I2(__1311__),
    .I1(__1319__),
    .I0(__1223__),
    .O(__1654__)
  );
  LUT5 #(
    .INIT(32'h3fc0aaaa)
  ) __5035__ (
    .I4(g35),
    .I3(__516__),
    .I2(__1311__),
    .I1(__1319__),
    .I0(__846__),
    .O(__1655__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __5036__ (
    .I1(__661__),
    .I0(__259__),
    .O(__1656__)
  );
  LUT6 #(
    .INIT(64'h0a03000000000000)
  ) __5037__ (
    .I5(g35),
    .I4(__1656__),
    .I3(__45__),
    .I2(__442__),
    .I1(__160__),
    .I0(__502__),
    .O(__1657__)
  );
  LUT6 #(
    .INIT(64'h00dfdf00ffff0000)
  ) __5038__ (
    .I5(g35),
    .I4(__457__),
    .I3(__1264__),
    .I2(__1303__),
    .I1(__810__),
    .I0(__1294__),
    .O(__1658__)
  );
  LUT6 #(
    .INIT(64'heaaa2aaaffff0000)
  ) __5039__ (
    .I5(g35),
    .I4(__60__),
    .I3(__157__),
    .I2(__561__),
    .I1(__863__),
    .I0(__1198__),
    .O(__1659__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5040__ (
    .I1(__509__),
    .I0(__705__),
    .O(__1660__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5041__ (
    .I5(g35),
    .I4(__1621__),
    .I3(__1660__),
    .I2(__1185__),
    .I1(__24__),
    .I0(__1391__),
    .O(__1661__)
  );
  LUT6 #(
    .INIT(64'h8000000000000000)
  ) __5042__ (
    .I5(__1004__),
    .I4(__1147__),
    .I3(__637__),
    .I2(__914__),
    .I1(__342__),
    .I0(__564__),
    .O(__1662__)
  );
  LUT4 #(
    .INIT(16'h8000)
  ) __5043__ (
    .I3(__592__),
    .I2(__890__),
    .I1(__1662__),
    .I0(__496__),
    .O(__1663__)
  );
  LUT5 #(
    .INIT(32'h0af0cccc)
  ) __5044__ (
    .I4(g35),
    .I3(__997__),
    .I2(__1663__),
    .I1(__496__),
    .I0(__1147__),
    .O(__1664__)
  );
  LUT6 #(
    .INIT(64'h8000000000000000)
  ) __5045__ (
    .I5(__606__),
    .I4(__214__),
    .I3(__719__),
    .I2(__546__),
    .I1(__285__),
    .I0(__1117__),
    .O(__1665__)
  );
  LUT6 #(
    .INIT(64'h7f33b3b3cc000000)
  ) __5046__ (
    .I5(__197__),
    .I4(__211__),
    .I3(__214__),
    .I2(__777__),
    .I1(g35),
    .I0(__1665__),
    .O(__1666__)
  );
  LUT5 #(
    .INIT(32'h00000080)
  ) __5047__ (
    .I4(g113),
    .I3(__1283__),
    .I2(__972__),
    .I1(__1446__),
    .I0(__1459__),
    .O(__1667__)
  );
  LUT6 #(
    .INIT(64'hf30caaaaf0f0f0f0)
  ) __5048__ (
    .I5(g35),
    .I4(__1667__),
    .I3(__749__),
    .I2(__469__),
    .I1(__784__),
    .I0(__1201__),
    .O(__1668__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __5049__ (
    .I2(g35),
    .I1(__223__),
    .I0(__232__),
    .O(__1669__)
  );
  LUT6 #(
    .INIT(64'h0000000000008421)
  ) __5050__ (
    .I5(__757__),
    .I4(__605__),
    .I3(g72),
    .I2(g73),
    .I1(__629__),
    .I0(__664__),
    .O(__1670__)
  );
  LUT6 #(
    .INIT(64'h06666666aaaaaaaa)
  ) __5051__ (
    .I5(g35),
    .I4(__1303__),
    .I3(__810__),
    .I2(__1670__),
    .I1(__357__),
    .I0(__613__),
    .O(__1671__)
  );
  LUT6 #(
    .INIT(64'h0000000000008000)
  ) __5052__ (
    .I5(__32__),
    .I4(__452__),
    .I3(__1235__),
    .I2(__153__),
    .I1(__347__),
    .I0(__203__),
    .O(__1672__)
  );
  LUT5 #(
    .INIT(32'hbfff0000)
  ) __5053__ (
    .I4(__52__),
    .I3(__282__),
    .I2(__374__),
    .I1(__1672__),
    .I0(__132__),
    .O(__1673__)
  );
  LUT4 #(
    .INIT(16'h8000)
  ) __5054__ (
    .I3(__359__),
    .I2(__1187__),
    .I1(__511__),
    .I0(__820__),
    .O(__1674__)
  );
  LUT5 #(
    .INIT(32'h3fc0aaaa)
  ) __5055__ (
    .I4(g35),
    .I3(__60__),
    .I2(__1674__),
    .I1(__1673__),
    .I0(__167__),
    .O(__1675__)
  );
  LUT5 #(
    .INIT(32'h00cef0f0)
  ) __5056__ (
    .I4(g35),
    .I3(__542__),
    .I2(__586__),
    .I1(__362__),
    .I0(__128__),
    .O(__1676__)
  );
  LUT3 #(
    .INIT(8'h08)
  ) __5057__ (
    .I2(__1236__),
    .I1(__1440__),
    .I0(__1052__),
    .O(__1677__)
  );
  LUT6 #(
    .INIT(64'hbfffffff00000000)
  ) __5058__ (
    .I5(__640__),
    .I4(__1310__),
    .I3(__1077__),
    .I2(__1309__),
    .I1(__222__),
    .I0(__69__),
    .O(__1678__)
  );
  LUT6 #(
    .INIT(64'h0077ff00f0f0f0f0)
  ) __5059__ (
    .I5(g35),
    .I4(__1678__),
    .I3(__1211__),
    .I2(__471__),
    .I1(__1338__),
    .I0(__1677__),
    .O(__1679__)
  );
  LUT6 #(
    .INIT(64'h0305000000000000)
  ) __5060__ (
    .I5(__11__),
    .I4(__492__),
    .I3(g84),
    .I2(__1193__),
    .I1(__143__),
    .I0(__246__),
    .O(__1680__)
  );
  LUT6 #(
    .INIT(64'h0c0a000000000000)
  ) __5061__ (
    .I5(__1193__),
    .I4(__959__),
    .I3(g84),
    .I2(__11__),
    .I1(__143__),
    .I0(__246__),
    .O(__1681__)
  );
  LUT6 #(
    .INIT(64'h00110c1cf0f0f0f0)
  ) __5062__ (
    .I5(g35),
    .I4(__959__),
    .I3(__1681__),
    .I2(__492__),
    .I1(__1205__),
    .I0(__1680__),
    .O(__1682__)
  );
  LUT6 #(
    .INIT(64'h06666666aaaaaaaa)
  ) __5063__ (
    .I5(g35),
    .I4(__1303__),
    .I3(__810__),
    .I2(__1302__),
    .I1(__548__),
    .I0(__566__),
    .O(__1683__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5064__ (
    .I1(__901__),
    .I0(__68__),
    .O(__1684__)
  );
  LUT6 #(
    .INIT(64'h7fffffff00000000)
  ) __5065__ (
    .I5(__12__),
    .I4(g35),
    .I3(__723__),
    .I2(__518__),
    .I1(__816__),
    .I0(__1684__),
    .O(__1685__)
  );
  LUT5 #(
    .INIT(32'hc3aaf0f0)
  ) __5066__ (
    .I4(g35),
    .I3(__1525__),
    .I2(__1244__),
    .I1(__516__),
    .I0(__1133__),
    .O(__1686__)
  );
  LUT4 #(
    .INIT(16'h8000)
  ) __5067__ (
    .I3(__1087__),
    .I2(__682__),
    .I1(__140__),
    .I0(__524__),
    .O(__1687__)
  );
  LUT5 #(
    .INIT(32'hfefeff00)
  ) __5068__ (
    .I4(__341__),
    .I3(__1165__),
    .I2(g72),
    .I1(g73),
    .I0(__1280__),
    .O(__1688__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __5069__ (
    .I1(g72),
    .I0(g73),
    .O(__1689__)
  );
  LUT6 #(
    .INIT(64'heeeef0f0ff00ff00)
  ) __5070__ (
    .I5(g35),
    .I4(__1689__),
    .I3(__682__),
    .I2(__1688__),
    .I1(__1687__),
    .I0(__796__),
    .O(__1690__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5071__ (
    .I1(g35),
    .I0(__569__),
    .O(__1691__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5072__ (
    .I1(__874__),
    .I0(__1264__),
    .O(__1692__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5073__ (
    .I5(g35),
    .I4(__457__),
    .I3(__1692__),
    .I2(__37__),
    .I1(__144__),
    .I0(__1391__),
    .O(__1693__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __5074__ (
    .I2(__507__),
    .I1(__1032__),
    .I0(__709__),
    .O(__1694__)
  );
  LUT6 #(
    .INIT(64'hdfff7555aaaa0000)
  ) __5075__ (
    .I5(__731__),
    .I4(__245__),
    .I3(__1694__),
    .I2(__88__),
    .I1(__835__),
    .I0(g35),
    .O(__1695__)
  );
  LUT5 #(
    .INIT(32'h0000f800)
  ) __5076__ (
    .I4(g113),
    .I3(__15__),
    .I2(g134),
    .I1(__884__),
    .I0(g99),
    .O(__1696__)
  );
  LUT6 #(
    .INIT(64'h0000000082000082)
  ) __5077__ (
    .I5(__1240__),
    .I4(g72),
    .I3(__976__),
    .I2(g73),
    .I1(__738__),
    .I0(__1696__),
    .O(__1697__)
  );
  LUT4 #(
    .INIT(16'h8000)
  ) __5078__ (
    .I3(__1235__),
    .I2(__203__),
    .I1(__153__),
    .I0(__706__),
    .O(__1698__)
  );
  LUT6 #(
    .INIT(64'h0000000000000004)
  ) __5079__ (
    .I5(__1698__),
    .I4(__1697__),
    .I3(__52__),
    .I2(__124__),
    .I1(g35),
    .I0(__21__),
    .O(__1699__)
  );
  LUT3 #(
    .INIT(8'h01)
  ) __5080__ (
    .I2(__364__),
    .I1(__321__),
    .I0(__646__),
    .O(__1700__)
  );
  LUT6 #(
    .INIT(64'h0000000000000580)
  ) __5081__ (
    .I5(__1207__),
    .I4(__936__),
    .I3(__544__),
    .I2(__396__),
    .I1(__646__),
    .I0(__262__),
    .O(__1701__)
  );
  LUT6 #(
    .INIT(64'hfcff0300aaaaaaaa)
  ) __5082__ (
    .I5(g35),
    .I4(__1701__),
    .I3(__1700__),
    .I2(__709__),
    .I1(__802__),
    .I0(__396__),
    .O(__1702__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5083__ (
    .I1(g35),
    .I0(__962__),
    .O(__1703__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5084__ (
    .I1(__688__),
    .I0(__636__),
    .O(__1704__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5085__ (
    .I5(g35),
    .I4(__1692__),
    .I3(__1704__),
    .I2(__144__),
    .I1(__948__),
    .I0(__1391__),
    .O(__1705__)
  );
  LUT6 #(
    .INIT(64'hfffc0003aaaaaaaa)
  ) __5086__ (
    .I5(g35),
    .I4(__850__),
    .I3(__196__),
    .I2(__1028__),
    .I1(__1489__),
    .I0(__697__),
    .O(__1706__)
  );
  LUT5 #(
    .INIT(32'h00000080)
  ) __5087__ (
    .I4(__917__),
    .I3(__353__),
    .I2(__972__),
    .I1(__1444__),
    .I0(__1443__),
    .O(__1707__)
  );
  LUT6 #(
    .INIT(64'h00000000fff40000)
  ) __5088__ (
    .I5(__795__),
    .I4(__718__),
    .I3(__465__),
    .I2(__842__),
    .I1(__1285__),
    .I0(__1158__),
    .O(__1708__)
  );
  LUT6 #(
    .INIT(64'heeeef0f0ff00ff00)
  ) __5089__ (
    .I5(g35),
    .I4(__1708__),
    .I3(__174__),
    .I2(__1237__),
    .I1(__934__),
    .I0(__1707__),
    .O(__1709__)
  );
  LUT5 #(
    .INIT(32'h00000008)
  ) __5090__ (
    .I4(__972__),
    .I3(g113),
    .I2(__1283__),
    .I1(__749__),
    .I0(__1298__),
    .O(__1710__)
  );
  LUT5 #(
    .INIT(32'hffa0cfc0)
  ) __5091__ (
    .I4(__1299__),
    .I3(__1197__),
    .I2(g35),
    .I1(__760__),
    .I0(__1710__),
    .O(__1711__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5092__ (
    .I1(__548__),
    .I0(__566__),
    .O(__1712__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5093__ (
    .I5(g35),
    .I4(__1712__),
    .I3(__1416__),
    .I2(__849__),
    .I1(__782__),
    .I0(__1391__),
    .O(__1713__)
  );
  LUT3 #(
    .INIT(8'h2c)
  ) __5094__ (
    .I2(g35),
    .I1(__912__),
    .I0(__66__),
    .O(__1714__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5095__ (
    .I1(__962__),
    .I0(__1034__),
    .O(__1715__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5096__ (
    .I5(g35),
    .I4(__1558__),
    .I3(__1715__),
    .I2(__856__),
    .I1(__703__),
    .I0(__1391__),
    .O(__1716__)
  );
  LUT4 #(
    .INIT(16'h8000)
  ) __5097__ (
    .I3(__917__),
    .I2(__972__),
    .I1(__1444__),
    .I0(__1282__),
    .O(__1717__)
  );
  LUT6 #(
    .INIT(64'hfff4000000000000)
  ) __5098__ (
    .I5(__795__),
    .I4(__718__),
    .I3(__465__),
    .I2(__842__),
    .I1(__1285__),
    .I0(__38__),
    .O(__1718__)
  );
  LUT6 #(
    .INIT(64'heeeef0f0ff00ff00)
  ) __5099__ (
    .I5(g35),
    .I4(__1718__),
    .I3(__792__),
    .I2(__13__),
    .I1(__91__),
    .I0(__1717__),
    .O(__1719__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __5100__ (
    .I1(__1091__),
    .I0(__1058__),
    .O(__1720__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __5101__ (
    .I1(__1045__),
    .I0(__483__),
    .O(__1721__)
  );
  LUT6 #(
    .INIT(64'h0000000000000008)
  ) __5102__ (
    .I5(__1149__),
    .I4(__602__),
    .I3(__1274__),
    .I2(__534__),
    .I1(__1721__),
    .I0(__1720__),
    .O(__1722__)
  );
  LUT4 #(
    .INIT(16'h0001)
  ) __5103__ (
    .I3(__965__),
    .I2(__861__),
    .I1(__231__),
    .I0(__1026__),
    .O(__1723__)
  );
  LUT6 #(
    .INIT(64'hfffeffff00000000)
  ) __5104__ (
    .I5(g35),
    .I4(__1723__),
    .I3(__697__),
    .I2(__836__),
    .I1(__183__),
    .I0(__928__),
    .O(__1724__)
  );
  LUT2 #(
    .INIT(4'hb)
  ) __5105__ (
    .I1(__1724__),
    .I0(__1722__),
    .O(__1725__)
  );
  LUT6 #(
    .INIT(64'h0000007f00000000)
  ) __5106__ (
    .I5(g35),
    .I4(__306__),
    .I3(__120__),
    .I2(__1303__),
    .I1(__810__),
    .I0(__1294__),
    .O(__1726__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5107__ (
    .I1(__613__),
    .I0(__357__),
    .O(__1727__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5108__ (
    .I1(__253__),
    .I0(__689__),
    .O(__1728__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5109__ (
    .I5(g35),
    .I4(__1728__),
    .I3(__1727__),
    .I2(__686__),
    .I1(__135__),
    .I0(__1391__),
    .O(__1729__)
  );
  LUT3 #(
    .INIT(8'h01)
  ) __5110__ (
    .I2(__170__),
    .I1(__1085__),
    .I0(__736__),
    .O(__1730__)
  );
  LUT6 #(
    .INIT(64'h55df557500aa0000)
  ) __5111__ (
    .I5(__896__),
    .I4(__1019__),
    .I3(__631__),
    .I2(__214__),
    .I1(__1730__),
    .I0(g35),
    .O(__1731__)
  );
  LUT6 #(
    .INIT(64'h00003fff00001555)
  ) __5112__ (
    .I5(__1118__),
    .I4(__1342__),
    .I3(__493__),
    .I2(__65__),
    .I1(__895__),
    .I0(__1022__),
    .O(__1732__)
  );
  LUT6 #(
    .INIT(64'h88d8888888d888d8)
  ) __5113__ (
    .I5(__1022__),
    .I4(__1118__),
    .I3(__1342__),
    .I2(__1248__),
    .I1(__739__),
    .I0(__1732__),
    .O(__1733__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __5114__ (
    .I1(__1638__),
    .I0(__318__),
    .O(__1734__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5115__ (
    .I5(g35),
    .I4(__617__),
    .I3(__1734__),
    .I2(__839__),
    .I1(__1252__),
    .I0(__1733__),
    .O(__1735__)
  );
  LUT4 #(
    .INIT(16'h77f0)
  ) __5116__ (
    .I3(g35),
    .I2(__1165__),
    .I1(__341__),
    .I0(__327__),
    .O(__1736__)
  );
  LUT3 #(
    .INIT(8'he0)
  ) __5117__ (
    .I2(g35),
    .I1(__1121__),
    .I0(__478__),
    .O(__1737__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5118__ (
    .I1(__13__),
    .I0(__711__),
    .O(__1738__)
  );
  LUT6 #(
    .INIT(64'hc3aaaaaaf0f0f0f0)
  ) __5119__ (
    .I5(g35),
    .I4(__1738__),
    .I3(__1718__),
    .I2(__1140__),
    .I1(__460__),
    .I0(__1026__),
    .O(__1739__)
  );
  LUT5 #(
    .INIT(32'hefefff00)
  ) __5120__ (
    .I4(g35),
    .I3(__130__),
    .I2(__1722__),
    .I1(__1061__),
    .I0(__1724__),
    .O(__1740__)
  );
  LUT6 #(
    .INIT(64'h0000007f00000000)
  ) __5121__ (
    .I5(g35),
    .I4(__613__),
    .I3(__623__),
    .I2(__1303__),
    .I1(__810__),
    .I0(__1670__),
    .O(__1741__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5122__ (
    .I1(__509__),
    .I0(__705__),
    .O(__1742__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5123__ (
    .I1(__463__),
    .I0(__120__),
    .O(__1743__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5124__ (
    .I5(g35),
    .I4(__1743__),
    .I3(__1742__),
    .I2(__911__),
    .I1(__670__),
    .I0(__1391__),
    .O(__1744__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __5125__ (
    .I2(g35),
    .I1(__796__),
    .I0(__1012__),
    .O(__1745__)
  );
  LUT6 #(
    .INIT(64'hff07ffffffffffff)
  ) __5126__ (
    .I5(g113),
    .I4(__1567__),
    .I3(__1578__),
    .I2(g134),
    .I1(__884__),
    .I0(g99),
    .O(__1746__)
  );
  LUT6 #(
    .INIT(64'h000000ff0000efef)
  ) __5127__ (
    .I5(__1343__),
    .I4(__1348__),
    .I3(__804__),
    .I2(__1248__),
    .I1(__1347__),
    .I0(__1342__),
    .O(__1747__)
  );
  LUT6 #(
    .INIT(64'h6666666affff0000)
  ) __5128__ (
    .I5(g35),
    .I4(__728__),
    .I3(__1348__),
    .I2(__801__),
    .I1(__673__),
    .I0(__1747__),
    .O(__1748__)
  );
  LUT6 #(
    .INIT(64'h6c206c6cf0f0f0f0)
  ) __5129__ (
    .I5(g35),
    .I4(__751__),
    .I3(__869__),
    .I2(__764__),
    .I1(__880__),
    .I0(__1454__),
    .O(__1749__)
  );
  LUT6 #(
    .INIT(64'h0000000080000000)
  ) __5130__ (
    .I5(__465__),
    .I4(__842__),
    .I3(__1227__),
    .I2(__917__),
    .I1(__353__),
    .I0(__972__),
    .O(__1750__)
  );
  LUT5 #(
    .INIT(32'hccaa0f0f)
  ) __5131__ (
    .I4(__1750__),
    .I3(__1503__),
    .I2(__864__),
    .I1(__1098__),
    .I0(__278__),
    .O(__1751__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __5132__ (
    .I2(g35),
    .I1(__1751__),
    .I0(__38__),
    .O(__1752__)
  );
  LUT3 #(
    .INIT(8'h08)
  ) __5133__ (
    .I2(__342__),
    .I1(g35),
    .I0(__1147__),
    .O(__1753__)
  );
  LUT5 #(
    .INIT(32'h00000001)
  ) __5134__ (
    .I4(__1103__),
    .I3(__485__),
    .I2(__284__),
    .I1(__192__),
    .I0(__481__),
    .O(__1754__)
  );
  LUT6 #(
    .INIT(64'h0f00afaacccccccc)
  ) __5135__ (
    .I5(g35),
    .I4(__659__),
    .I3(__284__),
    .I2(__479__),
    .I1(__192__),
    .I0(__1754__),
    .O(__1755__)
  );
  LUT2 #(
    .INIT(4'h9)
  ) __5136__ (
    .I1(__427__),
    .I0(__479__),
    .O(__1756__)
  );
  LUT5 #(
    .INIT(32'h00000001)
  ) __5137__ (
    .I4(__320__),
    .I3(__239__),
    .I2(__427__),
    .I1(__685__),
    .I0(__967__),
    .O(__1757__)
  );
  LUT6 #(
    .INIT(64'h11110f0fff00ff00)
  ) __5138__ (
    .I5(g35),
    .I4(__1757__),
    .I3(__604__),
    .I2(__1756__),
    .I1(__659__),
    .I0(__1144__),
    .O(__1758__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __5139__ (
    .I2(__881__),
    .I1(__660__),
    .I0(__580__),
    .O(__1759__)
  );
  LUT6 #(
    .INIT(64'hdfff7555aaaa0000)
  ) __5140__ (
    .I5(__137__),
    .I4(__943__),
    .I3(__152__),
    .I2(__1759__),
    .I1(__985__),
    .I0(g35),
    .O(__1760__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5141__ (
    .I1(__1264__),
    .I0(__874__),
    .O(__1761__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5142__ (
    .I5(g35),
    .I4(__1761__),
    .I3(__1704__),
    .I2(__593__),
    .I1(__138__),
    .I0(__1391__),
    .O(__1762__)
  );
  LUT6 #(
    .INIT(64'h0000000000000008)
  ) __5143__ (
    .I5(__445__),
    .I4(__519__),
    .I3(__1224__),
    .I2(__1190__),
    .I1(__614__),
    .I0(__1615__),
    .O(__1763__)
  );
  LUT5 #(
    .INIT(32'hccaaf0f0)
  ) __5144__ (
    .I4(g35),
    .I3(__1763__),
    .I2(__1025__),
    .I1(__1108__),
    .I0(__94__),
    .O(__1764__)
  );
  LUT6 #(
    .INIT(64'h3fffc000aaaaaaaa)
  ) __5145__ (
    .I5(g35),
    .I4(__376__),
    .I3(__1123__),
    .I2(__1074__),
    .I1(__1627__),
    .I0(__920__),
    .O(__1765__)
  );
  LUT5 #(
    .INIT(32'h7fff0000)
  ) __5146__ (
    .I4(g35),
    .I3(__1043__),
    .I2(__1110__),
    .I1(__762__),
    .I0(__1251__),
    .O(__1766__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __5147__ (
    .I2(__1766__),
    .I1(__159__),
    .I0(__495__),
    .O(__1767__)
  );
  LUT6 #(
    .INIT(64'h77ff0800ff00ff00)
  ) __5148__ (
    .I5(g35),
    .I4(__1181__),
    .I3(__770__),
    .I2(__1072__),
    .I1(__1233__),
    .I0(__385__),
    .O(__1768__)
  );
  LUT6 #(
    .INIT(64'h5adaaa2affff0000)
  ) __5149__ (
    .I5(g35),
    .I4(__963__),
    .I3(__958__),
    .I2(__1643__),
    .I1(__1208__),
    .I0(__1152__),
    .O(__1769__)
  );
  LUT6 #(
    .INIT(64'h0000000000000001)
  ) __5150__ (
    .I5(__659__),
    .I4(__1103__),
    .I3(__485__),
    .I2(__284__),
    .I1(__192__),
    .I0(__481__),
    .O(__1770__)
  );
  LUT4 #(
    .INIT(16'hff80)
  ) __5151__ (
    .I3(__485__),
    .I2(g35),
    .I1(__337__),
    .I0(__1770__),
    .O(__1771__)
  );
  LUT4 #(
    .INIT(16'h7da0)
  ) __5152__ (
    .I3(__725__),
    .I2(__1095__),
    .I1(__734__),
    .I0(g35),
    .O(__1772__)
  );
  LUT6 #(
    .INIT(64'h0000000082410000)
  ) __5153__ (
    .I5(__605__),
    .I4(__757__),
    .I3(g72),
    .I2(g73),
    .I1(__664__),
    .I0(__629__),
    .O(__1773__)
  );
  LUT6 #(
    .INIT(64'h06666666aaaaaaaa)
  ) __5154__ (
    .I5(g35),
    .I4(__1773__),
    .I3(__1303__),
    .I2(__810__),
    .I1(__832__),
    .I0(__791__),
    .O(__1774__)
  );
  LUT6 #(
    .INIT(64'h0000000080000000)
  ) __5155__ (
    .I5(__794__),
    .I4(__1268__),
    .I3(__1052__),
    .I2(__1236__),
    .I1(__702__),
    .I0(__482__),
    .O(__1775__)
  );
  LUT6 #(
    .INIT(64'h44444444ccccc444)
  ) __5156__ (
    .I5(g113),
    .I4(g134),
    .I3(__884__),
    .I2(g99),
    .I1(__473__),
    .I0(__1689__),
    .O(__1776__)
  );
  LUT6 #(
    .INIT(64'h0000000022220888)
  ) __5157__ (
    .I5(__1776__),
    .I4(__1240__),
    .I3(__738__),
    .I2(__976__),
    .I1(__1775__),
    .I0(g35),
    .O(__1777__)
  );
  LUT5 #(
    .INIT(32'h0000f800)
  ) __5158__ (
    .I4(g113),
    .I3(__1060__),
    .I2(g134),
    .I1(__884__),
    .I0(g99),
    .O(__1778__)
  );
  LUT5 #(
    .INIT(32'h00008000)
  ) __5159__ (
    .I4(__639__),
    .I3(__1778__),
    .I2(__779__),
    .I1(__1414__),
    .I0(__845__),
    .O(__1779__)
  );
  LUT4 #(
    .INIT(16'hbf00)
  ) __5160__ (
    .I3(__380__),
    .I2(__1487__),
    .I1(__507__),
    .I0(__1032__),
    .O(__1780__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5161__ (
    .I1(__583__),
    .I0(__441__),
    .O(__1781__)
  );
  LUT6 #(
    .INIT(64'h00000000000000f7)
  ) __5162__ (
    .I5(__1485__),
    .I4(__1781__),
    .I3(__1780__),
    .I2(__1143__),
    .I1(__1186__),
    .I0(__961__),
    .O(__1782__)
  );
  LUT6 #(
    .INIT(64'hf0f04444ff00ff00)
  ) __5163__ (
    .I5(g35),
    .I4(__1782__),
    .I3(__753__),
    .I2(__908__),
    .I1(__860__),
    .I0(__1779__),
    .O(__1783__)
  );
  LUT4 #(
    .INIT(16'hcacc)
  ) __5164__ (
    .I3(g35),
    .I2(__1532__),
    .I1(__781__),
    .I0(__244__),
    .O(__1784__)
  );
  LUT6 #(
    .INIT(64'h0000f3ff00005155)
  ) __5165__ (
    .I5(__1118__),
    .I4(__1342__),
    .I3(__493__),
    .I2(__65__),
    .I1(__895__),
    .I0(__943__),
    .O(__1785__)
  );
  LUT6 #(
    .INIT(64'h0000ff000000efef)
  ) __5166__ (
    .I5(__1785__),
    .I4(__1521__),
    .I3(__804__),
    .I2(__1248__),
    .I1(__1342__),
    .I0(__1519__),
    .O(__1786__)
  );
  LUT6 #(
    .INIT(64'h6666666affff0000)
  ) __5167__ (
    .I5(g35),
    .I4(__595__),
    .I3(__112__),
    .I2(__1521__),
    .I1(__58__),
    .I0(__1786__),
    .O(__1787__)
  );
  LUT2 #(
    .INIT(4'h2)
  ) __5168__ (
    .I1(__869__),
    .I0(__751__),
    .O(__1788__)
  );
  LUT6 #(
    .INIT(64'h337fb3b300cc0000)
  ) __5169__ (
    .I5(__880__),
    .I4(__207__),
    .I3(__1788__),
    .I2(__764__),
    .I1(g35),
    .I0(__1454__),
    .O(__1789__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5170__ (
    .I1(__561__),
    .I0(__863__),
    .O(__1790__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5171__ (
    .I1(__267__),
    .I0(__425__),
    .O(__1791__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5172__ (
    .I5(g35),
    .I4(__1791__),
    .I3(__1790__),
    .I2(__324__),
    .I1(__905__),
    .I0(__1391__),
    .O(__1792__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5173__ (
    .I1(__569__),
    .I0(__313__),
    .O(__1793__)
  );
  LUT3 #(
    .INIT(8'h01)
  ) __5174__ (
    .I2(__989__),
    .I1(__418__),
    .I0(__1173__),
    .O(__1794__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5175__ (
    .I5(g35),
    .I4(__1794__),
    .I3(__1793__),
    .I2(__234__),
    .I1(__937__),
    .I0(__1391__),
    .O(__1795__)
  );
  LUT6 #(
    .INIT(64'hf0f04444ff00ff00)
  ) __5176__ (
    .I5(g35),
    .I4(__1489__),
    .I3(__1128__),
    .I2(__190__),
    .I1(__1028__),
    .I0(__1484__),
    .O(__1796__)
  );
  LUT5 #(
    .INIT(32'hc3aaf0f0)
  ) __5177__ (
    .I4(g35),
    .I3(__1493__),
    .I2(__625__),
    .I1(__630__),
    .I0(__292__),
    .O(__1797__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5178__ (
    .I1(__801__),
    .I0(__1348__),
    .O(__1798__)
  );
  LUT6 #(
    .INIT(64'hf055f0f0cccccccc)
  ) __5179__ (
    .I5(g35),
    .I4(__1798__),
    .I3(__179__),
    .I2(__506__),
    .I1(__1131__),
    .I0(__1344__),
    .O(__1799__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5180__ (
    .I1(__1014__),
    .I0(__950__),
    .O(__1800__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5181__ (
    .I1(__1208__),
    .I0(__191__),
    .O(__1801__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5182__ (
    .I5(g35),
    .I4(__1643__),
    .I3(__1801__),
    .I2(__41__),
    .I1(__1059__),
    .I0(__1800__),
    .O(__1802__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5183__ (
    .I1(__469__),
    .I0(__462__),
    .O(__1803__)
  );
  LUT6 #(
    .INIT(64'h3caaaaaaf0f0f0f0)
  ) __5184__ (
    .I5(g35),
    .I4(__1446__),
    .I3(__1803__),
    .I2(__108__),
    .I1(__273__),
    .I0(__322__),
    .O(__1804__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5185__ (
    .I1(__817__),
    .I0(__900__),
    .O(__1805__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5186__ (
    .I5(g35),
    .I4(__1417__),
    .I3(__1805__),
    .I2(__1259__),
    .I1(__1075__),
    .I0(__1391__),
    .O(__1806__)
  );
  LUT3 #(
    .INIT(8'h81)
  ) __5187__ (
    .I2(__584__),
    .I1(__244__),
    .I0(__77__),
    .O(__1807__)
  );
  LUT6 #(
    .INIT(64'h000d0d0d00000000)
  ) __5188__ (
    .I5(__1532__),
    .I4(__786__),
    .I3(__693__),
    .I2(__1807__),
    .I1(__973__),
    .I0(__28__),
    .O(__1808__)
  );
  LUT5 #(
    .INIT(32'h0dd0cccc)
  ) __5189__ (
    .I4(g35),
    .I3(__497__),
    .I2(__1808__),
    .I1(__279__),
    .I0(__973__),
    .O(__1809__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5190__ (
    .I1(__91__),
    .I0(__711__),
    .O(__1810__)
  );
  LUT6 #(
    .INIT(64'h3caaaaaaf0f0f0f0)
  ) __5191__ (
    .I5(g35),
    .I4(__1718__),
    .I3(__1810__),
    .I2(__708__),
    .I1(__332__),
    .I0(__470__),
    .O(__1811__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __5192__ (
    .I1(__544__),
    .I0(__396__),
    .O(__1812__)
  );
  LUT6 #(
    .INIT(64'h0000553f000000ff)
  ) __5193__ (
    .I5(__1207__),
    .I4(__936__),
    .I3(__1812__),
    .I2(__775__),
    .I1(__766__),
    .I0(__594__),
    .O(__1813__)
  );
  LUT6 #(
    .INIT(64'h0a380a38ffff0000)
  ) __5194__ (
    .I5(g35),
    .I4(__1207__),
    .I3(__544__),
    .I2(__1036__),
    .I1(__646__),
    .I0(__1813__),
    .O(__1814__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5195__ (
    .I5(g35),
    .I4(__1611__),
    .I3(__1727__),
    .I2(__761__),
    .I1(__405__),
    .I0(__1391__),
    .O(__1815__)
  );
  LUT6 #(
    .INIT(64'h000d000000000000)
  ) __5196__ (
    .I5(__1532__),
    .I4(__497__),
    .I3(__1530__),
    .I2(__1807__),
    .I1(__973__),
    .I0(__28__),
    .O(__1816__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5197__ (
    .I1(__973__),
    .I0(__279__),
    .O(__1817__)
  );
  LUT6 #(
    .INIT(64'h0000000080000000)
  ) __5198__ (
    .I5(__1817__),
    .I4(__633__),
    .I3(__126__),
    .I2(__587__),
    .I1(__175__),
    .I0(__1816__),
    .O(__1818__)
  );
  LUT6 #(
    .INIT(64'h8000000000000000)
  ) __5199__ (
    .I5(__252__),
    .I4(__1818__),
    .I3(__642__),
    .I2(__790__),
    .I1(__459__),
    .I0(__525__),
    .O(__1819__)
  );
  LUT6 #(
    .INIT(64'h557f55d500aa0000)
  ) __5200__ (
    .I5(__251__),
    .I4(__693__),
    .I3(__1817__),
    .I2(__1078__),
    .I1(__1819__),
    .I0(g35),
    .O(__1820__)
  );
  LUT6 #(
    .INIT(64'heaaa2aaaffff0000)
  ) __5201__ (
    .I5(g35),
    .I4(__539__),
    .I3(__253__),
    .I2(__689__),
    .I1(__623__),
    .I0(__240__),
    .O(__1821__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __5202__ (
    .I2(g35),
    .I1(__938__),
    .I0(__789__),
    .O(__1822__)
  );
  LUT3 #(
    .INIT(8'h01)
  ) __5203__ (
    .I2(__306__),
    .I1(__463__),
    .I0(__120__),
    .O(__1823__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5204__ (
    .I5(g35),
    .I4(__1823__),
    .I3(__1742__),
    .I2(__421__),
    .I1(__1137__),
    .I0(__1391__),
    .O(__1824__)
  );
  LUT5 #(
    .INIT(32'h7d55a000)
  ) __5205__ (
    .I4(__1227__),
    .I3(__650__),
    .I2(__972__),
    .I1(__1462__),
    .I0(g35),
    .O(__1825__)
  );
  LUT6 #(
    .INIT(64'hfffc0003aaaaaaaa)
  ) __5206__ (
    .I5(g35),
    .I4(__931__),
    .I3(__860__),
    .I2(__1111__),
    .I1(__1782__),
    .I0(__861__),
    .O(__1826__)
  );
  LUT6 #(
    .INIT(64'h0a0a5f0a0a0a1b0a)
  ) __5207__ (
    .I5(__1118__),
    .I4(__1342__),
    .I3(__1248__),
    .I2(__739__),
    .I1(__943__),
    .I0(__1785__),
    .O(__1827__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5208__ (
    .I1(__595__),
    .I0(__1521__),
    .O(__1828__)
  );
  LUT6 #(
    .INIT(64'hf055f0f0cccccccc)
  ) __5209__ (
    .I5(g35),
    .I4(__1828__),
    .I3(__540__),
    .I2(__26__),
    .I1(__1277__),
    .I0(__1827__),
    .O(__1829__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5210__ (
    .I1(__934__),
    .I0(__653__),
    .O(__1830__)
  );
  LUT6 #(
    .INIT(64'h3caaaaaaf0f0f0f0)
  ) __5211__ (
    .I5(g35),
    .I4(__1708__),
    .I3(__1830__),
    .I2(__894__),
    .I1(__1001__),
    .I0(__947__),
    .O(__1831__)
  );
  LUT6 #(
    .INIT(64'h0000553f000000ff)
  ) __5212__ (
    .I5(__437__),
    .I4(__35__),
    .I3(__1398__),
    .I2(__413__),
    .I1(__116__),
    .I0(__1029__),
    .O(__1832__)
  );
  LUT6 #(
    .INIT(64'h0a380a38ffff0000)
  ) __5213__ (
    .I5(g35),
    .I4(__437__),
    .I3(__631__),
    .I2(__555__),
    .I1(__736__),
    .I0(__1832__),
    .O(__1833__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __5214__ (
    .I2(g35),
    .I1(g64),
    .I0(__244__),
    .O(__1834__)
  );
  LUT6 #(
    .INIT(64'h0000000000008000)
  ) __5215__ (
    .I5(g113),
    .I4(__1283__),
    .I3(__757__),
    .I2(__1385__),
    .I1(__236__),
    .I0(__810__),
    .O(__1835__)
  );
  LUT5 #(
    .INIT(32'h575d0a00)
  ) __5216__ (
    .I4(__704__),
    .I3(__468__),
    .I2(__1835__),
    .I1(__898__),
    .I0(g35),
    .O(__1836__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5217__ (
    .I1(__798__),
    .I0(__386__),
    .O(__1837__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5218__ (
    .I5(g35),
    .I4(__1837__),
    .I3(__1394__),
    .I2(__1163__),
    .I1(__574__),
    .I0(__1391__),
    .O(__1838__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __5219__ (
    .I1(__141__),
    .I0(__812__),
    .O(__1839__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __5220__ (
    .I1(__984__),
    .I0(__980__),
    .O(__1840__)
  );
  LUT6 #(
    .INIT(64'h0000000000000008)
  ) __5221__ (
    .I5(__907__),
    .I4(__651__),
    .I3(__174__),
    .I2(__957__),
    .I1(__1840__),
    .I0(__1839__),
    .O(__1841__)
  );
  LUT4 #(
    .INIT(16'h0001)
  ) __5222__ (
    .I3(__422__),
    .I2(__792__),
    .I1(__228__),
    .I0(__753__),
    .O(__1842__)
  );
  LUT6 #(
    .INIT(64'hfffeffff00000000)
  ) __5223__ (
    .I5(g35),
    .I4(__1842__),
    .I3(__1128__),
    .I2(__543__),
    .I1(__925__),
    .I0(__1201__),
    .O(__1843__)
  );
  LUT2 #(
    .INIT(4'hb)
  ) __5224__ (
    .I1(__1843__),
    .I0(__1841__),
    .O(__1844__)
  );
  LUT6 #(
    .INIT(64'heaaa2aaaffff0000)
  ) __5225__ (
    .I5(g35),
    .I4(__1024__),
    .I3(__157__),
    .I2(__561__),
    .I1(__863__),
    .I0(__787__),
    .O(__1845__)
  );
  LUT6 #(
    .INIT(64'heaaa2aaaffff0000)
  ) __5226__ (
    .I5(g35),
    .I4(__969__),
    .I3(__653__),
    .I2(__1237__),
    .I1(__1708__),
    .I0(__877__),
    .O(__1846__)
  );
  LUT4 #(
    .INIT(16'h8000)
  ) __5227__ (
    .I3(__1063__),
    .I2(__376__),
    .I1(__527__),
    .I0(__254__),
    .O(__1847__)
  );
  LUT5 #(
    .INIT(32'hbf80aaaa)
  ) __5228__ (
    .I4(g35),
    .I3(__258__),
    .I2(__1847__),
    .I1(__1630__),
    .I0(__235__),
    .O(__1848__)
  );
  LUT6 #(
    .INIT(64'h000000ff0000efef)
  ) __5229__ (
    .I5(__1551__),
    .I4(__1555__),
    .I3(__666__),
    .I2(__1248__),
    .I1(__1485__),
    .I0(__1553__),
    .O(__1849__)
  );
  LUT6 #(
    .INIT(64'h6666666affff0000)
  ) __5230__ (
    .I5(g35),
    .I4(__746__),
    .I3(__793__),
    .I2(__1555__),
    .I1(__855__),
    .I0(__1849__),
    .O(__1850__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __5231__ (
    .I2(g35),
    .I1(g6749),
    .I0(__524__),
    .O(__1851__)
  );
  LUT3 #(
    .INIT(8'h01)
  ) __5232__ (
    .I2(__412__),
    .I1(__566__),
    .I0(__548__),
    .O(__1852__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5233__ (
    .I1(__900__),
    .I0(__817__),
    .O(__1853__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5234__ (
    .I5(g35),
    .I4(__1853__),
    .I3(__1852__),
    .I2(__1246__),
    .I1(__1136__),
    .I0(__1391__),
    .O(__1854__)
  );
  LUT4 #(
    .INIT(16'h7da0)
  ) __5235__ (
    .I3(__585__),
    .I2(__652__),
    .I1(__1068__),
    .I0(g35),
    .O(__1855__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __5236__ (
    .I2(__1766__),
    .I1(__996__),
    .I0(__1183__),
    .O(__1856__)
  );
  LUT5 #(
    .INIT(32'h80000000)
  ) __5237__ (
    .I4(__151__),
    .I3(__926__),
    .I2(__995__),
    .I1(__1192__),
    .I0(__288__),
    .O(__1857__)
  );
  LUT6 #(
    .INIT(64'h112055a0f0f0f0f0)
  ) __5238__ (
    .I5(g35),
    .I4(__1440__),
    .I3(__788__),
    .I2(__721__),
    .I1(__1696__),
    .I0(__1857__),
    .O(__1858__)
  );
  LUT5 #(
    .INIT(32'h80000000)
  ) __5239__ (
    .I4(__1235__),
    .I3(__203__),
    .I2(__153__),
    .I1(__706__),
    .I0(__32__),
    .O(__1859__)
  );
  LUT6 #(
    .INIT(64'h00787878cccccccc)
  ) __5240__ (
    .I5(g35),
    .I4(__1696__),
    .I3(__1396__),
    .I2(__132__),
    .I1(__347__),
    .I0(__1859__),
    .O(__1860__)
  );
  LUT6 #(
    .INIT(64'heaaa2aaaffff0000)
  ) __5241__ (
    .I5(g35),
    .I4(__516__),
    .I3(__509__),
    .I2(__306__),
    .I1(__705__),
    .I0(__1244__),
    .O(__1861__)
  );
  LUT6 #(
    .INIT(64'h78f070f0ffff0000)
  ) __5242__ (
    .I5(g35),
    .I4(__1181__),
    .I3(__770__),
    .I2(__1072__),
    .I1(__1233__),
    .I0(__385__),
    .O(__1862__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5243__ (
    .I5(g35),
    .I4(__1852__),
    .I3(__1416__),
    .I2(__1086__),
    .I1(__1215__),
    .I0(__1391__),
    .O(__1863__)
  );
  LUT3 #(
    .INIT(8'h04)
  ) __5244__ (
    .I2(__188__),
    .I1(__315__),
    .I0(__891__),
    .O(__1864__)
  );
  LUT5 #(
    .INIT(32'hccaaf0f0)
  ) __5245__ (
    .I4(g35),
    .I3(__1864__),
    .I2(__34__),
    .I1(__528__),
    .I0(__198__),
    .O(__1865__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5246__ (
    .I1(__468__),
    .I0(__704__),
    .O(__1866__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5247__ (
    .I5(g35),
    .I4(__1866__),
    .I3(__898__),
    .I2(__194__),
    .I1(__1010__),
    .I0(__1391__),
    .O(__1867__)
  );
  LUT6 #(
    .INIT(64'heaaa2aaaffff0000)
  ) __5248__ (
    .I5(g35),
    .I4(__1073__),
    .I3(__509__),
    .I2(__306__),
    .I1(__705__),
    .I0(__754__),
    .O(__1868__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5249__ (
    .I1(__760__),
    .I0(__1197__),
    .O(__1869__)
  );
  LUT6 #(
    .INIT(64'h3caaaaaaf0f0f0f0)
  ) __5250__ (
    .I5(g35),
    .I4(__1299__),
    .I3(__1869__),
    .I2(__692__),
    .I1(__372__),
    .I0(__260__),
    .O(__1870__)
  );
  LUT4 #(
    .INIT(16'h8000)
  ) __5251__ (
    .I3(__738__),
    .I2(__976__),
    .I1(__1775__),
    .I0(__871__),
    .O(__1871__)
  );
  LUT4 #(
    .INIT(16'h8000)
  ) __5252__ (
    .I3(__343__),
    .I2(__114__),
    .I1(__92__),
    .I0(__1871__),
    .O(__1872__)
  );
  LUT6 #(
    .INIT(64'h00003a3aff00ff00)
  ) __5253__ (
    .I5(g35),
    .I4(__1776__),
    .I3(__92__),
    .I2(__301__),
    .I1(__1871__),
    .I0(__1872__),
    .O(__1873__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __5254__ (
    .I1(__313__),
    .I0(__569__),
    .O(__1874__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5255__ (
    .I5(g35),
    .I4(__989__),
    .I3(__1874__),
    .I2(__147__),
    .I1(__121__),
    .I0(__1391__),
    .O(__1875__)
  );
  LUT4 #(
    .INIT(16'h8000)
  ) __5256__ (
    .I3(__151__),
    .I2(__926__),
    .I1(__995__),
    .I0(__1192__),
    .O(__1876__)
  );
  LUT6 #(
    .INIT(64'h03300ff0aaaaaaaa)
  ) __5257__ (
    .I5(g35),
    .I4(__1440__),
    .I3(__1876__),
    .I2(__288__),
    .I1(__1696__),
    .I0(__1055__),
    .O(__1877__)
  );
  LUT6 #(
    .INIT(64'hbfffffff00000000)
  ) __5258__ (
    .I5(__124__),
    .I4(g35),
    .I3(__1503__),
    .I2(__1567__),
    .I1(__15__),
    .I0(__1240__),
    .O(__1878__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __5259__ (
    .I2(g35),
    .I1(__1187__),
    .I0(__227__),
    .O(__1879__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5260__ (
    .I1(__832__),
    .I0(__791__),
    .O(__1880__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5261__ (
    .I5(g35),
    .I4(__1880__),
    .I3(__1632__),
    .I2(__1229__),
    .I1(__556__),
    .I0(__1391__),
    .O(__1881__)
  );
  LUT6 #(
    .INIT(64'h13034c0caaaaaaaa)
  ) __5262__ (
    .I5(g35),
    .I4(__1451__),
    .I3(__875__),
    .I2(__671__),
    .I1(__265__),
    .I0(__177__),
    .O(__1882__)
  );
  LUT3 #(
    .INIT(8'h08)
  ) __5263__ (
    .I2(__1032__),
    .I1(__507__),
    .I0(__709__),
    .O(__1883__)
  );
  LUT6 #(
    .INIT(64'hdfff7555aaaa0000)
  ) __5264__ (
    .I5(__275__),
    .I4(__583__),
    .I3(__88__),
    .I2(__1883__),
    .I1(__835__),
    .I0(g35),
    .O(__1884__)
  );
  LUT4 #(
    .INIT(16'h8000)
  ) __5265__ (
    .I3(__115__),
    .I2(__612__),
    .I1(__394__),
    .I0(__873__),
    .O(__1885__)
  );
  LUT4 #(
    .INIT(16'h3caa)
  ) __5266__ (
    .I3(g35),
    .I2(__1187__),
    .I1(__1885__),
    .I0(__681__),
    .O(__1886__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5267__ (
    .I1(__944__),
    .I0(__1600__),
    .O(__1887__)
  );
  LUT6 #(
    .INIT(64'hf055f0f0cccccccc)
  ) __5268__ (
    .I5(g35),
    .I4(__1887__),
    .I3(__1027__),
    .I2(__1021__),
    .I1(__927__),
    .I0(__1597__),
    .O(__1888__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5269__ (
    .I5(g35),
    .I4(__296__),
    .I3(__1887__),
    .I2(__923__),
    .I1(__70__),
    .I0(__1597__),
    .O(__1889__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __5270__ (
    .I2(__770__),
    .I1(__1233__),
    .I0(__385__),
    .O(__1890__)
  );
  LUT5 #(
    .INIT(32'h0000002c)
  ) __5271__ (
    .I4(__1207__),
    .I3(__936__),
    .I2(__396__),
    .I1(__544__),
    .I0(__646__),
    .O(__1891__)
  );
  LUT6 #(
    .INIT(64'h00000000000000f7)
  ) __5272__ (
    .I5(__998__),
    .I4(__380__),
    .I3(__674__),
    .I2(__1891__),
    .I1(__1072__),
    .I0(__1890__),
    .O(__1892__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5273__ (
    .I1(g35),
    .I0(__1892__),
    .O(__1893__)
  );
  LUT5 #(
    .INIT(32'h00000008)
  ) __5274__ (
    .I4(g113),
    .I3(__1283__),
    .I2(__810__),
    .I1(__1773__),
    .I0(__236__),
    .O(__1894__)
  );
  LUT5 #(
    .INIT(32'h575d0a00)
  ) __5275__ (
    .I4(__863__),
    .I3(__561__),
    .I2(__1894__),
    .I1(__157__),
    .I0(g35),
    .O(__1895__)
  );
  LUT5 #(
    .INIT(32'hefff0000)
  ) __5276__ (
    .I4(__21__),
    .I3(__1672__),
    .I2(__1179__),
    .I1(__282__),
    .I0(__132__),
    .O(__1896__)
  );
  LUT5 #(
    .INIT(32'h80000000)
  ) __5277__ (
    .I4(__847__),
    .I3(__870__),
    .I2(__648__),
    .I1(__1896__),
    .I0(__155__),
    .O(__1897__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5278__ (
    .I1(__870__),
    .I0(__648__),
    .O(__1898__)
  );
  LUT6 #(
    .INIT(64'h0fffffffffff7777)
  ) __5279__ (
    .I5(__870__),
    .I4(__648__),
    .I3(__565__),
    .I2(__724__),
    .I1(__1262__),
    .I0(__759__),
    .O(__1899__)
  );
  LUT6 #(
    .INIT(64'h7f00000000007f00)
  ) __5280__ (
    .I5(__847__),
    .I4(__379__),
    .I3(__1899__),
    .I2(__474__),
    .I1(__1898__),
    .I0(__1064__),
    .O(__1900__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5281__ (
    .I1(__648__),
    .I0(__870__),
    .O(__1901__)
  );
  LUT6 #(
    .INIT(64'hffff0fffffff7777)
  ) __5282__ (
    .I5(__870__),
    .I4(__648__),
    .I3(__109__),
    .I2(__759__),
    .I1(__474__),
    .I0(__47__),
    .O(__1902__)
  );
  LUT6 #(
    .INIT(64'h00007f007f000000)
  ) __5283__ (
    .I5(__847__),
    .I4(__379__),
    .I3(__1902__),
    .I2(__724__),
    .I1(__1901__),
    .I0(__986__),
    .O(__1903__)
  );
  LUT4 #(
    .INIT(16'h8000)
  ) __5284__ (
    .I3(__847__),
    .I2(__870__),
    .I1(__648__),
    .I0(__155__),
    .O(__1904__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5285__ (
    .I1(__208__),
    .I0(__513__),
    .O(__1905__)
  );
  LUT6 #(
    .INIT(64'h007f7f7f00000000)
  ) __5286__ (
    .I5(__847__),
    .I4(__1898__),
    .I3(__1905__),
    .I2(__181__),
    .I1(__1566__),
    .I0(__121__),
    .O(__1906__)
  );
  LUT6 #(
    .INIT(64'h000000f800000088)
  ) __5287__ (
    .I5(__122__),
    .I4(__870__),
    .I3(__648__),
    .I2(__598__),
    .I1(__885__),
    .I0(__147__),
    .O(__1907__)
  );
  LUT6 #(
    .INIT(64'h000007770000ffff)
  ) __5288__ (
    .I5(__1901__),
    .I4(__1907__),
    .I3(__133__),
    .I2(__601__),
    .I1(__379__),
    .I0(__1191__),
    .O(__1908__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __5289__ (
    .I1(__870__),
    .I0(__648__),
    .O(__1909__)
  );
  LUT6 #(
    .INIT(64'h0000f88800000000)
  ) __5290__ (
    .I5(__870__),
    .I4(__648__),
    .I3(__122__),
    .I2(__234__),
    .I1(__885__),
    .I0(__883__),
    .O(__1910__)
  );
  LUT6 #(
    .INIT(64'h0000f88800000000)
  ) __5291__ (
    .I5(__648__),
    .I4(__870__),
    .I3(__181__),
    .I2(__570__),
    .I1(__155__),
    .I0(__937__),
    .O(__1911__)
  );
  LUT6 #(
    .INIT(64'h000007770000ffff)
  ) __5292__ (
    .I5(__1566__),
    .I4(__1911__),
    .I3(__133__),
    .I2(__807__),
    .I1(__379__),
    .I0(__808__),
    .O(__1912__)
  );
  LUT6 #(
    .INIT(64'h0000007f00000000)
  ) __5293__ (
    .I5(__1912__),
    .I4(__847__),
    .I3(__1910__),
    .I2(__1909__),
    .I1(__1090__),
    .I0(__208__),
    .O(__1913__)
  );
  LUT3 #(
    .INIT(8'h07)
  ) __5294__ (
    .I2(__1913__),
    .I1(__1908__),
    .I0(__1906__),
    .O(__1914__)
  );
  LUT6 #(
    .INIT(64'hfffff11100000000)
  ) __5295__ (
    .I5(__1896__),
    .I4(__1914__),
    .I3(__1226__),
    .I2(__1904__),
    .I1(__1903__),
    .I0(__1900__),
    .O(__1915__)
  );
  LUT5 #(
    .INIT(32'hcf30aaaa)
  ) __5296__ (
    .I4(g35),
    .I3(__1915__),
    .I2(__1210__),
    .I1(__1897__),
    .I0(__449__),
    .O(__1916__)
  );
  LUT6 #(
    .INIT(64'hc3aaaaaaf0f0f0f0)
  ) __5297__ (
    .I5(g35),
    .I4(__1896__),
    .I3(__1904__),
    .I2(__765__),
    .I1(__1232__),
    .I0(__368__),
    .O(__1917__)
  );
  LUT4 #(
    .INIT(16'h0008)
  ) __5298__ (
    .I3(__1107__),
    .I2(__118__),
    .I1(__50__),
    .I0(__1359__),
    .O(__1918__)
  );
  LUT3 #(
    .INIT(8'h04)
  ) __5299__ (
    .I2(__50__),
    .I1(__118__),
    .I0(__1107__),
    .O(__1919__)
  );
  LUT5 #(
    .INIT(32'h0777ffff)
  ) __5300__ (
    .I4(__1919__),
    .I3(__1357__),
    .I2(g127),
    .I1(__1355__),
    .I0(g92),
    .O(__1920__)
  );
  LUT5 #(
    .INIT(32'h00008000)
  ) __5301__ (
    .I4(__1107__),
    .I3(__50__),
    .I2(__118__),
    .I1(__1353__),
    .I0(__904__),
    .O(__1921__)
  );
  LUT5 #(
    .INIT(32'h00000080)
  ) __5302__ (
    .I4(__1107__),
    .I3(__118__),
    .I2(__50__),
    .I1(__1357__),
    .I0(__806__),
    .O(__1922__)
  );
  LUT5 #(
    .INIT(32'h00000080)
  ) __5303__ (
    .I4(__1107__),
    .I3(__118__),
    .I2(__50__),
    .I1(__1353__),
    .I0(__209__),
    .O(__1923__)
  );
  LUT6 #(
    .INIT(64'h0000000000000070)
  ) __5304__ (
    .I5(__1923__),
    .I4(__1922__),
    .I3(__1921__),
    .I2(__1920__),
    .I1(__1918__),
    .I0(__1260__),
    .O(__1924__)
  );
  LUT6 #(
    .INIT(64'h0000000000000004)
  ) __5305__ (
    .I5(__96__),
    .I4(__1100__),
    .I3(__876__),
    .I2(__720__),
    .I1(__1367__),
    .I0(__825__),
    .O(__1925__)
  );
  LUT3 #(
    .INIT(8'hd0)
  ) __5306__ (
    .I2(__1362__),
    .I1(__886__),
    .I0(g35),
    .O(__1926__)
  );
  LUT6 #(
    .INIT(64'h000d000000000000)
  ) __5307__ (
    .I5(__1364__),
    .I4(__1107__),
    .I3(__50__),
    .I2(__118__),
    .I1(__744__),
    .I0(g35),
    .O(__1927__)
  );
  LUT5 #(
    .INIT(32'h35003f0f)
  ) __5308__ (
    .I4(__1357__),
    .I3(g35),
    .I2(__1355__),
    .I1(__587__),
    .I0(__525__),
    .O(__1928__)
  );
  LUT6 #(
    .INIT(64'hf0f0f080f0f0f0f0)
  ) __5309__ (
    .I5(__1928__),
    .I4(__1927__),
    .I3(__1926__),
    .I2(__1371__),
    .I1(__1925__),
    .I0(__221__),
    .O(__1929__)
  );
  LUT5 #(
    .INIT(32'h00008000)
  ) __5310__ (
    .I4(__118__),
    .I3(__50__),
    .I2(__1107__),
    .I1(__1370__),
    .I0(__1362__),
    .O(__1930__)
  );
  LUT6 #(
    .INIT(64'h0000000080000000)
  ) __5311__ (
    .I5(__118__),
    .I4(__493__),
    .I3(__1364__),
    .I2(__50__),
    .I1(__1107__),
    .I0(__1370__),
    .O(__1931__)
  );
  LUT6 #(
    .INIT(64'h0000000080000000)
  ) __5312__ (
    .I5(__118__),
    .I4(__50__),
    .I3(__1107__),
    .I2(__1370__),
    .I1(__1357__),
    .I0(__789__),
    .O(__1932__)
  );
  LUT6 #(
    .INIT(64'h0000000000000777)
  ) __5313__ (
    .I5(__1932__),
    .I4(__1931__),
    .I3(__620__),
    .I2(__1374__),
    .I1(__1143__),
    .I0(__1930__),
    .O(__1933__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5314__ (
    .I5(__1379__),
    .I4(__638__),
    .I3(__1378__),
    .I2(__626__),
    .I1(__1373__),
    .I0(__432__),
    .O(__1934__)
  );
  LUT5 #(
    .INIT(32'hf4ffffff)
  ) __5315__ (
    .I4(__1934__),
    .I3(__1933__),
    .I2(__1929__),
    .I1(__1370__),
    .I0(__1924__),
    .O(__1935__)
  );
  LUT3 #(
    .INIT(8'h01)
  ) __5316__ (
    .I2(__944__),
    .I1(__296__),
    .I0(__1600__),
    .O(__1936__)
  );
  LUT5 #(
    .INIT(32'h33aaf0f0)
  ) __5317__ (
    .I4(g35),
    .I3(__1936__),
    .I2(__946__),
    .I1(__1597__),
    .I0(__987__),
    .O(__1937__)
  );
  LUT6 #(
    .INIT(64'h3fc0ff00aaaaaaaa)
  ) __5318__ (
    .I5(g35),
    .I4(__1430__),
    .I3(__491__),
    .I2(__142__),
    .I1(__243__),
    .I0(__1094__),
    .O(__1938__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5319__ (
    .I1(__659__),
    .I0(g35),
    .O(__1939__)
  );
  LUT5 #(
    .INIT(32'hccaaf0f0)
  ) __5320__ (
    .I4(g35),
    .I3(__1009__),
    .I2(__804__),
    .I1(__214__),
    .I0(__42__),
    .O(__1940__)
  );
  LUT6 #(
    .INIT(64'h1a303030ff00ff00)
  ) __5321__ (
    .I5(g35),
    .I4(__252__),
    .I3(__790__),
    .I2(__642__),
    .I1(__1817__),
    .I0(__1818__),
    .O(__1941__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __5322__ (
    .I2(__1211__),
    .I1(__471__),
    .I0(__741__),
    .O(__1942__)
  );
  LUT5 #(
    .INIT(32'h00000008)
  ) __5323__ (
    .I4(__69__),
    .I3(__1077__),
    .I2(__721__),
    .I1(__288__),
    .I0(__788__),
    .O(__1943__)
  );
  LUT6 #(
    .INIT(64'hebaa00aa00000000)
  ) __5324__ (
    .I5(g35),
    .I4(__1943__),
    .I3(__1678__),
    .I2(__46__),
    .I1(__1942__),
    .I0(__1084__),
    .O(__1944__)
  );
  LUT5 #(
    .INIT(32'h0000b400)
  ) __5325__ (
    .I4(__544__),
    .I3(g35),
    .I2(__776__),
    .I1(__1147__),
    .I0(__1700__),
    .O(__1945__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5326__ (
    .I1(__689__),
    .I0(__253__),
    .O(__1946__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5327__ (
    .I5(g35),
    .I4(__1946__),
    .I3(__1727__),
    .I2(__853__),
    .I1(__628__),
    .I0(__1391__),
    .O(__1947__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5328__ (
    .I1(__645__),
    .I0(__1014__),
    .O(__1948__)
  );
  LUT4 #(
    .INIT(16'h0004)
  ) __5329__ (
    .I3(__779__),
    .I2(__845__),
    .I1(__1414__),
    .I0(__639__),
    .O(__1949__)
  );
  LUT6 #(
    .INIT(64'h990f0f0f0f0f0f0f)
  ) __5330__ (
    .I5(__1503__),
    .I4(__1471__),
    .I3(__1949__),
    .I2(__980__),
    .I1(__1060__),
    .I0(__1948__),
    .O(__1950__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __5331__ (
    .I2(g35),
    .I1(__1950__),
    .I0(__950__),
    .O(__1951__)
  );
  LUT5 #(
    .INIT(32'hefefff00)
  ) __5332__ (
    .I4(g35),
    .I3(__722__),
    .I2(__1841__),
    .I1(__467__),
    .I0(__1843__),
    .O(__1952__)
  );
  LUT6 #(
    .INIT(64'h0000000000009009)
  ) __5333__ (
    .I5(__917__),
    .I4(__353__),
    .I3(g72),
    .I2(__591__),
    .I1(g73),
    .I0(__851__),
    .O(__1953__)
  );
  LUT6 #(
    .INIT(64'h3f3f002affff00aa)
  ) __5334__ (
    .I5(__972__),
    .I4(__1237__),
    .I3(__653__),
    .I2(__1444__),
    .I1(__1953__),
    .I0(__934__),
    .O(__1954__)
  );
  LUT5 #(
    .INIT(32'h33aaf0f0)
  ) __5335__ (
    .I4(g35),
    .I3(__1708__),
    .I2(__732__),
    .I1(__1954__),
    .I0(__653__),
    .O(__1955__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5336__ (
    .I1(__191__),
    .I0(__958__),
    .O(__1956__)
  );
  LUT6 #(
    .INIT(64'hc3aaaaaaf0f0f0f0)
  ) __5337__ (
    .I5(g35),
    .I4(__1643__),
    .I3(__1956__),
    .I2(__1104__),
    .I1(__578__),
    .I0(__1274__),
    .O(__1957__)
  );
  LUT3 #(
    .INIT(8'h01)
  ) __5338__ (
    .I2(__595__),
    .I1(__112__),
    .I0(__1521__),
    .O(__1958__)
  );
  LUT5 #(
    .INIT(32'hc3aaf0f0)
  ) __5339__ (
    .I4(g35),
    .I3(__1958__),
    .I2(__17__),
    .I1(__491__),
    .I0(__1058__),
    .O(__1959__)
  );
  LUT6 #(
    .INIT(64'h5ffffffffffffff3)
  ) __5340__ (
    .I5(__1205__),
    .I4(__838__),
    .I3(__1070__),
    .I2(__392__),
    .I1(__492__),
    .I0(__959__),
    .O(__1960__)
  );
  LUT6 #(
    .INIT(64'h000a5555cccccccc)
  ) __5341__ (
    .I5(g35),
    .I4(__143__),
    .I3(__1681__),
    .I2(__1680__),
    .I1(__392__),
    .I0(__1960__),
    .O(__1961__)
  );
  LUT3 #(
    .INIT(8'hb4)
  ) __5342__ (
    .I2(__891__),
    .I1(g35),
    .I0(__315__),
    .O(__1962__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5343__ (
    .I1(g35),
    .I0(g64),
    .O(__1963__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5344__ (
    .I1(__313__),
    .I0(__569__),
    .O(__1964__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5345__ (
    .I1(__418__),
    .I0(__1173__),
    .O(__1965__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5346__ (
    .I5(g35),
    .I4(__1965__),
    .I3(__1964__),
    .I2(__109__),
    .I1(__986__),
    .I0(__1391__),
    .O(__1966__)
  );
  LUT5 #(
    .INIT(32'h575d0a00)
  ) __5347__ (
    .I4(__1264__),
    .I3(__874__),
    .I2(__1295__),
    .I1(__457__),
    .I0(g35),
    .O(__1967__)
  );
  LUT6 #(
    .INIT(64'h000000000000bf00)
  ) __5348__ (
    .I5(__989__),
    .I4(__418__),
    .I3(g35),
    .I2(__1303__),
    .I1(__1670__),
    .I0(__810__),
    .O(__1968__)
  );
  LUT2 #(
    .INIT(4'h2)
  ) __5349__ (
    .I1(__962__),
    .I0(__1034__),
    .O(__1969__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5350__ (
    .I5(g35),
    .I4(__1969__),
    .I3(__1393__),
    .I2(__929__),
    .I1(__634__),
    .I0(__1391__),
    .O(__1970__)
  );
  LUT6 #(
    .INIT(64'hc3aaaaaaf0f0f0f0)
  ) __5351__ (
    .I5(g35),
    .I4(__1311__),
    .I3(__1319__),
    .I2(__622__),
    .I1(__1223__),
    .I0(__846__),
    .O(__1971__)
  );
  LUT6 #(
    .INIT(64'hfffc0003aaaaaaaa)
  ) __5352__ (
    .I5(g35),
    .I4(__1134__),
    .I3(__1269__),
    .I2(__1638__),
    .I1(__318__),
    .I0(__483__),
    .O(__1972__)
  );
  LUT6 #(
    .INIT(64'h00000000bf000000)
  ) __5353__ (
    .I5(__660__),
    .I4(__881__),
    .I3(__170__),
    .I2(__204__),
    .I1(__299__),
    .I0(__717__),
    .O(__1973__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5354__ (
    .I1(__134__),
    .I0(__1973__),
    .O(__1974__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5355__ (
    .I1(__170__),
    .I0(__1401__),
    .O(__1975__)
  );
  LUT6 #(
    .INIT(64'h7777f0f0ff00ff00)
  ) __5356__ (
    .I5(g35),
    .I4(__1115__),
    .I3(__717__),
    .I2(__1975__),
    .I1(__148__),
    .I0(__1974__),
    .O(__1976__)
  );
  LUT5 #(
    .INIT(32'h0000b400)
  ) __5357__ (
    .I4(__631__),
    .I3(g35),
    .I2(__896__),
    .I1(__214__),
    .I0(__1730__),
    .O(__1977__)
  );
  LUT6 #(
    .INIT(64'hffffff22f0f0f0f0)
  ) __5358__ (
    .I5(g35),
    .I4(__100__),
    .I3(__1512__),
    .I2(__862__),
    .I1(__84__),
    .I0(__913__),
    .O(__1978__)
  );
  LUT6 #(
    .INIT(64'h0000f3ff00005155)
  ) __5359__ (
    .I5(__441__),
    .I4(__1485__),
    .I3(__1143__),
    .I2(__1186__),
    .I1(__961__),
    .I0(__245__),
    .O(__1979__)
  );
  LUT6 #(
    .INIT(64'h0a0a5f0a0a0a1b0a)
  ) __5360__ (
    .I5(__441__),
    .I4(__1485__),
    .I3(__1248__),
    .I2(__768__),
    .I1(__245__),
    .I0(__1979__),
    .O(__1980__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __5361__ (
    .I1(__196__),
    .I0(__1489__),
    .O(__1981__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5362__ (
    .I5(g35),
    .I4(__190__),
    .I3(__1981__),
    .I2(__64__),
    .I1(__431__),
    .I0(__1980__),
    .O(__1982__)
  );
  LUT6 #(
    .INIT(64'h0000000000000080)
  ) __5363__ (
    .I5(g113),
    .I4(__1283__),
    .I3(__639__),
    .I2(__1060__),
    .I1(__779__),
    .I0(__1522__),
    .O(__1983__)
  );
  LUT5 #(
    .INIT(32'haaf030f0)
  ) __5364__ (
    .I4(__1348__),
    .I3(g35),
    .I2(__179__),
    .I1(__1983__),
    .I0(__728__),
    .O(__1984__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5365__ (
    .I1(g35),
    .I0(g113),
    .O(__1985__)
  );
  LUT5 #(
    .INIT(32'hffa0cfc0)
  ) __5366__ (
    .I4(__1452__),
    .I3(__1228__),
    .I2(g35),
    .I1(__941__),
    .I0(__579__),
    .O(__1986__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __5367__ (
    .I2(g35),
    .I1(__1688__),
    .I0(__1271__),
    .O(__1987__)
  );
  LUT6 #(
    .INIT(64'hdfdfdfdfdfffffff)
  ) __5368__ (
    .I5(g134),
    .I4(__884__),
    .I3(g99),
    .I2(__1005__),
    .I1(__1292__),
    .I0(__230__),
    .O(__1988__)
  );
  LUT5 #(
    .INIT(32'h73bbc000)
  ) __5369__ (
    .I4(__777__),
    .I3(__197__),
    .I2(__214__),
    .I1(g35),
    .I0(__1665__),
    .O(__1989__)
  );
  LUT6 #(
    .INIT(64'h3fffc000aaaaaaaa)
  ) __5370__ (
    .I5(g35),
    .I4(__1230__),
    .I3(__13__),
    .I2(__711__),
    .I1(__1718__),
    .I0(__470__),
    .O(__1990__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5371__ (
    .I1(g35),
    .I0(__707__),
    .O(__1991__)
  );
  LUT6 #(
    .INIT(64'h7fd55555aa000000)
  ) __5372__ (
    .I5(__972__),
    .I4(__650__),
    .I3(__917__),
    .I2(__1227__),
    .I1(__1462__),
    .I0(g35),
    .O(__1992__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5373__ (
    .I1(__296__),
    .I0(__1600__),
    .O(__1993__)
  );
  LUT6 #(
    .INIT(64'hf055f0f0cccccccc)
  ) __5374__ (
    .I5(g35),
    .I4(__1993__),
    .I3(__1027__),
    .I2(__1109__),
    .I1(__987__),
    .I0(__1597__),
    .O(__1994__)
  );
  LUT5 #(
    .INIT(32'h00009009)
  ) __5375__ (
    .I4(__353__),
    .I3(g72),
    .I2(__591__),
    .I1(g73),
    .I0(__851__),
    .O(__1995__)
  );
  LUT6 #(
    .INIT(64'h0000000000000008)
  ) __5376__ (
    .I5(__917__),
    .I4(__972__),
    .I3(g113),
    .I2(__1283__),
    .I1(__1995__),
    .I0(__1643__),
    .O(__1996__)
  );
  LUT6 #(
    .INIT(64'hf30caaaaf0f0f0f0)
  ) __5377__ (
    .I5(g35),
    .I4(__1996__),
    .I3(__749__),
    .I2(__1208__),
    .I1(__191__),
    .I0(__141__),
    .O(__1997__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5378__ (
    .I5(g35),
    .I4(__1145__),
    .I3(__1969__),
    .I2(__1054__),
    .I1(__89__),
    .I0(__1391__),
    .O(__1998__)
  );
  LUT6 #(
    .INIT(64'hffff44f400f000f0)
  ) __5379__ (
    .I5(__1389__),
    .I4(__1101__),
    .I3(g35),
    .I2(__933__),
    .I1(__1388__),
    .I0(__732__),
    .O(__1999__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5380__ (
    .I1(__705__),
    .I0(__509__),
    .O(__2000__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5381__ (
    .I5(g35),
    .I4(__2000__),
    .I3(__1823__),
    .I2(__119__),
    .I1(__458__),
    .I0(__1391__),
    .O(__2001__)
  );
  LUT6 #(
    .INIT(64'hff75aa20ff00ff00)
  ) __5382__ (
    .I5(g35),
    .I4(__779__),
    .I3(__53__),
    .I2(__599__),
    .I1(__461__),
    .I0(__1586__),
    .O(__2002__)
  );
  LUT5 #(
    .INIT(32'hfefeff00)
  ) __5383__ (
    .I4(g35),
    .I3(__388__),
    .I2(__44__),
    .I1(__200__),
    .I0(__610__),
    .O(__2003__)
  );
  LUT6 #(
    .INIT(64'h3fffc000aaaaaaaa)
  ) __5384__ (
    .I5(g35),
    .I4(__235__),
    .I3(__962__),
    .I2(__1145__),
    .I1(__1034__),
    .I0(__298__),
    .O(__2004__)
  );
  LUT4 #(
    .INIT(16'h8000)
  ) __5385__ (
    .I3(__519__),
    .I2(__1224__),
    .I1(__1190__),
    .I0(__614__),
    .O(__2005__)
  );
  LUT4 #(
    .INIT(16'h8000)
  ) __5386__ (
    .I3(__757__),
    .I2(__810__),
    .I1(__445__),
    .I0(__2005__),
    .O(__2006__)
  );
  LUT5 #(
    .INIT(32'h78ccffcc)
  ) __5387__ (
    .I4(__752__),
    .I3(g35),
    .I2(__629__),
    .I1(__605__),
    .I0(__2006__),
    .O(__2007__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __5388__ (
    .I2(g35),
    .I1(__778__),
    .I0(__954__),
    .O(__2008__)
  );
  LUT6 #(
    .INIT(64'hccccccacaaaaaaaa)
  ) __5389__ (
    .I5(g35),
    .I4(__507__),
    .I3(__1032__),
    .I2(__709__),
    .I1(__88__),
    .I0(__835__),
    .O(__2009__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5390__ (
    .I5(g35),
    .I4(__1837__),
    .I3(__1715__),
    .I2(__703__),
    .I1(__1049__),
    .I0(__1391__),
    .O(__2010__)
  );
  LUT5 #(
    .INIT(32'hacaacccc)
  ) __5391__ (
    .I4(g35),
    .I3(__1531__),
    .I2(__1476__),
    .I1(__939__),
    .I0(__560__),
    .O(__2011__)
  );
  LUT4 #(
    .INIT(16'h8000)
  ) __5392__ (
    .I3(__935__),
    .I2(__451__),
    .I1(__1162__),
    .I0(__302__),
    .O(__2012__)
  );
  LUT4 #(
    .INIT(16'h3caa)
  ) __5393__ (
    .I3(g35),
    .I2(__840__),
    .I1(__2012__),
    .I0(__1172__),
    .O(__2013__)
  );
  LUT6 #(
    .INIT(64'h00001cccf0f0f0f0)
  ) __5394__ (
    .I5(g35),
    .I4(__1441__),
    .I3(__1876__),
    .I2(__288__),
    .I1(__721__),
    .I0(__788__),
    .O(__2014__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5395__ (
    .I1(g35),
    .I0(__1039__),
    .O(__2015__)
  );
  LUT6 #(
    .INIT(64'hff00ccccf0f0aaaa)
  ) __5396__ (
    .I5(__69__),
    .I4(__1077__),
    .I3(__780__),
    .I2(__222__),
    .I1(__727__),
    .I0(__39__),
    .O(__2016__)
  );
  LUT6 #(
    .INIT(64'hdfdfdfdfdfffffff)
  ) __5397__ (
    .I5(g134),
    .I4(__884__),
    .I3(g99),
    .I2(__287__),
    .I1(__2016__),
    .I0(__990__),
    .O(__2017__)
  );
  LUT6 #(
    .INIT(64'haaaaaaaccccccccc)
  ) __5398__ (
    .I5(g35),
    .I4(__728__),
    .I3(__1348__),
    .I2(__801__),
    .I1(__673__),
    .I0(__1001__),
    .O(__2018__)
  );
  LUT6 #(
    .INIT(64'h2000000000000000)
  ) __5399__ (
    .I5(__465__),
    .I4(__1227__),
    .I3(__917__),
    .I2(__353__),
    .I1(__842__),
    .I0(__972__),
    .O(__2019__)
  );
  LUT5 #(
    .INIT(32'hccaa0f0f)
  ) __5400__ (
    .I4(__2019__),
    .I3(__1503__),
    .I2(__503__),
    .I1(__1098__),
    .I0(__611__),
    .O(__2020__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __5401__ (
    .I2(g35),
    .I1(__2020__),
    .I0(__864__),
    .O(__2021__)
  );
  LUT3 #(
    .INIT(8'h78)
  ) __5402__ (
    .I2(__385__),
    .I1(g35),
    .I0(__1233__),
    .O(__2022__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5403__ (
    .I1(__196__),
    .I0(__1489__),
    .O(__2023__)
  );
  LUT6 #(
    .INIT(64'hf055f0f0cccccccc)
  ) __5404__ (
    .I5(g35),
    .I4(__2023__),
    .I3(__190__),
    .I2(__411__),
    .I1(__64__),
    .I0(__1980__),
    .O(__2024__)
  );
  LUT6 #(
    .INIT(64'h557f55d500aa0000)
  ) __5405__ (
    .I5(__633__),
    .I4(__126__),
    .I3(__1817__),
    .I2(__587__),
    .I1(__1816__),
    .I0(g35),
    .O(__2025__)
  );
  LUT2 #(
    .INIT(4'h2)
  ) __5406__ (
    .I1(__561__),
    .I0(__863__),
    .O(__2026__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5407__ (
    .I1(__425__),
    .I0(__267__),
    .O(__2027__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5408__ (
    .I5(g35),
    .I4(__2027__),
    .I3(__2026__),
    .I2(__953__),
    .I1(__1161__),
    .I0(__1391__),
    .O(__2028__)
  );
  LUT3 #(
    .INIT(8'h2c)
  ) __5409__ (
    .I2(__299__),
    .I1(__631__),
    .I0(__736__),
    .O(__2029__)
  );
  LUT5 #(
    .INIT(32'h0af0cccc)
  ) __5410__ (
    .I4(g35),
    .I3(__2029__),
    .I2(__319__),
    .I1(__713__),
    .I0(__437__),
    .O(__2030__)
  );
  LUT5 #(
    .INIT(32'h00ccf0aa)
  ) __5411__ (
    .I4(g72),
    .I3(g73),
    .I2(__439__),
    .I1(__501__),
    .I0(__34__),
    .O(__2031__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __5412__ (
    .I2(g35),
    .I1(__2031__),
    .I0(__73__),
    .O(__2032__)
  );
  LUT6 #(
    .INIT(64'h0000f3ff00005155)
  ) __5413__ (
    .I5(__441__),
    .I4(__1485__),
    .I3(__1186__),
    .I2(__1143__),
    .I1(__961__),
    .I0(__583__),
    .O(__2033__)
  );
  LUT6 #(
    .INIT(64'h88d8888888d888d8)
  ) __5414__ (
    .I5(__583__),
    .I4(__441__),
    .I3(__1485__),
    .I2(__1248__),
    .I1(__768__),
    .I0(__2033__),
    .O(__2034__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5415__ (
    .I1(__860__),
    .I0(__1782__),
    .O(__2035__)
  );
  LUT6 #(
    .INIT(64'hf055f0f0cccccccc)
  ) __5416__ (
    .I5(g35),
    .I4(__2035__),
    .I3(__908__),
    .I2(__336__),
    .I1(__7__),
    .I0(__2034__),
    .O(__2036__)
  );
  LUT6 #(
    .INIT(64'h0000333fccfcffaa)
  ) __5417__ (
    .I5(__384__),
    .I4(__448__),
    .I3(__1195__),
    .I2(__550__),
    .I1(__1142__),
    .I0(__1033__),
    .O(__2037__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __5418__ (
    .I2(g35),
    .I1(__2037__),
    .I0(__1033__),
    .O(__2038__)
  );
  LUT4 #(
    .INIT(16'h7580)
  ) __5419__ (
    .I3(__546__),
    .I2(__214__),
    .I1(__606__),
    .I0(g35),
    .O(__2039__)
  );
  LUT4 #(
    .INIT(16'h8000)
  ) __5420__ (
    .I3(__442__),
    .I2(__502__),
    .I1(__45__),
    .I0(__160__),
    .O(__2040__)
  );
  LUT4 #(
    .INIT(16'h1f30)
  ) __5421__ (
    .I3(__897__),
    .I2(g35),
    .I1(__18__),
    .I0(__2040__),
    .O(__2041__)
  );
  LUT6 #(
    .INIT(64'h6c206c6cf0f0f0f0)
  ) __5422__ (
    .I5(g35),
    .I4(__973__),
    .I3(__279__),
    .I2(__1078__),
    .I1(__251__),
    .I0(__1819__),
    .O(__2042__)
  );
  LUT6 #(
    .INIT(64'h0000007f00000000)
  ) __5423__ (
    .I5(g35),
    .I4(__412__),
    .I3(__566__),
    .I2(__1303__),
    .I1(__810__),
    .I0(__1302__),
    .O(__2043__)
  );
  LUT6 #(
    .INIT(64'h0000000500000080)
  ) __5424__ (
    .I5(__631__),
    .I4(__35__),
    .I3(__437__),
    .I2(__299__),
    .I1(__736__),
    .I0(__90__),
    .O(__2044__)
  );
  LUT6 #(
    .INIT(64'hfcff0300aaaaaaaa)
  ) __5425__ (
    .I5(g35),
    .I4(__2044__),
    .I3(__1730__),
    .I2(__580__),
    .I1(__1177__),
    .I0(__299__),
    .O(__2045__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5426__ (
    .I1(__313__),
    .I0(__569__),
    .O(__2046__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5427__ (
    .I5(g35),
    .I4(__989__),
    .I3(__2046__),
    .I2(__937__),
    .I1(__1262__),
    .I0(__1391__),
    .O(__2047__)
  );
  LUT6 #(
    .INIT(64'h48888888ffff0000)
  ) __5428__ (
    .I5(g35),
    .I4(__926__),
    .I3(__151__),
    .I2(__1192__),
    .I1(__1517__),
    .I0(__241__),
    .O(__2048__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5429__ (
    .I5(g35),
    .I4(__2046__),
    .I3(__1794__),
    .I2(__1191__),
    .I1(__147__),
    .I0(__1391__),
    .O(__2049__)
  );
  LUT4 #(
    .INIT(16'h7580)
  ) __5430__ (
    .I3(__342__),
    .I2(__1147__),
    .I1(__914__),
    .I0(g35),
    .O(__2050__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __5431__ (
    .I2(__313__),
    .I1(__569__),
    .I0(__989__),
    .O(__2051__)
  );
  LUT4 #(
    .INIT(16'h9009)
  ) __5432__ (
    .I3(g72),
    .I2(__629__),
    .I1(g73),
    .I0(__664__),
    .O(__2052__)
  );
  LUT6 #(
    .INIT(64'h5ffffff3ffffffff)
  ) __5433__ (
    .I5(__2052__),
    .I4(__757__),
    .I3(__605__),
    .I2(__810__),
    .I1(__2051__),
    .I0(__1525__),
    .O(__2053__)
  );
  LUT5 #(
    .INIT(32'h82000082)
  ) __5434__ (
    .I4(g72),
    .I3(__629__),
    .I2(g73),
    .I1(__664__),
    .I0(__605__),
    .O(__2054__)
  );
  LUT6 #(
    .INIT(64'hf030f050f0f0f0f0)
  ) __5435__ (
    .I5(__2054__),
    .I4(__757__),
    .I3(__810__),
    .I2(__2053__),
    .I1(__1493__),
    .I0(__1506__),
    .O(__2055__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __5436__ (
    .I2(__412__),
    .I1(__900__),
    .I0(__817__),
    .O(__2056__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __5437__ (
    .I2(__253__),
    .I1(__689__),
    .I0(__623__),
    .O(__2057__)
  );
  LUT6 #(
    .INIT(64'hffffffff135fffff)
  ) __5438__ (
    .I5(__757__),
    .I4(__810__),
    .I3(__1385__),
    .I2(__2054__),
    .I1(__2057__),
    .I0(__2056__),
    .O(__2058__)
  );
  LUT6 #(
    .INIT(64'hc0a0ffffffffffff)
  ) __5439__ (
    .I5(__2058__),
    .I4(__2055__),
    .I3(__810__),
    .I2(__1773__),
    .I1(__1584__),
    .I0(__1528__),
    .O(__2059__)
  );
  LUT6 #(
    .INIT(64'hff07ffffffffffff)
  ) __5440__ (
    .I5(g113),
    .I4(__2052__),
    .I3(__2059__),
    .I2(g134),
    .I1(__884__),
    .I0(g99),
    .O(__2060__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5441__ (
    .I1(__566__),
    .I0(__548__),
    .O(__2061__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5442__ (
    .I5(g35),
    .I4(__2061__),
    .I3(__1805__),
    .I2(__1151__),
    .I1(__568__),
    .I0(__1391__),
    .O(__2062__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __5443__ (
    .I2(g35),
    .I1(__789__),
    .I0(__1204__),
    .O(__2063__)
  );
  LUT6 #(
    .INIT(64'haaaaaaaccccccccc)
  ) __5444__ (
    .I5(g35),
    .I4(__944__),
    .I3(__296__),
    .I2(__1600__),
    .I1(__454__),
    .I0(__139__),
    .O(__2064__)
  );
  LUT5 #(
    .INIT(32'h80000000)
  ) __5445__ (
    .I4(__606__),
    .I3(__214__),
    .I2(__719__),
    .I1(__546__),
    .I0(__1117__),
    .O(__2065__)
  );
  LUT5 #(
    .INIT(32'h73bbc000)
  ) __5446__ (
    .I4(__285__),
    .I3(__777__),
    .I2(__214__),
    .I1(g35),
    .I0(__2065__),
    .O(__2066__)
  );
  LUT3 #(
    .INIT(8'h08)
  ) __5447__ (
    .I2(__118__),
    .I1(__50__),
    .I0(__1107__),
    .O(__2067__)
  );
  LUT3 #(
    .INIT(8'h04)
  ) __5448__ (
    .I2(__1107__),
    .I1(__50__),
    .I0(__118__),
    .O(__2068__)
  );
  LUT6 #(
    .INIT(64'h050f153f0f0fffff)
  ) __5449__ (
    .I5(__2068__),
    .I4(__2067__),
    .I3(__1353__),
    .I2(__1359__),
    .I1(__1153__),
    .I0(__44__),
    .O(__2069__)
  );
  LUT6 #(
    .INIT(64'h553355ff550f55ff)
  ) __5450__ (
    .I5(__50__),
    .I4(__1357__),
    .I3(__1364__),
    .I2(__796__),
    .I1(__722__),
    .I0(__1220__),
    .O(__2070__)
  );
  LUT5 #(
    .INIT(32'hfff3ff1f)
  ) __5451__ (
    .I4(__50__),
    .I3(__1107__),
    .I2(__118__),
    .I1(__1357__),
    .I0(__1355__),
    .O(__2071__)
  );
  LUT5 #(
    .INIT(32'h0f8f8f8f)
  ) __5452__ (
    .I4(__1364__),
    .I3(__2068__),
    .I2(__1370__),
    .I1(__2071__),
    .I0(__0__),
    .O(__2072__)
  );
  LUT3 #(
    .INIT(8'hd0)
  ) __5453__ (
    .I2(__1362__),
    .I1(__207__),
    .I0(g35),
    .O(__2073__)
  );
  LUT6 #(
    .INIT(64'h000d000000000000)
  ) __5454__ (
    .I5(__1364__),
    .I4(__1107__),
    .I3(__50__),
    .I2(__118__),
    .I1(__716__),
    .I0(g35),
    .O(__2074__)
  );
  LUT5 #(
    .INIT(32'h35003f0f)
  ) __5455__ (
    .I4(__1357__),
    .I3(g35),
    .I2(__1355__),
    .I1(__175__),
    .I0(__693__),
    .O(__2075__)
  );
  LUT6 #(
    .INIT(64'hf0f0f080f0f0f0f0)
  ) __5456__ (
    .I5(__2075__),
    .I4(__2074__),
    .I3(__2073__),
    .I2(__1371__),
    .I1(__1925__),
    .I0(__563__),
    .O(__2076__)
  );
  LUT6 #(
    .INIT(64'h0000000080000000)
  ) __5457__ (
    .I5(__50__),
    .I4(__1107__),
    .I3(__118__),
    .I2(__1370__),
    .I1(__1357__),
    .I0(__232__),
    .O(__2077__)
  );
  LUT6 #(
    .INIT(64'h000000000fff0777)
  ) __5458__ (
    .I5(__2077__),
    .I4(__1118__),
    .I3(__1380__),
    .I2(__672__),
    .I1(__500__),
    .I0(__1373__),
    .O(__2078__)
  );
  LUT3 #(
    .INIT(8'h08)
  ) __5459__ (
    .I2(__50__),
    .I1(__1107__),
    .I0(__118__),
    .O(__2079__)
  );
  LUT6 #(
    .INIT(64'h0777ffffffffffff)
  ) __5460__ (
    .I5(__1364__),
    .I4(__1370__),
    .I3(__1919__),
    .I2(__1599__),
    .I1(__2079__),
    .I0(__161__),
    .O(__2080__)
  );
  LUT5 #(
    .INIT(32'h07770000)
  ) __5461__ (
    .I4(__2080__),
    .I3(__1378__),
    .I2(__443__),
    .I1(__1930__),
    .I0(__892__),
    .O(__2081__)
  );
  LUT6 #(
    .INIT(64'hff07ffffffffffff)
  ) __5462__ (
    .I5(__2081__),
    .I4(__2078__),
    .I3(__2076__),
    .I2(__2072__),
    .I1(__2070__),
    .I0(__2069__),
    .O(__2082__)
  );
  LUT4 #(
    .INIT(16'h0008)
  ) __5463__ (
    .I3(__1107__),
    .I2(__118__),
    .I1(__50__),
    .I0(__1353__),
    .O(__2083__)
  );
  LUT5 #(
    .INIT(32'h00000080)
  ) __5464__ (
    .I4(__1107__),
    .I3(__118__),
    .I2(__50__),
    .I1(__1357__),
    .I0(__1061__),
    .O(__2084__)
  );
  LUT5 #(
    .INIT(32'hc0f7f7f7)
  ) __5465__ (
    .I4(__1364__),
    .I3(__316__),
    .I2(__2068__),
    .I1(__1357__),
    .I0(__1121__),
    .O(__2085__)
  );
  LUT6 #(
    .INIT(64'h0000153f00000000)
  ) __5466__ (
    .I5(__2085__),
    .I4(__2084__),
    .I3(__1200__),
    .I2(__2083__),
    .I1(__345__),
    .I0(__1918__),
    .O(__2086__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5467__ (
    .I1(g35),
    .I0(__790__),
    .O(__2087__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5468__ (
    .I1(g35),
    .I0(__854__),
    .O(__2088__)
  );
  LUT6 #(
    .INIT(64'h0020000000300000)
  ) __5469__ (
    .I5(g35),
    .I4(__1364__),
    .I3(__50__),
    .I2(__1107__),
    .I1(__118__),
    .I0(__799__),
    .O(__2089__)
  );
  LUT6 #(
    .INIT(64'hff4f0000ff440000)
  ) __5470__ (
    .I5(__1362__),
    .I4(__1371__),
    .I3(__2089__),
    .I2(__2088__),
    .I1(__1355__),
    .I0(__2087__),
    .O(__2090__)
  );
  LUT6 #(
    .INIT(64'h0777ffffffffffff)
  ) __5471__ (
    .I5(__1364__),
    .I4(__1370__),
    .I3(__508__),
    .I2(__2079__),
    .I1(__1486__),
    .I0(__1919__),
    .O(__2091__)
  );
  LUT6 #(
    .INIT(64'h7f7f7f7fffff00ff)
  ) __5472__ (
    .I5(__1370__),
    .I4(g53),
    .I3(__205__),
    .I2(__1357__),
    .I1(__1369__),
    .I0(__1519__),
    .O(__2092__)
  );
  LUT6 #(
    .INIT(64'h0000000080000000)
  ) __5473__ (
    .I5(__50__),
    .I4(__1107__),
    .I3(__118__),
    .I2(__1370__),
    .I1(__1357__),
    .I0(__104__),
    .O(__2093__)
  );
  LUT6 #(
    .INIT(64'h0000000080000000)
  ) __5474__ (
    .I5(__118__),
    .I4(__242__),
    .I3(__1364__),
    .I2(__50__),
    .I1(__1107__),
    .I0(__1370__),
    .O(__2094__)
  );
  LUT6 #(
    .INIT(64'h0000000000007000)
  ) __5475__ (
    .I5(__2094__),
    .I4(__2093__),
    .I3(__2092__),
    .I2(__2091__),
    .I1(__1930__),
    .I0(__818__),
    .O(__2095__)
  );
  LUT4 #(
    .INIT(16'hf1ff)
  ) __5476__ (
    .I3(__2095__),
    .I2(__2090__),
    .I1(__2072__),
    .I0(__2086__),
    .O(__2096__)
  );
  LUT5 #(
    .INIT(32'h00000080)
  ) __5477__ (
    .I4(__1107__),
    .I3(__118__),
    .I2(__50__),
    .I1(__1357__),
    .I0(__429__),
    .O(__2097__)
  );
  LUT5 #(
    .INIT(32'hc8fbfbfb)
  ) __5478__ (
    .I4(__1364__),
    .I3(__363__),
    .I2(__2068__),
    .I1(__1357__),
    .I0(__1012__),
    .O(__2098__)
  );
  LUT6 #(
    .INIT(64'h0000153f00000000)
  ) __5479__ (
    .I5(__2098__),
    .I4(__2097__),
    .I3(__1159__),
    .I2(__2083__),
    .I1(__388__),
    .I0(__1918__),
    .O(__2099__)
  );
  LUT3 #(
    .INIT(8'hd0)
  ) __5480__ (
    .I2(__1362__),
    .I1(__1113__),
    .I0(g35),
    .O(__2100__)
  );
  LUT6 #(
    .INIT(64'h000d000000000000)
  ) __5481__ (
    .I5(__1364__),
    .I4(__1107__),
    .I3(__50__),
    .I2(__118__),
    .I1(__226__),
    .I0(g35),
    .O(__2101__)
  );
  LUT5 #(
    .INIT(32'h35003f0f)
  ) __5482__ (
    .I4(__1357__),
    .I3(g35),
    .I2(__1355__),
    .I1(__252__),
    .I0(__786__),
    .O(__2102__)
  );
  LUT6 #(
    .INIT(64'hf0f0f080f0f0f0f0)
  ) __5483__ (
    .I5(__2102__),
    .I4(__2101__),
    .I3(__2100__),
    .I2(__1371__),
    .I1(__1925__),
    .I0(__1127__),
    .O(__2103__)
  );
  LUT6 #(
    .INIT(64'h0000000080000000)
  ) __5484__ (
    .I5(__118__),
    .I4(__1364__),
    .I3(__50__),
    .I2(__1107__),
    .I1(__1370__),
    .I0(__219__),
    .O(__2104__)
  );
  LUT6 #(
    .INIT(64'h0000000080000000)
  ) __5485__ (
    .I5(__50__),
    .I4(__1107__),
    .I3(__118__),
    .I2(__1370__),
    .I1(__1357__),
    .I0(__415__),
    .O(__2105__)
  );
  LUT6 #(
    .INIT(64'h0000000080000000)
  ) __5486__ (
    .I5(__50__),
    .I4(__1364__),
    .I3(__1107__),
    .I2(__118__),
    .I1(__1370__),
    .I0(__1071__),
    .O(__2106__)
  );
  LUT6 #(
    .INIT(64'h7f7f7f7fffff00ff)
  ) __5487__ (
    .I5(__1370__),
    .I4(g53),
    .I3(__472__),
    .I2(__1347__),
    .I1(__1357__),
    .I0(__1369__),
    .O(__2107__)
  );
  LUT6 #(
    .INIT(64'h0000153f00000000)
  ) __5488__ (
    .I5(__2107__),
    .I4(__2106__),
    .I3(__1374__),
    .I2(__1930__),
    .I1(__310__),
    .I0(__1781__),
    .O(__2108__)
  );
  LUT6 #(
    .INIT(64'hfffffff1ffffffff)
  ) __5489__ (
    .I5(__2108__),
    .I4(__2105__),
    .I3(__2104__),
    .I2(__2103__),
    .I1(__2072__),
    .I0(__2099__),
    .O(__2109__)
  );
  LUT6 #(
    .INIT(64'h0000000000000004)
  ) __5490__ (
    .I5(__96__),
    .I4(__1100__),
    .I3(__876__),
    .I2(__720__),
    .I1(__297__),
    .I0(__825__),
    .O(__2110__)
  );
  LUT5 #(
    .INIT(32'h00000080)
  ) __5491__ (
    .I4(__1107__),
    .I3(__118__),
    .I2(__50__),
    .I1(__1357__),
    .I0(__130__),
    .O(__2111__)
  );
  LUT6 #(
    .INIT(64'h0000000000000777)
  ) __5492__ (
    .I5(__2111__),
    .I4(__2110__),
    .I3(__2083__),
    .I2(__40__),
    .I1(__1918__),
    .I0(__773__),
    .O(__2112__)
  );
  LUT3 #(
    .INIT(8'hd0)
  ) __5493__ (
    .I2(__1355__),
    .I1(__642__),
    .I0(g35),
    .O(__2113__)
  );
  LUT5 #(
    .INIT(32'h440fffff)
  ) __5494__ (
    .I4(__1364__),
    .I3(__1369__),
    .I2(__426__),
    .I1(g35),
    .I0(__123__),
    .O(__2114__)
  );
  LUT6 #(
    .INIT(64'hff00b000ff00ff00)
  ) __5495__ (
    .I5(__2114__),
    .I4(__2113__),
    .I3(__1371__),
    .I2(__1362__),
    .I1(g35),
    .I0(__981__),
    .O(__2115__)
  );
  LUT6 #(
    .INIT(64'h0000000080000000)
  ) __5496__ (
    .I5(__118__),
    .I4(__1364__),
    .I3(__50__),
    .I2(__1107__),
    .I1(__1370__),
    .I0(__590__),
    .O(__2116__)
  );
  LUT6 #(
    .INIT(64'h0000000080000000)
  ) __5497__ (
    .I5(__50__),
    .I4(__1107__),
    .I3(__118__),
    .I2(__1370__),
    .I1(__1357__),
    .I0(__494__),
    .O(__2117__)
  );
  LUT6 #(
    .INIT(64'h0000000080000000)
  ) __5498__ (
    .I5(__50__),
    .I4(__1039__),
    .I3(__1364__),
    .I2(__1107__),
    .I1(__118__),
    .I0(__1370__),
    .O(__2118__)
  );
  LUT6 #(
    .INIT(64'h7f7f7f7fffff00ff)
  ) __5499__ (
    .I5(__1370__),
    .I4(g53),
    .I3(__325__),
    .I2(__1637__),
    .I1(__1357__),
    .I0(__1369__),
    .O(__2119__)
  );
  LUT6 #(
    .INIT(64'h0000153f00000000)
  ) __5500__ (
    .I5(__2119__),
    .I4(__2118__),
    .I3(__1374__),
    .I2(__270__),
    .I1(__1930__),
    .I0(__1553__),
    .O(__2120__)
  );
  LUT6 #(
    .INIT(64'hfffffff1ffffffff)
  ) __5501__ (
    .I5(__2120__),
    .I4(__2117__),
    .I3(__2116__),
    .I2(__2115__),
    .I1(__2072__),
    .I0(__2112__),
    .O(__2121__)
  );
  LUT4 #(
    .INIT(16'h6996)
  ) __5502__ (
    .I3(__2121__),
    .I2(__2109__),
    .I1(__2096__),
    .I0(__2082__),
    .O(__2122__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5503__ (
    .I1(g54),
    .I0(g56),
    .O(__2123__)
  );
  LUT5 #(
    .INIT(32'hf4ffffff)
  ) __5504__ (
    .I4(__1381__),
    .I3(__1377__),
    .I2(__1372__),
    .I1(__1370__),
    .I0(__1361__),
    .O(__2124__)
  );
  LUT3 #(
    .INIT(8'hd0)
  ) __5505__ (
    .I2(__1362__),
    .I1(__880__),
    .I0(g35),
    .O(__2125__)
  );
  LUT6 #(
    .INIT(64'h000d000000000000)
  ) __5506__ (
    .I5(__1364__),
    .I4(__1107__),
    .I3(__50__),
    .I2(__118__),
    .I1(__407__),
    .I0(g35),
    .O(__2126__)
  );
  LUT5 #(
    .INIT(32'h35003f0f)
  ) __5507__ (
    .I4(__1357__),
    .I3(g35),
    .I2(__1355__),
    .I1(__126__),
    .I0(__251__),
    .O(__2127__)
  );
  LUT6 #(
    .INIT(64'hf0f0f080f0f0f0f0)
  ) __5508__ (
    .I5(__2127__),
    .I4(__2126__),
    .I3(__2125__),
    .I2(__1371__),
    .I1(__1925__),
    .I0(__1250__),
    .O(__2128__)
  );
  LUT6 #(
    .INIT(64'h0000000000000080)
  ) __5509__ (
    .I5(__1100__),
    .I4(__876__),
    .I3(__825__),
    .I2(__884__),
    .I1(__96__),
    .I0(__720__),
    .O(__2129__)
  );
  LUT6 #(
    .INIT(64'h5f5f5f3f5f5f5f5f)
  ) __5510__ (
    .I5(__50__),
    .I4(__1107__),
    .I3(__118__),
    .I2(__1357__),
    .I1(__467__),
    .I0(__932__),
    .O(__2130__)
  );
  LUT4 #(
    .INIT(16'h0080)
  ) __5511__ (
    .I3(__720__),
    .I2(__1100__),
    .I1(__876__),
    .I0(__825__),
    .O(__2131__)
  );
  LUT6 #(
    .INIT(64'h030f55ffffffffff)
  ) __5512__ (
    .I5(__2131__),
    .I4(__96__),
    .I3(__2068__),
    .I2(__2067__),
    .I1(__1035__),
    .I0(__264__),
    .O(__2132__)
  );
  LUT5 #(
    .INIT(32'h0fbf0000)
  ) __5513__ (
    .I4(__1370__),
    .I3(__2071__),
    .I2(__2132__),
    .I1(__2130__),
    .I0(__2129__),
    .O(__2133__)
  );
  LUT5 #(
    .INIT(32'h00008000)
  ) __5514__ (
    .I4(__50__),
    .I3(__1107__),
    .I2(__118__),
    .I1(__1370__),
    .I0(__1357__),
    .O(__2134__)
  );
  LUT6 #(
    .INIT(64'h0000000080000000)
  ) __5515__ (
    .I5(__118__),
    .I4(__50__),
    .I3(__1107__),
    .I2(__1370__),
    .I1(__1357__),
    .I0(__1273__),
    .O(__2135__)
  );
  LUT6 #(
    .INIT(64'h0000000000008000)
  ) __5516__ (
    .I5(__50__),
    .I4(__356__),
    .I3(__1364__),
    .I2(__1107__),
    .I1(__118__),
    .I0(__1370__),
    .O(__2136__)
  );
  LUT6 #(
    .INIT(64'h0000000000005f13)
  ) __5517__ (
    .I5(__2136__),
    .I4(__2135__),
    .I3(__223__),
    .I2(__1118__),
    .I1(__2134__),
    .I0(__1373__),
    .O(__2137__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5518__ (
    .I5(__441__),
    .I4(__1374__),
    .I3(__662__),
    .I2(__1379__),
    .I1(__1378__),
    .I0(__1188__),
    .O(__2138__)
  );
  LUT4 #(
    .INIT(16'hefff)
  ) __5519__ (
    .I3(__2138__),
    .I2(__2137__),
    .I1(__2133__),
    .I0(__2128__),
    .O(__2139__)
  );
  LUT5 #(
    .INIT(32'h00000080)
  ) __5520__ (
    .I4(__1107__),
    .I3(__118__),
    .I2(__50__),
    .I1(__1357__),
    .I0(__822__),
    .O(__2140__)
  );
  LUT5 #(
    .INIT(32'h0777ffff)
  ) __5521__ (
    .I4(__1919__),
    .I3(__1357__),
    .I2(__399__),
    .I1(__1355__),
    .I0(__1170__),
    .O(__2141__)
  );
  LUT6 #(
    .INIT(64'h0000153f00000000)
  ) __5522__ (
    .I5(__2141__),
    .I4(__2140__),
    .I3(__291__),
    .I2(__694__),
    .I1(__2083__),
    .I0(__1918__),
    .O(__2142__)
  );
  LUT3 #(
    .INIT(8'hd0)
  ) __5523__ (
    .I2(__1362__),
    .I1(__764__),
    .I0(g35),
    .O(__2143__)
  );
  LUT6 #(
    .INIT(64'h000d000000000000)
  ) __5524__ (
    .I5(__1364__),
    .I4(__1107__),
    .I3(__50__),
    .I2(__118__),
    .I1(__199__),
    .I0(g35),
    .O(__2144__)
  );
  LUT5 #(
    .INIT(32'h35003f0f)
  ) __5525__ (
    .I4(__1357__),
    .I3(g35),
    .I2(__1355__),
    .I1(__633__),
    .I0(__1078__),
    .O(__2145__)
  );
  LUT6 #(
    .INIT(64'hf0f0f040f0f0f0f0)
  ) __5526__ (
    .I5(__2145__),
    .I4(__2144__),
    .I3(__2143__),
    .I2(__1371__),
    .I1(__1925__),
    .I0(__340__),
    .O(__2146__)
  );
  LUT6 #(
    .INIT(64'h0000000080000000)
  ) __5527__ (
    .I5(__118__),
    .I4(__50__),
    .I3(__1107__),
    .I2(__1370__),
    .I1(__1204__),
    .I0(__1357__),
    .O(__2147__)
  );
  LUT6 #(
    .INIT(64'h0000000080000000)
  ) __5528__ (
    .I5(__118__),
    .I4(__961__),
    .I3(__50__),
    .I2(__1107__),
    .I1(__1370__),
    .I0(__1362__),
    .O(__2148__)
  );
  LUT6 #(
    .INIT(64'h000000000000f351)
  ) __5529__ (
    .I5(__2148__),
    .I4(__2147__),
    .I3(__428__),
    .I2(__224__),
    .I1(__1374__),
    .I0(__1373__),
    .O(__2149__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __5530__ (
    .I5(__895__),
    .I4(__1380__),
    .I3(__888__),
    .I2(__1379__),
    .I1(__910__),
    .I0(__1378__),
    .O(__2150__)
  );
  LUT5 #(
    .INIT(32'hf4ffffff)
  ) __5531__ (
    .I4(__2150__),
    .I3(__2149__),
    .I2(__2146__),
    .I1(__1370__),
    .I0(__2142__),
    .O(__2151__)
  );
  LUT6 #(
    .INIT(64'hb44b4bb44bb4b44b)
  ) __5532__ (
    .I5(__2151__),
    .I4(__2139__),
    .I3(__2124__),
    .I2(__1935__),
    .I1(__171__),
    .I0(__2123__),
    .O(__2152__)
  );
  LUT3 #(
    .INIT(8'h01)
  ) __5533__ (
    .I2(g56),
    .I1(g54),
    .I0(g53),
    .O(__2153__)
  );
  LUT6 #(
    .INIT(64'hcffcccccaaaaaaaa)
  ) __5534__ (
    .I5(g35),
    .I4(__2153__),
    .I3(__2152__),
    .I2(__2122__),
    .I1(__505__),
    .I0(__904__),
    .O(__2154__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5535__ (
    .I1(__758__),
    .I0(__916__),
    .O(__2155__)
  );
  LUT6 #(
    .INIT(64'h00000000bf000000)
  ) __5536__ (
    .I5(__1110__),
    .I4(__762__),
    .I3(__1251__),
    .I2(__758__),
    .I1(__1450__),
    .I0(__1249__),
    .O(__2156__)
  );
  LUT6 #(
    .INIT(64'haaff00ccf0f0f0f0)
  ) __5537__ (
    .I5(g35),
    .I4(__1249__),
    .I3(__2156__),
    .I2(__941__),
    .I1(__1586__),
    .I0(__2155__),
    .O(__2157__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5538__ (
    .I1(__636__),
    .I0(__688__),
    .O(__2158__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5539__ (
    .I5(g35),
    .I4(__1692__),
    .I3(__2158__),
    .I2(__948__),
    .I1(__533__),
    .I0(__1391__),
    .O(__2159__)
  );
  LUT3 #(
    .INIT(8'h04)
  ) __5540__ (
    .I2(__762__),
    .I1(g35),
    .I0(__547__),
    .O(__2160__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5541__ (
    .I5(g35),
    .I4(__457__),
    .I3(__1761__),
    .I2(__715__),
    .I1(__593__),
    .I0(__1391__),
    .O(__2161__)
  );
  LUT6 #(
    .INIT(64'hfffc0003aaaaaaaa)
  ) __5542__ (
    .I5(g35),
    .I4(__1062__),
    .I3(__595__),
    .I2(__112__),
    .I1(__1521__),
    .I0(__1058__),
    .O(__2162__)
  );
  LUT3 #(
    .INIT(8'h01)
  ) __5543__ (
    .I2(__267__),
    .I1(__425__),
    .I0(__157__),
    .O(__2163__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5544__ (
    .I5(g35),
    .I4(__2163__),
    .I3(__1790__),
    .I2(__735__),
    .I1(__1079__),
    .I0(__1391__),
    .O(__2164__)
  );
  LUT5 #(
    .INIT(32'h3caaf0f0)
  ) __5545__ (
    .I4(g35),
    .I3(__1312__),
    .I2(__361__),
    .I1(__754__),
    .I0(__20__),
    .O(__2165__)
  );
  LUT4 #(
    .INIT(16'heef0)
  ) __5546__ (
    .I3(g35),
    .I2(__822__),
    .I1(__806__),
    .I0(__249__),
    .O(__2166__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5547__ (
    .I1(g35),
    .I0(g125),
    .O(__2167__)
  );
  LUT6 #(
    .INIT(64'h7fffffff00000000)
  ) __5548__ (
    .I5(__1092__),
    .I4(g35),
    .I3(__395__),
    .I2(__635__),
    .I1(__1491__),
    .I0(__56__),
    .O(__2168__)
  );
  LUT6 #(
    .INIT(64'h00dfdf00ffff0000)
  ) __5549__ (
    .I5(g35),
    .I4(__418__),
    .I3(__1173__),
    .I2(__1303__),
    .I1(__810__),
    .I0(__1670__),
    .O(__2169__)
  );
  LUT6 #(
    .INIT(64'hffff44f400f000f0)
  ) __5550__ (
    .I5(__1389__),
    .I4(__81__),
    .I3(g35),
    .I2(__607__),
    .I1(__1388__),
    .I0(__581__),
    .O(__2170__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5551__ (
    .I1(g35),
    .I0(__672__),
    .O(__2171__)
  );
  LUT4 #(
    .INIT(16'he0ee)
  ) __5552__ (
    .I3(__1832__),
    .I2(__555__),
    .I1(__631__),
    .I0(__736__),
    .O(__2172__)
  );
  LUT6 #(
    .INIT(64'h8000aaaa7fffffff)
  ) __5553__ (
    .I5(__713__),
    .I4(__1832__),
    .I3(__289__),
    .I2(__413__),
    .I1(__116__),
    .I0(__2172__),
    .O(__2173__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __5554__ (
    .I2(g35),
    .I1(__2173__),
    .I0(__116__),
    .O(__2174__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __5555__ (
    .I1(__645__),
    .I0(__1473__),
    .O(__2175__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5556__ (
    .I5(g35),
    .I4(__1014__),
    .I3(__2175__),
    .I2(__63__),
    .I1(__589__),
    .I0(__1470__),
    .O(__2176__)
  );
  LUT6 #(
    .INIT(64'hee22eeeef0f0f0f0)
  ) __5557__ (
    .I5(g35),
    .I4(__1248__),
    .I3(__1245__),
    .I2(__1088__),
    .I1(__2056__),
    .I0(__740__),
    .O(__2177__)
  );
  LUT5 #(
    .INIT(32'h00008000)
  ) __5558__ (
    .I4(__721__),
    .I3(__69__),
    .I2(__1077__),
    .I1(__288__),
    .I0(__788__),
    .O(__2178__)
  );
  LUT5 #(
    .INIT(32'h000000f8)
  ) __5559__ (
    .I4(__186__),
    .I3(__1055__),
    .I2(g134),
    .I1(__884__),
    .I0(g99),
    .O(__2179__)
  );
  LUT6 #(
    .INIT(64'hccccf0aaf0f0f0f0)
  ) __5560__ (
    .I5(g35),
    .I4(__2179__),
    .I3(__2178__),
    .I2(__889__),
    .I1(__1279__),
    .I0(__39__),
    .O(__2180__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __5561__ (
    .I2(g35),
    .I1(__1200__),
    .I0(__773__),
    .O(__2181__)
  );
  LUT5 #(
    .INIT(32'h00008000)
  ) __5562__ (
    .I4(__757__),
    .I3(__2052__),
    .I2(__605__),
    .I1(__1303__),
    .I0(__810__),
    .O(__2182__)
  );
  LUT5 #(
    .INIT(32'h10ff0000)
  ) __5563__ (
    .I4(__548__),
    .I3(g35),
    .I2(__566__),
    .I1(__412__),
    .I0(__2182__),
    .O(__2183__)
  );
  LUT3 #(
    .INIT(8'h01)
  ) __5564__ (
    .I2(__688__),
    .I1(__457__),
    .I0(__636__),
    .O(__2184__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5565__ (
    .I5(g35),
    .I4(__2184__),
    .I3(__1761__),
    .I2(__827__),
    .I1(__164__),
    .I0(__1391__),
    .O(__2185__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5566__ (
    .I5(g35),
    .I4(__2061__),
    .I3(__1416__),
    .I2(__1088__),
    .I1(__849__),
    .I0(__1391__),
    .O(__2186__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __5567__ (
    .I1(__1207__),
    .I0(__936__),
    .O(__2187__)
  );
  LUT3 #(
    .INIT(8'h08)
  ) __5568__ (
    .I2(__293__),
    .I1(__1263__),
    .I0(__396__),
    .O(__2188__)
  );
  LUT6 #(
    .INIT(64'h4000ffff00000000)
  ) __5569__ (
    .I5(__2188__),
    .I4(__2187__),
    .I3(__1105__),
    .I2(__1036__),
    .I1(__1275__),
    .I0(__1812__),
    .O(__2189__)
  );
  LUT5 #(
    .INIT(32'h08880808)
  ) __5570__ (
    .I4(__507__),
    .I3(__1032__),
    .I2(__1041__),
    .I1(__364__),
    .I0(__2189__),
    .O(__2190__)
  );
  LUT6 #(
    .INIT(64'h00000000bf000000)
  ) __5571__ (
    .I5(__1032__),
    .I4(__507__),
    .I3(__364__),
    .I2(__1263__),
    .I1(__396__),
    .I0(__293__),
    .O(__2191__)
  );
  LUT5 #(
    .INIT(32'h0330aaaa)
  ) __5572__ (
    .I4(g35),
    .I3(__1067__),
    .I2(__2191__),
    .I1(__2190__),
    .I0(__1041__),
    .O(__2192__)
  );
  LUT4 #(
    .INIT(16'h070c)
  ) __5573__ (
    .I3(__69__),
    .I2(__721__),
    .I1(__1077__),
    .I0(__223__),
    .O(__2193__)
  );
  LUT6 #(
    .INIT(64'h00ff33330f0f5555)
  ) __5574__ (
    .I5(__69__),
    .I4(__1077__),
    .I3(__494__),
    .I2(__415__),
    .I1(__104__),
    .I0(__232__),
    .O(__2194__)
  );
  LUT6 #(
    .INIT(64'hcccccffc00ff5555)
  ) __5575__ (
    .I5(__788__),
    .I4(__288__),
    .I3(__2016__),
    .I2(__2194__),
    .I1(__721__),
    .I0(__2193__),
    .O(__2195__)
  );
  LUT3 #(
    .INIT(8'h01)
  ) __5576__ (
    .I2(__640__),
    .I1(__678__),
    .I0(__747__),
    .O(__2196__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5577__ (
    .I1(__640__),
    .I0(__250__),
    .O(__2197__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5578__ (
    .I1(__747__),
    .I0(__733__),
    .O(__2198__)
  );
  LUT6 #(
    .INIT(64'h0000000000005f13)
  ) __5579__ (
    .I5(__2198__),
    .I4(__2197__),
    .I3(__663__),
    .I2(__678__),
    .I1(__151__),
    .I0(__382__),
    .O(__2199__)
  );
  LUT6 #(
    .INIT(64'h0f0f4f4fff00ff00)
  ) __5580__ (
    .I5(g35),
    .I4(__151__),
    .I3(__390__),
    .I2(__2199__),
    .I1(__2196__),
    .I0(__2195__),
    .O(__2200__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __5581__ (
    .I2(g35),
    .I1(__1220__),
    .I0(__363__),
    .O(__2201__)
  );
  LUT6 #(
    .INIT(64'h04000000f4ffffff)
  ) __5582__ (
    .I5(__1116__),
    .I4(__1446__),
    .I3(__469__),
    .I2(__784__),
    .I1(__908__),
    .I0(__860__),
    .O(__2202__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __5583__ (
    .I2(g35),
    .I1(__2202__),
    .I0(__233__),
    .O(__2203__)
  );
  LUT5 #(
    .INIT(32'hf888ff00)
  ) __5584__ (
    .I4(g35),
    .I3(__427__),
    .I2(__479__),
    .I1(__1757__),
    .I0(__659__),
    .O(__2204__)
  );
  LUT6 #(
    .INIT(64'h0fff7f0070ff0000)
  ) __5585__ (
    .I5(__557__),
    .I4(__696__),
    .I3(g35),
    .I2(__1311__),
    .I1(__1338__),
    .I0(__1337__),
    .O(__2205__)
  );
  LUT6 #(
    .INIT(64'heaaa2aaaffff0000)
  ) __5586__ (
    .I5(g35),
    .I4(__931__),
    .I3(__784__),
    .I2(__462__),
    .I1(__1446__),
    .I0(__1148__),
    .O(__2206__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __5587__ (
    .I2(g35),
    .I1(g6744),
    .I0(__384__),
    .O(__2207__)
  );
  LUT6 #(
    .INIT(64'h00ff33330f0f5555)
  ) __5588__ (
    .I5(__795__),
    .I4(__718__),
    .I3(__38__),
    .I2(__503__),
    .I1(__864__),
    .I0(__1000__),
    .O(__2208__)
  );
  LUT3 #(
    .INIT(8'h01)
  ) __5589__ (
    .I2(__917__),
    .I1(__353__),
    .I0(__972__),
    .O(__2209__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __5590__ (
    .I1(__465__),
    .I0(__842__),
    .O(__2210__)
  );
  LUT6 #(
    .INIT(64'hff00ccccf0f0aaaa)
  ) __5591__ (
    .I5(__795__),
    .I4(__718__),
    .I3(__974__),
    .I2(__369__),
    .I1(__295__),
    .I0(__552__),
    .O(__2211__)
  );
  LUT6 #(
    .INIT(64'hefff200000000000)
  ) __5592__ (
    .I5(g35),
    .I4(__2211__),
    .I3(__2210__),
    .I2(__2209__),
    .I1(__1227__),
    .I0(__2208__),
    .O(__2212__)
  );
  LUT3 #(
    .INIT(8'hf4)
  ) __5593__ (
    .I2(__2212__),
    .I1(__1000__),
    .I0(g35),
    .O(__2213__)
  );
  LUT5 #(
    .INIT(32'h3cffaaaa)
  ) __5594__ (
    .I4(g35),
    .I3(__752__),
    .I2(__605__),
    .I1(__2006__),
    .I0(__757__),
    .O(__2214__)
  );
  LUT5 #(
    .INIT(32'h00000008)
  ) __5595__ (
    .I4(g113),
    .I3(__1283__),
    .I2(__779__),
    .I1(__1060__),
    .I0(__1405__),
    .O(__2215__)
  );
  LUT6 #(
    .INIT(64'hf0f04444ff00ff00)
  ) __5596__ (
    .I5(g35),
    .I4(__1473__),
    .I3(__980__),
    .I2(__1014__),
    .I1(__950__),
    .I0(__2215__),
    .O(__2216__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __5597__ (
    .I2(g35),
    .I1(__161__),
    .I0(__1071__),
    .O(__2217__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5598__ (
    .I5(g35),
    .I4(__1715__),
    .I3(__1393__),
    .I2(__1049__),
    .I1(__921__),
    .I0(__1391__),
    .O(__2218__)
  );
  LUT6 #(
    .INIT(64'h15405500cccccccc)
  ) __5599__ (
    .I5(g35),
    .I4(__185__),
    .I3(__764__),
    .I2(__1351__),
    .I1(__886__),
    .I0(__1788__),
    .O(__2219__)
  );
  LUT5 #(
    .INIT(32'h80000000)
  ) __5600__ (
    .I4(__359__),
    .I3(__1187__),
    .I2(__511__),
    .I1(__820__),
    .I0(__1673__),
    .O(__2220__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5601__ (
    .I1(__820__),
    .I0(__511__),
    .O(__2221__)
  );
  LUT6 #(
    .INIT(64'h0fffffffffff7777)
  ) __5602__ (
    .I5(__511__),
    .I4(__820__),
    .I3(__408__),
    .I2(__873__),
    .I1(__115__),
    .I0(__1129__),
    .O(__2222__)
  );
  LUT6 #(
    .INIT(64'h7f00000000007f00)
  ) __5603__ (
    .I5(__1187__),
    .I4(__612__),
    .I3(__2222__),
    .I2(__953__),
    .I1(__394__),
    .I0(__2221__),
    .O(__2223__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5604__ (
    .I1(__511__),
    .I0(__820__),
    .O(__2224__)
  );
  LUT6 #(
    .INIT(64'hffff0fffffff7777)
  ) __5605__ (
    .I5(__820__),
    .I4(__511__),
    .I3(__115__),
    .I2(__420__),
    .I1(__394__),
    .I0(__905__),
    .O(__2225__)
  );
  LUT6 #(
    .INIT(64'h00007f007f000000)
  ) __5606__ (
    .I5(__1187__),
    .I4(__612__),
    .I3(__2225__),
    .I2(__873__),
    .I1(__2224__),
    .I0(__324__),
    .O(__2226__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5607__ (
    .I1(__991__),
    .I0(__444__),
    .O(__2227__)
  );
  LUT6 #(
    .INIT(64'h007f7f7f00000000)
  ) __5608__ (
    .I5(__1187__),
    .I4(__2221__),
    .I3(__2227__),
    .I2(__1574__),
    .I1(__105__),
    .I0(__57__),
    .O(__2228__)
  );
  LUT6 #(
    .INIT(64'h000000f800000088)
  ) __5609__ (
    .I5(__29__),
    .I4(__511__),
    .I3(__820__),
    .I2(__979__),
    .I1(__681__),
    .I0(__255__),
    .O(__2229__)
  );
  LUT6 #(
    .INIT(64'h000007770000ffff)
  ) __5610__ (
    .I5(__2224__),
    .I4(__2229__),
    .I3(__95__),
    .I2(__349__),
    .I1(__612__),
    .I0(__1161__),
    .O(__2230__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __5611__ (
    .I1(__511__),
    .I0(__820__),
    .O(__2231__)
  );
  LUT6 #(
    .INIT(64'h0000f88800000000)
  ) __5612__ (
    .I5(__820__),
    .I4(__511__),
    .I3(__647__),
    .I2(__979__),
    .I1(__1079__),
    .I0(__681__),
    .O(__2232__)
  );
  LUT6 #(
    .INIT(64'h0000f88800000000)
  ) __5613__ (
    .I5(__511__),
    .I4(__820__),
    .I3(__359__),
    .I2(__176__),
    .I1(__335__),
    .I0(__105__),
    .O(__2233__)
  );
  LUT6 #(
    .INIT(64'h000007770000ffff)
  ) __5614__ (
    .I5(__1574__),
    .I4(__2233__),
    .I3(__79__),
    .I2(__349__),
    .I1(__612__),
    .I0(__735__),
    .O(__2234__)
  );
  LUT6 #(
    .INIT(64'h0000007f00000000)
  ) __5615__ (
    .I5(__2234__),
    .I4(__1187__),
    .I3(__2232__),
    .I2(__977__),
    .I1(__2231__),
    .I0(__991__),
    .O(__2235__)
  );
  LUT3 #(
    .INIT(8'h07)
  ) __5616__ (
    .I2(__2235__),
    .I1(__2230__),
    .I0(__2228__),
    .O(__2236__)
  );
  LUT6 #(
    .INIT(64'hfffff11100000000)
  ) __5617__ (
    .I5(__1673__),
    .I4(__2236__),
    .I3(__1674__),
    .I2(__899__),
    .I1(__2226__),
    .I0(__2223__),
    .O(__2237__)
  );
  LUT5 #(
    .INIT(32'hcf30aaaa)
  ) __5618__ (
    .I4(g35),
    .I3(__2237__),
    .I2(__290__),
    .I1(__2220__),
    .I0(__787__),
    .O(__2238__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __5619__ (
    .I2(g35),
    .I1(__395__),
    .I0(__1167__),
    .O(__2239__)
  );
  LUT6 #(
    .INIT(64'heaaa2aaaffff0000)
  ) __5620__ (
    .I5(g35),
    .I4(__314__),
    .I3(__962__),
    .I2(__1145__),
    .I1(__1034__),
    .I0(__951__),
    .O(__2240__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5621__ (
    .I5(g35),
    .I4(__1712__),
    .I3(__1853__),
    .I2(__323__),
    .I1(__1047__),
    .I0(__1391__),
    .O(__2241__)
  );
  LUT5 #(
    .INIT(32'hd2dd0000)
  ) __5622__ (
    .I4(g35),
    .I3(__1248__),
    .I2(__1245__),
    .I1(__2056__),
    .I0(__154__),
    .O(__2242__)
  );
  LUT5 #(
    .INIT(32'haa3cf0f0)
  ) __5623__ (
    .I4(g35),
    .I3(__803__),
    .I2(__436__),
    .I1(__1687__),
    .I0(__1271__),
    .O(__2243__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __5624__ (
    .I2(g35),
    .I1(__399__),
    .I0(__932__),
    .O(__2244__)
  );
  LUT5 #(
    .INIT(32'hff44f0f0)
  ) __5625__ (
    .I4(g35),
    .I3(__384__),
    .I2(__550__),
    .I1(__1142__),
    .I0(__448__),
    .O(__2245__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __5626__ (
    .I2(__648__),
    .I1(__1156__),
    .I0(__1258__),
    .O(__2246__)
  );
  LUT6 #(
    .INIT(64'hebaa00aa00000000)
  ) __5627__ (
    .I5(g35),
    .I4(__1608__),
    .I3(__1896__),
    .I2(__870__),
    .I1(__2246__),
    .I0(__577__),
    .O(__2247__)
  );
  LUT6 #(
    .INIT(64'hfefeff00ff00ff00)
  ) __5628__ (
    .I5(g35),
    .I4(__341__),
    .I3(__1196__),
    .I2(g72),
    .I1(g73),
    .I0(__25__),
    .O(__2248__)
  );
  LUT5 #(
    .INIT(32'hccaaf0f0)
  ) __5629__ (
    .I4(g35),
    .I3(__1864__),
    .I2(__410__),
    .I1(__330__),
    .I0(__34__),
    .O(__2249__)
  );
  LUT6 #(
    .INIT(64'hf055f0f0cccccccc)
  ) __5630__ (
    .I5(g35),
    .I4(__1349__),
    .I3(__179__),
    .I2(__1023__),
    .I1(__763__),
    .I0(__1344__),
    .O(__2250__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5631__ (
    .I5(g35),
    .I4(__898__),
    .I3(__1632__),
    .I2(__311__),
    .I1(__1229__),
    .I0(__1391__),
    .O(__2251__)
  );
  LUT6 #(
    .INIT(64'h96696996ffffffff)
  ) __5632__ (
    .I5(__680__),
    .I4(__2121__),
    .I3(__2109__),
    .I2(__2096__),
    .I1(__2082__),
    .I0(__2152__),
    .O(__2252__)
  );
  LUT6 #(
    .INIT(64'haaaaaaaccccccccc)
  ) __5633__ (
    .I5(g35),
    .I4(__595__),
    .I3(__112__),
    .I2(__1521__),
    .I1(__58__),
    .I0(__829__),
    .O(__2253__)
  );
  LUT5 #(
    .INIT(32'h7fff0000)
  ) __5634__ (
    .I4(__706__),
    .I3(__282__),
    .I2(__132__),
    .I1(__1672__),
    .I0(__125__),
    .O(__2254__)
  );
  LUT4 #(
    .INIT(16'h8000)
  ) __5635__ (
    .I3(__644__),
    .I2(__816__),
    .I1(__726__),
    .I0(__830__),
    .O(__2255__)
  );
  LUT5 #(
    .INIT(32'hbf80aaaa)
  ) __5636__ (
    .I4(g35),
    .I3(__61__),
    .I2(__2255__),
    .I1(__2254__),
    .I0(__434__),
    .O(__2256__)
  );
  LUT6 #(
    .INIT(64'h0000000000008000)
  ) __5637__ (
    .I5(__465__),
    .I4(__842__),
    .I3(__1227__),
    .I2(__917__),
    .I1(__353__),
    .I0(__972__),
    .O(__2257__)
  );
  LUT6 #(
    .INIT(64'hcf03cf03cf038b8b)
  ) __5638__ (
    .I5(g113),
    .I4(__1283__),
    .I3(__348__),
    .I2(__1000__),
    .I1(__2257__),
    .I0(__1098__),
    .O(__2258__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __5639__ (
    .I2(g35),
    .I1(__2258__),
    .I0(__503__),
    .O(__2259__)
  );
  LUT3 #(
    .INIT(8'h08)
  ) __5640__ (
    .I2(__660__),
    .I1(__881__),
    .I0(__580__),
    .O(__2260__)
  );
  LUT6 #(
    .INIT(64'hdfff7555aaaa0000)
  ) __5641__ (
    .I5(__1160__),
    .I4(__710__),
    .I3(__152__),
    .I2(__2260__),
    .I1(__985__),
    .I0(g35),
    .O(__2261__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5642__ (
    .I5(g35),
    .I4(__1743__),
    .I3(__1660__),
    .I2(__24__),
    .I1(__1015__),
    .I0(__1391__),
    .O(__2262__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5643__ (
    .I1(__688__),
    .I0(__636__),
    .O(__2263__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __5644__ (
    .I1(__874__),
    .I0(__1264__),
    .O(__2264__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5645__ (
    .I5(g35),
    .I4(__2264__),
    .I3(__2263__),
    .I2(__879__),
    .I1(__558__),
    .I0(__1391__),
    .O(__2265__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __5646__ (
    .I1(__561__),
    .I0(__863__),
    .O(__2266__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5647__ (
    .I5(g35),
    .I4(__157__),
    .I3(__2266__),
    .I2(__255__),
    .I1(__57__),
    .I0(__1391__),
    .O(__2267__)
  );
  LUT4 #(
    .INIT(16'h8000)
  ) __5648__ (
    .I3(__917__),
    .I2(__972__),
    .I1(__1444__),
    .I0(__1995__),
    .O(__2268__)
  );
  LUT5 #(
    .INIT(32'hffa0cfc0)
  ) __5649__ (
    .I4(__1383__),
    .I3(__964__),
    .I2(g35),
    .I1(__1114__),
    .I0(__2268__),
    .O(__2269__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __5650__ (
    .I2(__764__),
    .I1(__880__),
    .I0(__1454__),
    .O(__2270__)
  );
  LUT6 #(
    .INIT(64'h6c206c6cf0f0f0f0)
  ) __5651__ (
    .I5(g35),
    .I4(__751__),
    .I3(__869__),
    .I2(__207__),
    .I1(__1113__),
    .I0(__2270__),
    .O(__2271__)
  );
  LUT6 #(
    .INIT(64'h0000007f00000000)
  ) __5652__ (
    .I5(g35),
    .I4(__791__),
    .I3(__898__),
    .I2(__1773__),
    .I1(__1303__),
    .I0(__810__),
    .O(__2272__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5653__ (
    .I1(g35),
    .I0(__270__),
    .O(__2273__)
  );
  LUT6 #(
    .INIT(64'h00dfdf00ffff0000)
  ) __5654__ (
    .I5(g35),
    .I4(__1145__),
    .I3(__1034__),
    .I2(__1303__),
    .I1(__810__),
    .I0(__1302__),
    .O(__2274__)
  );
  LUT6 #(
    .INIT(64'h00088888cccccccc)
  ) __5655__ (
    .I5(g35),
    .I4(__1041__),
    .I3(__1207__),
    .I2(__936__),
    .I1(__997__),
    .I0(__1663__),
    .O(__2275__)
  );
  LUT6 #(
    .INIT(64'heaaa2aaaffff0000)
  ) __5656__ (
    .I5(g35),
    .I4(__308__),
    .I3(__769__),
    .I2(__1286__),
    .I1(__982__),
    .I0(__597__),
    .O(__2276__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5657__ (
    .I5(g35),
    .I4(__2264__),
    .I3(__1704__),
    .I2(__268__),
    .I1(__326__),
    .I0(__1391__),
    .O(__2277__)
  );
  LUT5 #(
    .INIT(32'haaf030f0)
  ) __5658__ (
    .I4(__1782__),
    .I3(g35),
    .I2(__908__),
    .I1(__1779__),
    .I0(__1111__),
    .O(__2278__)
  );
  LUT6 #(
    .INIT(64'hc0c0c0cd00000000)
  ) __5659__ (
    .I5(g35),
    .I4(__645__),
    .I3(__2215__),
    .I2(__1473__),
    .I1(__950__),
    .I0(__1014__),
    .O(__2279__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5660__ (
    .I5(g35),
    .I4(__1728__),
    .I3(__1612__),
    .I2(__404__),
    .I1(__1166__),
    .I0(__1391__),
    .O(__2280__)
  );
  LUT5 #(
    .INIT(32'h80000000)
  ) __5661__ (
    .I4(__1217__),
    .I3(__840__),
    .I2(__1211__),
    .I1(__46__),
    .I0(__1678__),
    .O(__2281__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5662__ (
    .I1(__46__),
    .I0(__1211__),
    .O(__2282__)
  );
  LUT6 #(
    .INIT(64'h0fffffffffff7777)
  ) __5663__ (
    .I5(__1211__),
    .I4(__46__),
    .I3(__935__),
    .I2(__323__),
    .I1(__1162__),
    .I0(__1266__),
    .O(__2283__)
  );
  LUT6 #(
    .INIT(64'h7f00000000007f00)
  ) __5664__ (
    .I5(__840__),
    .I4(__451__),
    .I3(__2283__),
    .I2(__2282__),
    .I1(__302__),
    .I0(__1047__),
    .O(__2284__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5665__ (
    .I1(__1211__),
    .I0(__46__),
    .O(__2285__)
  );
  LUT6 #(
    .INIT(64'hffff0fffffff7777)
  ) __5666__ (
    .I5(__46__),
    .I4(__1211__),
    .I3(__1088__),
    .I2(__1162__),
    .I1(__782__),
    .I0(__302__),
    .O(__2286__)
  );
  LUT6 #(
    .INIT(64'h00007f007f000000)
  ) __5667__ (
    .I5(__840__),
    .I4(__451__),
    .I3(__2286__),
    .I2(__935__),
    .I1(__2285__),
    .I0(__849__),
    .O(__2287__)
  );
  LUT4 #(
    .INIT(16'h8000)
  ) __5668__ (
    .I3(__1217__),
    .I2(__840__),
    .I1(__1211__),
    .I0(__46__),
    .O(__2288__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5669__ (
    .I1(__841__),
    .I0(__366__),
    .O(__2289__)
  );
  LUT6 #(
    .INIT(64'h007f7f7f00000000)
  ) __5670__ (
    .I5(__840__),
    .I4(__2282__),
    .I3(__2289__),
    .I2(__1571__),
    .I1(__283__),
    .I0(__1222__),
    .O(__2290__)
  );
  LUT6 #(
    .INIT(64'h000000f800000088)
  ) __5671__ (
    .I5(__1038__),
    .I4(__1211__),
    .I3(__46__),
    .I2(__1239__),
    .I1(__1172__),
    .I0(__1136__),
    .O(__2291__)
  );
  LUT6 #(
    .INIT(64'h000007770000ffff)
  ) __5672__ (
    .I5(__2285__),
    .I4(__2291__),
    .I3(__774__),
    .I2(__1096__),
    .I1(__451__),
    .I0(__1246__),
    .O(__2292__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __5673__ (
    .I1(__1211__),
    .I0(__46__),
    .O(__2293__)
  );
  LUT6 #(
    .INIT(64'h0000f88800000000)
  ) __5674__ (
    .I5(__46__),
    .I4(__1211__),
    .I3(__1038__),
    .I2(__1075__),
    .I1(__1172__),
    .I0(__1215__),
    .O(__2294__)
  );
  LUT6 #(
    .INIT(64'h0000f88800000000)
  ) __5675__ (
    .I5(__1211__),
    .I4(__46__),
    .I3(__1217__),
    .I2(__748__),
    .I1(__1222__),
    .I0(__1151__),
    .O(__2295__)
  );
  LUT6 #(
    .INIT(64'h000007770000ffff)
  ) __5676__ (
    .I5(__1571__),
    .I4(__2295__),
    .I3(__774__),
    .I2(__1259__),
    .I1(__451__),
    .I0(__1086__),
    .O(__2296__)
  );
  LUT6 #(
    .INIT(64'h0000007f00000000)
  ) __5677__ (
    .I5(__2296__),
    .I4(__840__),
    .I3(__2294__),
    .I2(__2293__),
    .I1(__568__),
    .I0(__366__),
    .O(__2297__)
  );
  LUT3 #(
    .INIT(8'h07)
  ) __5678__ (
    .I2(__2297__),
    .I1(__2292__),
    .I0(__2290__),
    .O(__2298__)
  );
  LUT6 #(
    .INIT(64'hfffff11100000000)
  ) __5679__ (
    .I5(__1678__),
    .I4(__2298__),
    .I3(__2288__),
    .I2(__740__),
    .I1(__2287__),
    .I0(__2284__),
    .O(__2299__)
  );
  LUT5 #(
    .INIT(32'hcf30aaaa)
  ) __5680__ (
    .I4(g35),
    .I3(__2299__),
    .I2(__1234__),
    .I1(__2281__),
    .I0(__178__),
    .O(__2300__)
  );
  LUT5 #(
    .INIT(32'hbfff0000)
  ) __5681__ (
    .I4(__124__),
    .I3(__132__),
    .I2(__1672__),
    .I1(__409__),
    .I0(__282__),
    .O(__2301__)
  );
  LUT6 #(
    .INIT(64'h0000000000008000)
  ) __5682__ (
    .I5(__1240__),
    .I4(__1236__),
    .I3(__1567__),
    .I2(__1052__),
    .I1(__2301__),
    .I0(__1338__),
    .O(__2302__)
  );
  LUT5 #(
    .INIT(32'h05f0cccc)
  ) __5683__ (
    .I4(g35),
    .I3(__2301__),
    .I2(__1126__),
    .I1(__1261__),
    .I0(__2302__),
    .O(__2303__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5684__ (
    .I1(__704__),
    .I0(__468__),
    .O(__2304__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5685__ (
    .I5(g35),
    .I4(__1880__),
    .I3(__2304__),
    .I2(__1176__),
    .I1(__309__),
    .I0(__1391__),
    .O(__2305__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5686__ (
    .I5(g35),
    .I4(__1621__),
    .I3(__1742__),
    .I2(__714__),
    .I1(__911__),
    .I0(__1391__),
    .O(__2306__)
  );
  LUT6 #(
    .INIT(64'h0000413000000c4d)
  ) __5687__ (
    .I5(__343__),
    .I4(g135),
    .I3(__114__),
    .I2(__871__),
    .I1(__92__),
    .I0(__301__),
    .O(__2307__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __5688__ (
    .I1(__1052__),
    .I0(__1236__),
    .O(__2308__)
  );
  LUT6 #(
    .INIT(64'h0000fbf000000000)
  ) __5689__ (
    .I5(__2308__),
    .I4(__702__),
    .I3(__1689__),
    .I2(__738__),
    .I1(__976__),
    .I0(__1271__),
    .O(__2309__)
  );
  LUT6 #(
    .INIT(64'hff000f00ff00bb00)
  ) __5690__ (
    .I5(__738__),
    .I4(__976__),
    .I3(__2309__),
    .I2(__1240__),
    .I1(g90),
    .I0(__1012__),
    .O(__2310__)
  );
  LUT5 #(
    .INIT(32'h0dfdfdcc)
  ) __5691__ (
    .I4(__1052__),
    .I3(__1236__),
    .I2(__702__),
    .I1(__2310__),
    .I0(__2307__),
    .O(__2311__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __5692__ (
    .I2(g35),
    .I1(__2311__),
    .I0(__1168__),
    .O(__2312__)
  );
  LUT6 #(
    .INIT(64'h7f80f0f0fffff0f0)
  ) __5693__ (
    .I5(__650__),
    .I4(g35),
    .I3(__851__),
    .I2(__591__),
    .I1(__353__),
    .I0(__1463__),
    .O(__2313__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5694__ (
    .I1(__908__),
    .I0(__1782__),
    .O(__2314__)
  );
  LUT6 #(
    .INIT(64'hf055f0f0cccccccc)
  ) __5695__ (
    .I5(g35),
    .I4(__2314__),
    .I3(__860__),
    .I2(__690__),
    .I1(__111__),
    .I0(__2034__),
    .O(__2315__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5696__ (
    .I1(g35),
    .I0(__310__),
    .O(__2316__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __5697__ (
    .I2(__1180__),
    .I1(__514__),
    .I0(__1092__),
    .O(__2317__)
  );
  LUT5 #(
    .INIT(32'h00000080)
  ) __5698__ (
    .I4(__69__),
    .I3(__721__),
    .I2(__1077__),
    .I1(__288__),
    .I0(__788__),
    .O(__2318__)
  );
  LUT6 #(
    .INIT(64'hebaa00aa00000000)
  ) __5699__ (
    .I5(g35),
    .I4(__2318__),
    .I3(__1438__),
    .I2(__691__),
    .I1(__2317__),
    .I0(__229__),
    .O(__2319__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __5700__ (
    .I1(__944__),
    .I0(__1600__),
    .O(__2320__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5701__ (
    .I5(g35),
    .I4(__1027__),
    .I3(__2320__),
    .I2(__927__),
    .I1(__1109__),
    .I0(__1597__),
    .O(__2321__)
  );
  LUT6 #(
    .INIT(64'hf055f0f0cccccccc)
  ) __5702__ (
    .I5(g35),
    .I4(__1605__),
    .I3(__352__),
    .I2(__1241__),
    .I1(__988__),
    .I0(__1552__),
    .O(__2322__)
  );
  LUT6 #(
    .INIT(64'h5adaaa2affff0000)
  ) __5703__ (
    .I5(g35),
    .I4(__974__),
    .I3(__711__),
    .I2(__1718__),
    .I1(__91__),
    .I0(__708__),
    .O(__2323__)
  );
  LUT6 #(
    .INIT(64'h0000000080000000)
  ) __5704__ (
    .I5(__1817__),
    .I4(__633__),
    .I3(__126__),
    .I2(__587__),
    .I1(__497__),
    .I0(__1808__),
    .O(__2324__)
  );
  LUT6 #(
    .INIT(64'h45aa45aaffff0000)
  ) __5705__ (
    .I5(g35),
    .I4(__126__),
    .I3(__175__),
    .I2(__973__),
    .I1(__279__),
    .I0(__2324__),
    .O(__2325__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __5706__ (
    .I2(__1766__),
    .I1(__671__),
    .I0(__480__),
    .O(__2326__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5707__ (
    .I5(g35),
    .I4(__1625__),
    .I3(__1558__),
    .I2(__67__),
    .I1(__150__),
    .I0(__1391__),
    .O(__2327__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __5708__ (
    .I2(g35),
    .I1(__1186__),
    .I0(__1143__),
    .O(__2328__)
  );
  LUT4 #(
    .INIT(16'h8000)
  ) __5709__ (
    .I3(__1503__),
    .I2(__779__),
    .I1(__1780__),
    .I0(__1404__),
    .O(__2329__)
  );
  LUT6 #(
    .INIT(64'h0ff0aaaacccccccc)
  ) __5710__ (
    .I5(g35),
    .I4(__2329__),
    .I3(__1060__),
    .I2(__1403__),
    .I1(__860__),
    .I0(__753__),
    .O(__2330__)
  );
  LUT5 #(
    .INIT(32'hbfff0000)
  ) __5711__ (
    .I4(g35),
    .I3(__1110__),
    .I2(__762__),
    .I1(__1251__),
    .I0(__1043__),
    .O(__2331__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __5712__ (
    .I2(__2331__),
    .I1(__127__),
    .I0(__446__),
    .O(__2332__)
  );
  LUT5 #(
    .INIT(32'h96696996)
  ) __5713__ (
    .I4(__2121__),
    .I3(__2109__),
    .I2(__2096__),
    .I1(__2082__),
    .I0(__2152__),
    .O(__2333__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __5714__ (
    .I2(__1766__),
    .I1(__700__),
    .I0(__949__),
    .O(__2334__)
  );
  LUT6 #(
    .INIT(64'h0000000000000080)
  ) __5715__ (
    .I5(__445__),
    .I4(__519__),
    .I3(__1224__),
    .I2(__1190__),
    .I1(__614__),
    .I0(__1615__),
    .O(__2335__)
  );
  LUT5 #(
    .INIT(32'hccaaf0f0)
  ) __5716__ (
    .I4(g35),
    .I3(__2335__),
    .I2(__1065__),
    .I1(__1108__),
    .I0(__975__),
    .O(__2336__)
  );
  LUT6 #(
    .INIT(64'haaaaaaaccccccccc)
  ) __5717__ (
    .I5(g35),
    .I4(__950__),
    .I3(__645__),
    .I2(__1473__),
    .I1(__632__),
    .I0(__1139__),
    .O(__2337__)
  );
  LUT6 #(
    .INIT(64'heaaa2aaaffff0000)
  ) __5718__ (
    .I5(g35),
    .I4(__578__),
    .I3(__1643__),
    .I2(__191__),
    .I1(__958__),
    .I0(__1104__),
    .O(__2338__)
  );
  LUT6 #(
    .INIT(64'h112055a0f0f0f0f0)
  ) __5719__ (
    .I5(g35),
    .I4(__1696__),
    .I3(__347__),
    .I2(__452__),
    .I1(__1396__),
    .I0(__1859__),
    .O(__2339__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5720__ (
    .I1(__1014__),
    .I0(__1473__),
    .O(__2340__)
  );
  LUT6 #(
    .INIT(64'hf055f0f0cccccccc)
  ) __5721__ (
    .I5(g35),
    .I4(__2340__),
    .I3(__950__),
    .I2(__834__),
    .I1(__828__),
    .I0(__1470__),
    .O(__2341__)
  );
  LUT4 #(
    .INIT(16'h77f0)
  ) __5722__ (
    .I3(g35),
    .I2(__200__),
    .I1(__752__),
    .I0(__614__),
    .O(__2342__)
  );
  LUT5 #(
    .INIT(32'h80000000)
  ) __5723__ (
    .I4(__833__),
    .I3(__62__),
    .I2(__1154__),
    .I1(__1126__),
    .I0(__2301__),
    .O(__2343__)
  );
  LUT5 #(
    .INIT(32'h3caaf0f0)
  ) __5724__ (
    .I4(g35),
    .I3(__2343__),
    .I2(__960__),
    .I1(__240__),
    .I0(__918__),
    .O(__2344__)
  );
  LUT6 #(
    .INIT(64'hccccf0aaf0f0f0f0)
  ) __5725__ (
    .I5(g35),
    .I4(__2179__),
    .I3(__1943__),
    .I2(__1084__),
    .I1(__1279__),
    .I0(__222__),
    .O(__2345__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5726__ (
    .I1(__413__),
    .I0(__116__),
    .O(__2346__)
  );
  LUT6 #(
    .INIT(64'h331100001f3f0000)
  ) __5727__ (
    .I5(__631__),
    .I4(__437__),
    .I3(__299__),
    .I2(__736__),
    .I1(__2346__),
    .I0(__1029__),
    .O(__2347__)
  );
  LUT6 #(
    .INIT(64'hafaaeaaaff00ff00)
  ) __5728__ (
    .I5(g35),
    .I4(__631__),
    .I3(__35__),
    .I2(__299__),
    .I1(__736__),
    .I0(__2347__),
    .O(__2348__)
  );
  LUT4 #(
    .INIT(16'hbbf0)
  ) __5729__ (
    .I3(g35),
    .I2(__467__),
    .I1(g91),
    .I0(__822__),
    .O(__2349__)
  );
  LUT3 #(
    .INIT(8'he0)
  ) __5730__ (
    .I2(__1115__),
    .I1(__35__),
    .I0(__437__),
    .O(__2350__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5731__ (
    .I1(__777__),
    .I0(__1665__),
    .O(__2351__)
  );
  LUT6 #(
    .INIT(64'h4000ffff00000000)
  ) __5732__ (
    .I5(__687__),
    .I4(g35),
    .I3(__211__),
    .I2(__197__),
    .I1(__2351__),
    .I0(__2350__),
    .O(__2352__)
  );
  LUT5 #(
    .INIT(32'h00000008)
  ) __5733__ (
    .I4(__972__),
    .I3(g113),
    .I2(__1283__),
    .I1(__1430__),
    .I0(__1465__),
    .O(__2353__)
  );
  LUT6 #(
    .INIT(64'hf30caaaaf0f0f0f0)
  ) __5734__ (
    .I5(g35),
    .I4(__2353__),
    .I3(__749__),
    .I2(__23__),
    .I1(__142__),
    .I0(__957__),
    .O(__2354__)
  );
  LUT5 #(
    .INIT(32'hacaacccc)
  ) __5735__ (
    .I4(g35),
    .I3(__1531__),
    .I2(__1476__),
    .I1(__579__),
    .I0(__1228__),
    .O(__2355__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __5736__ (
    .I2(__952__),
    .I1(__206__),
    .I0(__878__),
    .O(__2356__)
  );
  LUT5 #(
    .INIT(32'h0000002c)
  ) __5737__ (
    .I4(__35__),
    .I3(__437__),
    .I2(__299__),
    .I1(__631__),
    .I0(__736__),
    .O(__2357__)
  );
  LUT6 #(
    .INIT(64'h00000000000000f7)
  ) __5738__ (
    .I5(__168__),
    .I4(__1009__),
    .I3(__484__),
    .I2(__2357__),
    .I1(__992__),
    .I0(__2356__),
    .O(__2358__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5739__ (
    .I1(g35),
    .I0(__2358__),
    .O(__2359__)
  );
  LUT5 #(
    .INIT(32'h00cef0f0)
  ) __5740__ (
    .I4(g35),
    .I3(__1130__),
    .I2(__213__),
    .I1(__730__),
    .I0(__859__),
    .O(__2360__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5741__ (
    .I1(__253__),
    .I0(__689__),
    .O(__2361__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5742__ (
    .I5(g35),
    .I4(__2361__),
    .I3(__1612__),
    .I2(__162__),
    .I1(__1218__),
    .I0(__1391__),
    .O(__2362__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5743__ (
    .I1(__120__),
    .I0(__463__),
    .O(__2363__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5744__ (
    .I5(g35),
    .I4(__2000__),
    .I3(__2363__),
    .I2(__487__),
    .I1(__119__),
    .I0(__1391__),
    .O(__2364__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5745__ (
    .I1(__881__),
    .I0(__660__),
    .O(__2365__)
  );
  LUT6 #(
    .INIT(64'h06660066ffff0000)
  ) __5746__ (
    .I5(g35),
    .I4(__1115__),
    .I3(__1975__),
    .I2(__2365__),
    .I1(__134__),
    .I0(__1973__),
    .O(__2366__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __5747__ (
    .I1(__489__),
    .I0(__88__),
    .O(__2367__)
  );
  LUT5 #(
    .INIT(32'habff5400)
  ) __5748__ (
    .I4(__1189__),
    .I3(__1041__),
    .I2(__1207__),
    .I1(__936__),
    .I0(__983__),
    .O(__2368__)
  );
  LUT6 #(
    .INIT(64'hfa00f0f0cccccccc)
  ) __5749__ (
    .I5(g35),
    .I4(__1602__),
    .I3(__2368__),
    .I2(__107__),
    .I1(__245__),
    .I0(__2367__),
    .O(__2369__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __5750__ (
    .I2(__1766__),
    .I1(__184__),
    .I0(__783__),
    .O(__2370__)
  );
  LUT3 #(
    .INIT(8'h08)
  ) __5751__ (
    .I2(__596__),
    .I1(__639__),
    .I0(__163__),
    .O(__2371__)
  );
  LUT6 #(
    .INIT(64'h000001ff00000000)
  ) __5752__ (
    .I5(__1249__),
    .I4(__1540__),
    .I3(__2371__),
    .I2(__942__),
    .I1(__127__),
    .I0(__446__),
    .O(__2372__)
  );
  LUT6 #(
    .INIT(64'h8000000000000000)
  ) __5753__ (
    .I5(__2371__),
    .I4(__2372__),
    .I3(__641__),
    .I2(__955__),
    .I1(__1203__),
    .I0(__277__),
    .O(__2373__)
  );
  LUT4 #(
    .INIT(16'h8f00)
  ) __5754__ (
    .I3(__510__),
    .I2(g35),
    .I1(__575__),
    .I0(__2373__),
    .O(__2374__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5755__ (
    .I5(g35),
    .I4(__623__),
    .I3(__1611__),
    .I2(__858__),
    .I1(__805__),
    .I0(__1391__),
    .O(__2375__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __5756__ (
    .I2(g35),
    .I1(__356__),
    .I0(__161__),
    .O(__2376__)
  );
  LUT2 #(
    .INIT(4'h2)
  ) __5757__ (
    .I1(__824__),
    .I0(g73),
    .O(__2377__)
  );
  LUT6 #(
    .INIT(64'h7777f0f0ff00ff00)
  ) __5758__ (
    .I5(g35),
    .I4(__341__),
    .I3(__785__),
    .I2(__655__),
    .I1(g72),
    .I0(__2377__),
    .O(__2378__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5759__ (
    .I5(g35),
    .I4(__1965__),
    .I3(__1793__),
    .I2(__570__),
    .I1(__1090__),
    .I0(__1391__),
    .O(__2379__)
  );
  LUT6 #(
    .INIT(64'h2aaad55500000000)
  ) __5760__ (
    .I5(g35),
    .I4(__1391__),
    .I3(__468__),
    .I2(__704__),
    .I1(__898__),
    .I0(__76__),
    .O(__2380__)
  );
  LUT6 #(
    .INIT(64'hffff44f400f000f0)
  ) __5761__ (
    .I5(__1389__),
    .I4(__611__),
    .I3(g35),
    .I2(__348__),
    .I1(__1388__),
    .I0(__1116__),
    .O(__2381__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5762__ (
    .I1(__418__),
    .I0(__1173__),
    .O(__2382__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5763__ (
    .I5(g35),
    .I4(__2382__),
    .I3(__1874__),
    .I2(__601__),
    .I1(__598__),
    .I0(__1391__),
    .O(__2383__)
  );
  LUT4 #(
    .INIT(16'heef0)
  ) __5764__ (
    .I3(g35),
    .I2(__563__),
    .I1(__529__),
    .I0(__1250__),
    .O(__2384__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5765__ (
    .I1(__769__),
    .I0(__982__),
    .O(__2385__)
  );
  LUT6 #(
    .INIT(64'hc3aaaaaaf0f0f0f0)
  ) __5766__ (
    .I5(g35),
    .I4(__1286__),
    .I3(__2385__),
    .I2(__597__),
    .I1(__308__),
    .I0(__928__),
    .O(__2386__)
  );
  LUT6 #(
    .INIT(64'hdfffffffcfffffff)
  ) __5767__ (
    .I5(__1370__),
    .I4(__680__),
    .I3(__1934__),
    .I2(__1933__),
    .I1(__1929__),
    .I0(__1924__),
    .O(__2387__)
  );
  LUT6 #(
    .INIT(64'hf055f0f0cccccccc)
  ) __5768__ (
    .I5(g35),
    .I4(__2314__),
    .I3(__1111__),
    .I2(__1122__),
    .I1(__336__),
    .I0(__2034__),
    .O(__2388__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __5769__ (
    .I2(__2331__),
    .I1(__843__),
    .I0(__627__),
    .O(__2389__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5770__ (
    .I5(g35),
    .I4(__157__),
    .I3(__2026__),
    .I2(__176__),
    .I1(__1129__),
    .I0(__1391__),
    .O(__2390__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __5771__ (
    .I2(g35),
    .I1(__1147__),
    .I0(__262__),
    .O(__2391__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __5772__ (
    .I2(g35),
    .I1(__363__),
    .I0(__316__),
    .O(__2392__)
  );
  LUT6 #(
    .INIT(64'h00002300f0f0f0f0)
  ) __5773__ (
    .I5(g35),
    .I4(__182__),
    .I3(__1533__),
    .I2(__83__),
    .I1(__1538__),
    .I0(__1535__),
    .O(__2393__)
  );
  LUT6 #(
    .INIT(64'h45aa45aaffff0000)
  ) __5774__ (
    .I5(g35),
    .I4(__854__),
    .I3(__981__),
    .I2(__751__),
    .I1(__869__),
    .I0(__1455__),
    .O(__2394__)
  );
  LUT3 #(
    .INIT(8'hd0)
  ) __5775__ (
    .I2(__407__),
    .I1(__869__),
    .I0(__751__),
    .O(__2395__)
  );
  LUT5 #(
    .INIT(32'h7fd5aa00)
  ) __5776__ (
    .I4(__199__),
    .I3(__2395__),
    .I2(__744__),
    .I1(__1456__),
    .I0(g35),
    .O(__2396__)
  );
  LUT6 #(
    .INIT(64'hdfff7555aaaa0000)
  ) __5777__ (
    .I5(__107__),
    .I4(__1189__),
    .I3(__88__),
    .I2(__1602__),
    .I1(__835__),
    .I0(g35),
    .O(__2397__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5778__ (
    .I1(__1036__),
    .I0(__1275__),
    .O(__2398__)
  );
  LUT6 #(
    .INIT(64'hf0ff00ffffff7777)
  ) __5779__ (
    .I5(__1207__),
    .I4(__1812__),
    .I3(__1545__),
    .I2(__594__),
    .I1(__1105__),
    .I0(__2398__),
    .O(__2399__)
  );
  LUT6 #(
    .INIT(64'hf57f554400000000)
  ) __5780__ (
    .I5(g35),
    .I4(__936__),
    .I3(__544__),
    .I2(__396__),
    .I1(__646__),
    .I0(__2399__),
    .O(__2400__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __5781__ (
    .I2(g35),
    .I1(g6749),
    .I0(__882__),
    .O(__2401__)
  );
  LUT6 #(
    .INIT(64'h0000000000000004)
  ) __5782__ (
    .I5(__1103__),
    .I4(__485__),
    .I3(__284__),
    .I2(__192__),
    .I1(__659__),
    .I0(__481__),
    .O(__2402__)
  );
  LUT4 #(
    .INIT(16'hefa0)
  ) __5783__ (
    .I3(__284__),
    .I2(g35),
    .I1(__479__),
    .I0(__2402__),
    .O(__2403__)
  );
  LUT5 #(
    .INIT(32'hcceccccc)
  ) __5784__ (
    .I4(g35),
    .I3(__659__),
    .I2(__1757__),
    .I1(__685__),
    .I0(__604__),
    .O(__2404__)
  );
  LUT6 #(
    .INIT(64'h7f33b3b3cc000000)
  ) __5785__ (
    .I5(__890__),
    .I4(__496__),
    .I3(__1147__),
    .I2(__592__),
    .I1(g35),
    .I0(__1662__),
    .O(__2405__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __5786__ (
    .I2(g35),
    .I1(__54__),
    .I0(__638__),
    .O(__2406__)
  );
  LUT6 #(
    .INIT(64'h3fffc000aaaaaaaa)
  ) __5787__ (
    .I5(g35),
    .I4(__355__),
    .I3(__1164__),
    .I2(__964__),
    .I1(__1383__),
    .I0(__844__),
    .O(__2407__)
  );
  LUT6 #(
    .INIT(64'h333f33b300cc0000)
  ) __5788__ (
    .I5(__976__),
    .I4(__738__),
    .I3(__1776__),
    .I2(__1775__),
    .I1(g35),
    .I0(__1240__),
    .O(__2408__)
  );
  LUT6 #(
    .INIT(64'h000000ff0000efef)
  ) __5789__ (
    .I5(__1732__),
    .I4(__1638__),
    .I3(__804__),
    .I2(__1248__),
    .I1(__1342__),
    .I0(__1637__),
    .O(__2409__)
  );
  LUT6 #(
    .INIT(64'h6666666affff0000)
  ) __5790__ (
    .I5(g35),
    .I4(__318__),
    .I3(__1269__),
    .I2(__1638__),
    .I1(__1238__),
    .I0(__2409__),
    .O(__2410__)
  );
  LUT2 #(
    .INIT(4'h7)
  ) __5791__ (
    .I1(g113),
    .I0(__932__),
    .O(__2411__)
  );
  LUT6 #(
    .INIT(64'h0077ff00f0f0f0f0)
  ) __5792__ (
    .I5(g35),
    .I4(__1896__),
    .I3(__648__),
    .I2(__1156__),
    .I1(__1338__),
    .I0(__1568__),
    .O(__2412__)
  );
  LUT6 #(
    .INIT(64'hbfffffff00000000)
  ) __5793__ (
    .I5(__52__),
    .I4(g35),
    .I3(__1503__),
    .I2(__1567__),
    .I1(__15__),
    .I0(__1240__),
    .O(__2413__)
  );
  LUT6 #(
    .INIT(64'h00ff33330f0f5555)
  ) __5794__ (
    .I5(__795__),
    .I4(__718__),
    .I3(__101__),
    .I2(__1158__),
    .I1(__821__),
    .I0(__9__),
    .O(__2414__)
  );
  LUT6 #(
    .INIT(64'hff00ccccf0f0aaaa)
  ) __5795__ (
    .I5(__795__),
    .I4(__718__),
    .I3(__1178__),
    .I2(__1048__),
    .I1(__537__),
    .I0(__963__),
    .O(__2415__)
  );
  LUT6 #(
    .INIT(64'hefff200000000000)
  ) __5796__ (
    .I5(g35),
    .I4(__2415__),
    .I3(__2210__),
    .I2(__2209__),
    .I1(__1227__),
    .I0(__2414__),
    .O(__2416__)
  );
  LUT3 #(
    .INIT(8'hf4)
  ) __5797__ (
    .I2(__2416__),
    .I1(__868__),
    .I0(g35),
    .O(__2417__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5798__ (
    .I5(g35),
    .I4(__1794__),
    .I3(__1964__),
    .I2(__808__),
    .I1(__883__),
    .I0(__1391__),
    .O(__2418__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __5799__ (
    .I1(__519__),
    .I0(__1224__),
    .O(__2419__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __5800__ (
    .I1(__1190__),
    .I0(__614__),
    .O(__2420__)
  );
  LUT6 #(
    .INIT(64'h000080ff00000000)
  ) __5801__ (
    .I5(__2420__),
    .I4(__1082__),
    .I3(__2419__),
    .I2(__445__),
    .I1(__1025__),
    .I0(__1615__),
    .O(__2421__)
  );
  LUT6 #(
    .INIT(64'hff00df10ffff0000)
  ) __5802__ (
    .I5(g35),
    .I4(__561__),
    .I3(__29__),
    .I2(__2163__),
    .I1(__863__),
    .I0(__1391__),
    .O(__2422__)
  );
  LUT6 #(
    .INIT(64'h0000ff000000efef)
  ) __5803__ (
    .I5(__1979__),
    .I4(__1489__),
    .I3(__666__),
    .I2(__1248__),
    .I1(__1486__),
    .I0(__1485__),
    .O(__2423__)
  );
  LUT6 #(
    .INIT(64'h6666666affff0000)
  ) __5804__ (
    .I5(g35),
    .I4(__196__),
    .I3(__1028__),
    .I2(__1489__),
    .I1(__1002__),
    .I0(__2423__),
    .O(__2424__)
  );
  LUT6 #(
    .INIT(64'h78f070f0ffff0000)
  ) __5805__ (
    .I5(g35),
    .I4(__423__),
    .I3(__952__),
    .I2(__992__),
    .I1(__206__),
    .I0(__878__),
    .O(__2425__)
  );
  LUT4 #(
    .INIT(16'hb8cc)
  ) __5806__ (
    .I3(g35),
    .I2(__448__),
    .I1(__1142__),
    .I0(__384__),
    .O(__2426__)
  );
  LUT4 #(
    .INIT(16'h0001)
  ) __5807__ (
    .I3(__526__),
    .I2(__71__),
    .I1(__945__),
    .I0(__1272__),
    .O(__2427__)
  );
  LUT3 #(
    .INIT(8'h01)
  ) __5808__ (
    .I2(__1112__),
    .I1(__813__),
    .I0(__305__),
    .O(__2428__)
  );
  LUT6 #(
    .INIT(64'h00ffff88f0f0f0f0)
  ) __5809__ (
    .I5(g35),
    .I4(__1248__),
    .I3(__1102__),
    .I2(__249__),
    .I1(__2428__),
    .I0(__2427__),
    .O(__2429__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5810__ (
    .I5(g35),
    .I4(__412__),
    .I3(__1853__),
    .I2(__748__),
    .I1(__1266__),
    .I0(__1391__),
    .O(__2430__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5811__ (
    .I5(g35),
    .I4(__1965__),
    .I3(__1874__),
    .I2(__121__),
    .I1(__513__),
    .I0(__1391__),
    .O(__2431__)
  );
  LUT6 #(
    .INIT(64'h30fcfcb800000000)
  ) __5812__ (
    .I5(g35),
    .I4(__237__),
    .I3(__1648__),
    .I2(__480__),
    .I1(__1649__),
    .I0(__1647__),
    .O(__2432__)
  );
  LUT5 #(
    .INIT(32'h3535ff00)
  ) __5813__ (
    .I4(g35),
    .I3(__1248__),
    .I2(__1204__),
    .I1(__406__),
    .I0(__1108__),
    .O(__2433__)
  );
  LUT2 #(
    .INIT(4'h7)
  ) __5814__ (
    .I1(g113),
    .I0(__399__),
    .O(__2434__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __5815__ (
    .I2(__738__),
    .I1(__976__),
    .I0(__1775__),
    .O(__2435__)
  );
  LUT6 #(
    .INIT(64'h00001cccf0f0f0f0)
  ) __5816__ (
    .I5(g35),
    .I4(__1776__),
    .I3(__2435__),
    .I2(__871__),
    .I1(__343__),
    .I0(__301__),
    .O(__2436__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __5817__ (
    .I2(g35),
    .I1(__932__),
    .I0(__796__),
    .O(__2437__)
  );
  LUT4 #(
    .INIT(16'hbbf0)
  ) __5818__ (
    .I3(g35),
    .I2(__426__),
    .I1(__1249__),
    .I0(__1127__),
    .O(__2438__)
  );
  LUT6 #(
    .INIT(64'hcfcccfcc4544cfcc)
  ) __5819__ (
    .I5(__972__),
    .I4(__1444__),
    .I3(__819__),
    .I2(__769__),
    .I1(__982__),
    .I0(__1459__),
    .O(__2439__)
  );
  LUT5 #(
    .INIT(32'h33aaf0f0)
  ) __5820__ (
    .I4(g35),
    .I3(__1286__),
    .I2(__866__),
    .I1(__2439__),
    .I0(__769__),
    .O(__2440__)
  );
  LUT6 #(
    .INIT(64'h8000000000000000)
  ) __5821__ (
    .I5(__199__),
    .I4(__407__),
    .I3(__981__),
    .I2(__744__),
    .I1(__33__),
    .I0(__1455__),
    .O(__2441__)
  );
  LUT6 #(
    .INIT(64'h6c206c6cf0f0f0f0)
  ) __5822__ (
    .I5(g35),
    .I4(__751__),
    .I3(__869__),
    .I2(__716__),
    .I1(__226__),
    .I0(__2441__),
    .O(__2442__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __5823__ (
    .I2(g35),
    .I1(__276__),
    .I0(__938__),
    .O(__2443__)
  );
  LUT5 #(
    .INIT(32'h575d0a00)
  ) __5824__ (
    .I4(__1126__),
    .I3(__1154__),
    .I2(__2302__),
    .I1(__2301__),
    .I0(g35),
    .O(__2444__)
  );
  LUT4 #(
    .INIT(16'h0080)
  ) __5825__ (
    .I3(__794__),
    .I2(__1268__),
    .I1(__702__),
    .I0(__482__),
    .O(__2445__)
  );
  LUT5 #(
    .INIT(32'h575d0a00)
  ) __5826__ (
    .I4(__1052__),
    .I3(__1236__),
    .I2(__1776__),
    .I1(__2445__),
    .I0(g35),
    .O(__2446__)
  );
  LUT5 #(
    .INIT(32'he8000000)
  ) __5827__ (
    .I4(g35),
    .I3(__2371__),
    .I2(__942__),
    .I1(__127__),
    .I0(__446__),
    .O(__2447__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5828__ (
    .I1(__561__),
    .I0(__863__),
    .O(__2448__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5829__ (
    .I5(g35),
    .I4(__2448__),
    .I3(__1791__),
    .I2(__977__),
    .I1(__79__),
    .I0(__1391__),
    .O(__2449__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5830__ (
    .I1(__791__),
    .I0(__832__),
    .O(__2450__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5831__ (
    .I1(__468__),
    .I0(__704__),
    .O(__2451__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5832__ (
    .I5(g35),
    .I4(__2451__),
    .I3(__2450__),
    .I2(__136__),
    .I1(__281__),
    .I0(__1391__),
    .O(__2452__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5833__ (
    .I1(__252__),
    .I0(__1818__),
    .O(__2453__)
  );
  LUT6 #(
    .INIT(64'h337fb3b300cc0000)
  ) __5834__ (
    .I5(__642__),
    .I4(__459__),
    .I3(__1817__),
    .I2(__790__),
    .I1(g35),
    .I0(__2453__),
    .O(__2454__)
  );
  LUT5 #(
    .INIT(32'hccaaf0f0)
  ) __5835__ (
    .I4(g35),
    .I3(__638__),
    .I2(__664__),
    .I1(g124),
    .I0(g120),
    .O(__2455__)
  );
  LUT5 #(
    .INIT(32'h3cffaaaa)
  ) __5836__ (
    .I4(g35),
    .I3(__650__),
    .I2(__353__),
    .I1(__1463__),
    .I0(__917__),
    .O(__2456__)
  );
  LUT6 #(
    .INIT(64'h6c00cc00aaaaaaaa)
  ) __5837__ (
    .I5(g35),
    .I4(__2371__),
    .I3(__2372__),
    .I2(__955__),
    .I1(__641__),
    .I0(__1203__),
    .O(__2457__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5838__ (
    .I5(g35),
    .I4(__306__),
    .I3(__1620__),
    .I2(__238__),
    .I1(__615__),
    .I0(__1391__),
    .O(__2458__)
  );
  LUT3 #(
    .INIT(8'h01)
  ) __5839__ (
    .I2(__728__),
    .I1(__1348__),
    .I0(__801__),
    .O(__2459__)
  );
  LUT5 #(
    .INIT(32'h33aaf0f0)
  ) __5840__ (
    .I4(g35),
    .I3(__2459__),
    .I2(__1001__),
    .I1(__1344__),
    .I0(__1131__),
    .O(__2460__)
  );
  LUT5 #(
    .INIT(32'h00000008)
  ) __5841__ (
    .I4(g113),
    .I3(__1283__),
    .I2(__779__),
    .I1(__1060__),
    .I0(__1409__),
    .O(__2461__)
  );
  LUT5 #(
    .INIT(32'haaf030f0)
  ) __5842__ (
    .I4(__1638__),
    .I3(g35),
    .I2(__617__),
    .I1(__2461__),
    .I0(__318__),
    .O(__2462__)
  );
  LUT6 #(
    .INIT(64'h557f55d500aa0000)
  ) __5843__ (
    .I5(__1077__),
    .I4(__69__),
    .I3(__1441__),
    .I2(__788__),
    .I1(__1857__),
    .I0(g35),
    .O(__2463__)
  );
  LUT6 #(
    .INIT(64'h0000ffc0aaaaaaaa)
  ) __5844__ (
    .I5(g35),
    .I4(g113),
    .I3(g134),
    .I2(__884__),
    .I1(g99),
    .I0(__479__),
    .O(__2464__)
  );
  LUT4 #(
    .INIT(16'h8000)
  ) __5845__ (
    .I3(__833__),
    .I2(__62__),
    .I1(__1154__),
    .I0(__1126__),
    .O(__2465__)
  );
  LUT5 #(
    .INIT(32'hbf80aaaa)
  ) __5846__ (
    .I4(g35),
    .I3(__1093__),
    .I2(__2465__),
    .I1(__2301__),
    .I0(__658__),
    .O(__2466__)
  );
  LUT5 #(
    .INIT(32'h7fd5aa00)
  ) __5847__ (
    .I4(__1095__),
    .I3(__970__),
    .I2(__734__),
    .I1(__725__),
    .I0(g35),
    .O(__2467__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5848__ (
    .I5(g35),
    .I4(__412__),
    .I3(__1805__),
    .I2(__1215__),
    .I1(__1151__),
    .I0(__1391__),
    .O(__2468__)
  );
  LUT3 #(
    .INIT(8'h70)
  ) __5849__ (
    .I2(__315__),
    .I1(__1522__),
    .I0(__417__),
    .O(__2469__)
  );
  LUT6 #(
    .INIT(64'hcfcccfcc4544cfcc)
  ) __5850__ (
    .I5(__972__),
    .I4(__1444__),
    .I3(__760__),
    .I2(__1197__),
    .I1(__541__),
    .I0(__1298__),
    .O(__2470__)
  );
  LUT5 #(
    .INIT(32'h33aaf0f0)
  ) __5851__ (
    .I4(g35),
    .I3(__1299__),
    .I2(__453__),
    .I1(__2470__),
    .I0(__1197__),
    .O(__2471__)
  );
  LUT5 #(
    .INIT(32'hccaaf0f0)
  ) __5852__ (
    .I4(g35),
    .I3(__170__),
    .I2(__881__),
    .I1(__299__),
    .I0(__204__),
    .O(__2472__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5853__ (
    .I5(g35),
    .I4(__2361__),
    .I3(__1727__),
    .I2(__156__),
    .I1(__51__),
    .I0(__1391__),
    .O(__2473__)
  );
  LUT2 #(
    .INIT(4'h2)
  ) __5854__ (
    .I1(__1269__),
    .I0(__617__),
    .O(__2474__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5855__ (
    .I1(__1114__),
    .I0(__1164__),
    .O(__2475__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5856__ (
    .I5(g35),
    .I4(__1383__),
    .I3(__2475__),
    .I2(__581__),
    .I1(__742__),
    .I0(__2474__),
    .O(__2476__)
  );
  LUT6 #(
    .INIT(64'h0000000000008000)
  ) __5857__ (
    .I5(g113),
    .I4(__1283__),
    .I3(__757__),
    .I2(__236__),
    .I1(__810__),
    .I0(__2054__),
    .O(__2477__)
  );
  LUT5 #(
    .INIT(32'h10ff0000)
  ) __5858__ (
    .I4(__463__),
    .I3(g35),
    .I2(__120__),
    .I1(__306__),
    .I0(__2477__),
    .O(__2478__)
  );
  LUT6 #(
    .INIT(64'hff00df10ffff0000)
  ) __5859__ (
    .I5(g35),
    .I4(__705__),
    .I3(__317__),
    .I2(__1823__),
    .I1(__509__),
    .I0(__1391__),
    .O(__2479__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __5860__ (
    .I2(g35),
    .I1(__214__),
    .I0(__90__),
    .O(__2480__)
  );
  LUT6 #(
    .INIT(64'hc3aaaaaaf0f0f0f0)
  ) __5861__ (
    .I5(g35),
    .I4(__1674__),
    .I3(__1673__),
    .I2(__339__),
    .I1(__1175__),
    .I0(__167__),
    .O(__2481__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5862__ (
    .I5(g35),
    .I4(__2061__),
    .I3(__1853__),
    .I2(__1266__),
    .I1(__323__),
    .I0(__1391__),
    .O(__2482__)
  );
  LUT6 #(
    .INIT(64'hefefff00ff00ff00)
  ) __5863__ (
    .I5(g35),
    .I4(__341__),
    .I3(__603__),
    .I2(g72),
    .I1(g73),
    .I0(__390__),
    .O(__2483__)
  );
  LUT3 #(
    .INIT(8'h01)
  ) __5864__ (
    .I2(__950__),
    .I1(__645__),
    .I0(__1473__),
    .O(__2484__)
  );
  LUT5 #(
    .INIT(32'hc3aaf0f0)
  ) __5865__ (
    .I4(g35),
    .I3(__2484__),
    .I2(__146__),
    .I1(__102__),
    .I0(__1149__),
    .O(__2485__)
  );
  LUT6 #(
    .INIT(64'hccccccacaaaaaaaa)
  ) __5866__ (
    .I5(g35),
    .I4(__507__),
    .I3(__1032__),
    .I2(__709__),
    .I1(__835__),
    .I0(__489__),
    .O(__2486__)
  );
  LUT3 #(
    .INIT(8'h01)
  ) __5867__ (
    .I2(__1269__),
    .I1(__1638__),
    .I0(__318__),
    .O(__2487__)
  );
  LUT5 #(
    .INIT(32'hc3aaf0f0)
  ) __5868__ (
    .I4(g35),
    .I3(__2487__),
    .I2(__978__),
    .I1(__355__),
    .I0(__483__),
    .O(__2488__)
  );
  LUT5 #(
    .INIT(32'h00000008)
  ) __5869__ (
    .I4(g113),
    .I3(__1283__),
    .I2(__779__),
    .I1(__1060__),
    .I0(__1404__),
    .O(__2489__)
  );
  LUT6 #(
    .INIT(64'hf0f04444ff00ff00)
  ) __5870__ (
    .I5(g35),
    .I4(__1600__),
    .I3(__228__),
    .I2(__1027__),
    .I1(__296__),
    .I0(__2489__),
    .O(__2490__)
  );
  LUT4 #(
    .INIT(16'h7580)
  ) __5871__ (
    .I3(__794__),
    .I2(__1432__),
    .I1(__482__),
    .I0(g35),
    .O(__2491__)
  );
  LUT5 #(
    .INIT(32'hc3aaf0f0)
  ) __5872__ (
    .I4(g35),
    .I3(__1506__),
    .I2(__1037__),
    .I1(__1150__),
    .I0(__512__),
    .O(__2492__)
  );
  LUT5 #(
    .INIT(32'h3c00aaaa)
  ) __5873__ (
    .I4(g35),
    .I3(__2372__),
    .I2(__2371__),
    .I1(__955__),
    .I0(__381__),
    .O(__2493__)
  );
  LUT5 #(
    .INIT(32'hf8fff000)
  ) __5874__ (
    .I4(__1031__),
    .I3(g35),
    .I2(__320__),
    .I1(__1757__),
    .I0(__659__),
    .O(__2494__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5875__ (
    .I1(__728__),
    .I0(__179__),
    .O(__2495__)
  );
  LUT4 #(
    .INIT(16'h8000)
  ) __5876__ (
    .I3(__1503__),
    .I2(__779__),
    .I1(__1405__),
    .I0(__1346__),
    .O(__2496__)
  );
  LUT6 #(
    .INIT(64'h0ff0aaaacccccccc)
  ) __5877__ (
    .I5(g35),
    .I4(__2496__),
    .I3(__1060__),
    .I2(__2495__),
    .I1(__801__),
    .I0(__812__),
    .O(__2497__)
  );
  LUT6 #(
    .INIT(64'h3caaaaaaf0f0f0f0)
  ) __5878__ (
    .I5(g35),
    .I4(__712__),
    .I3(__956__),
    .I2(__466__),
    .I1(__294__),
    .I0(__304__),
    .O(__2498__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5879__ (
    .I1(__934__),
    .I0(__1237__),
    .O(__2499__)
  );
  LUT6 #(
    .INIT(64'h77770777ffffffff)
  ) __5880__ (
    .I5(__972__),
    .I4(__784__),
    .I3(__1459__),
    .I2(__469__),
    .I1(__1953__),
    .I0(__2499__),
    .O(__2500__)
  );
  LUT6 #(
    .INIT(64'hffffffff2a3f3f3f)
  ) __5881__ (
    .I5(__972__),
    .I4(__1953__),
    .I3(__1208__),
    .I2(__1459__),
    .I1(__1290__),
    .I0(__191__),
    .O(__2501__)
  );
  LUT6 #(
    .INIT(64'hcfffcfffffff55ff)
  ) __5882__ (
    .I5(__972__),
    .I4(__142__),
    .I3(__1465__),
    .I2(__1114__),
    .I1(__1164__),
    .I0(__23__),
    .O(__2502__)
  );
  LUT6 #(
    .INIT(64'hcfffcfffffff55ff)
  ) __5883__ (
    .I5(__972__),
    .I4(__541__),
    .I3(__1298__),
    .I2(__91__),
    .I1(__13__),
    .I0(__760__),
    .O(__2503__)
  );
  LUT6 #(
    .INIT(64'h7fffffffffffffff)
  ) __5884__ (
    .I5(__1413__),
    .I4(__1443__),
    .I3(__2503__),
    .I2(__2502__),
    .I1(__2501__),
    .I0(__2500__),
    .O(__2504__)
  );
  LUT3 #(
    .INIT(8'h78)
  ) __5885__ (
    .I2(__1068__),
    .I1(g35),
    .I0(__585__),
    .O(__2505__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5886__ (
    .I1(g35),
    .I0(__1068__),
    .O(__2506__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5887__ (
    .I5(g35),
    .I4(__2026__),
    .I3(__2163__),
    .I2(__1161__),
    .I1(__255__),
    .I0(__1391__),
    .O(__2507__)
  );
  LUT4 #(
    .INIT(16'h7fff)
  ) __5888__ (
    .I3(__2503__),
    .I2(__2502__),
    .I1(__2501__),
    .I0(__2500__),
    .O(__2508__)
  );
  LUT6 #(
    .INIT(64'h2aaad55500000000)
  ) __5889__ (
    .I5(g35),
    .I4(__1391__),
    .I3(__313__),
    .I2(__569__),
    .I1(__989__),
    .I0(__643__),
    .O(__2509__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5890__ (
    .I1(g35),
    .I0(__705__),
    .O(__2510__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5891__ (
    .I1(g35),
    .I0(__818__),
    .O(__2511__)
  );
  LUT3 #(
    .INIT(8'h01)
  ) __5892__ (
    .I2(__196__),
    .I1(__1028__),
    .I0(__1489__),
    .O(__2512__)
  );
  LUT5 #(
    .INIT(32'h33aaf0f0)
  ) __5893__ (
    .I4(g35),
    .I3(__2512__),
    .I2(__372__),
    .I1(__1980__),
    .I0(__800__),
    .O(__2513__)
  );
  LUT6 #(
    .INIT(64'hfefeff00ff00ff00)
  ) __5894__ (
    .I5(g35),
    .I4(__341__),
    .I3(__1213__),
    .I2(g72),
    .I1(g73),
    .I0(__824__),
    .O(__2514__)
  );
  LUT6 #(
    .INIT(64'hc0c0c0cd00000000)
  ) __5895__ (
    .I5(g35),
    .I4(__1111__),
    .I3(__1779__),
    .I2(__1782__),
    .I1(__860__),
    .I0(__908__),
    .O(__2515__)
  );
  LUT3 #(
    .INIT(8'h01)
  ) __5896__ (
    .I2(__357__),
    .I1(__613__),
    .I0(__623__),
    .O(__2516__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5897__ (
    .I5(g35),
    .I4(__1728__),
    .I3(__2516__),
    .I2(__135__),
    .I1(__27__),
    .I0(__1391__),
    .O(__2517__)
  );
  LUT4 #(
    .INIT(16'h0ef0)
  ) __5898__ (
    .I3(g35),
    .I2(__383__),
    .I1(__440__),
    .I0(__36__),
    .O(__2518__)
  );
  LUT6 #(
    .INIT(64'hb3bb8088aaaaaaaa)
  ) __5899__ (
    .I5(g35),
    .I4(__639__),
    .I3(__599__),
    .I2(__461__),
    .I1(__1586__),
    .I0(__596__),
    .O(__2519__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __5900__ (
    .I2(g35),
    .I1(__1147__),
    .I0(__768__),
    .O(__2520__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5901__ (
    .I1(__1154__),
    .I0(__1126__),
    .O(__2521__)
  );
  LUT6 #(
    .INIT(64'h0fffffffffff7777)
  ) __5902__ (
    .I5(__1154__),
    .I4(__1126__),
    .I3(__103__),
    .I2(__274__),
    .I1(__187__),
    .I0(__477__),
    .O(__2522__)
  );
  LUT6 #(
    .INIT(64'h7f00000000007f00)
  ) __5903__ (
    .I5(__62__),
    .I4(__823__),
    .I3(__2522__),
    .I2(__1199__),
    .I1(__853__),
    .I0(__2521__),
    .O(__2523__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5904__ (
    .I1(__1126__),
    .I0(__1154__),
    .O(__2524__)
  );
  LUT6 #(
    .INIT(64'hffff0fffffff7777)
  ) __5905__ (
    .I5(__1154__),
    .I4(__1126__),
    .I3(__404__),
    .I2(__187__),
    .I1(__686__),
    .I0(__1199__),
    .O(__2525__)
  );
  LUT6 #(
    .INIT(64'h00007f007f000000)
  ) __5906__ (
    .I5(__62__),
    .I4(__823__),
    .I3(__2525__),
    .I2(__1166__),
    .I1(__103__),
    .I0(__2524__),
    .O(__2526__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5907__ (
    .I1(__430__),
    .I0(__1135__),
    .O(__2527__)
  );
  LUT6 #(
    .INIT(64'h007f7f7f00000000)
  ) __5908__ (
    .I5(__62__),
    .I4(__2521__),
    .I3(__2527__),
    .I2(__1572__),
    .I1(__654__),
    .I0(__805__),
    .O(__2528__)
  );
  LUT6 #(
    .INIT(64'h000000f800000088)
  ) __5909__ (
    .I5(__1216__),
    .I4(__1154__),
    .I3(__1126__),
    .I2(__405__),
    .I1(__536__),
    .I0(__858__),
    .O(__2529__)
  );
  LUT6 #(
    .INIT(64'h000007770000ffff)
  ) __5910__ (
    .I5(__2524__),
    .I4(__2529__),
    .I3(__823__),
    .I2(__628__),
    .I1(__761__),
    .I0(__811__),
    .O(__2530__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __5911__ (
    .I1(__1154__),
    .I0(__1126__),
    .O(__2531__)
  );
  LUT6 #(
    .INIT(64'h0000f88800000000)
  ) __5912__ (
    .I5(__1154__),
    .I4(__1126__),
    .I3(__27__),
    .I2(__536__),
    .I1(__1216__),
    .I0(__51__),
    .O(__2532__)
  );
  LUT6 #(
    .INIT(64'h0000f88800000000)
  ) __5913__ (
    .I5(__1126__),
    .I4(__1154__),
    .I3(__833__),
    .I2(__202__),
    .I1(__162__),
    .I0(__654__),
    .O(__2533__)
  );
  LUT6 #(
    .INIT(64'h000007770000ffff)
  ) __5914__ (
    .I5(__1572__),
    .I4(__2533__),
    .I3(__156__),
    .I2(__811__),
    .I1(__823__),
    .I0(__135__),
    .O(__2534__)
  );
  LUT6 #(
    .INIT(64'h0000007f00000000)
  ) __5915__ (
    .I5(__2534__),
    .I4(__62__),
    .I3(__2532__),
    .I2(__1218__),
    .I1(__2531__),
    .I0(__1135__),
    .O(__2535__)
  );
  LUT3 #(
    .INIT(8'h07)
  ) __5916__ (
    .I2(__2535__),
    .I1(__2530__),
    .I0(__2528__),
    .O(__2536__)
  );
  LUT6 #(
    .INIT(64'hfffff11100000000)
  ) __5917__ (
    .I5(__2301__),
    .I4(__2536__),
    .I3(__2465__),
    .I2(__1278__),
    .I1(__2526__),
    .I0(__2523__),
    .O(__2537__)
  );
  LUT5 #(
    .INIT(32'hcf30aaaa)
  ) __5918__ (
    .I4(g35),
    .I3(__2537__),
    .I2(__960__),
    .I1(__2343__),
    .I0(__240__),
    .O(__2538__)
  );
  LUT6 #(
    .INIT(64'heaaa2aaaffff0000)
  ) __5919__ (
    .I5(g35),
    .I4(__630__),
    .I3(__457__),
    .I2(__874__),
    .I1(__1264__),
    .I0(__625__),
    .O(__2539__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5920__ (
    .I5(g35),
    .I4(__1852__),
    .I3(__1805__),
    .I2(__1075__),
    .I1(__748__),
    .I0(__1391__),
    .O(__2540__)
  );
  LUT5 #(
    .INIT(32'h00000008)
  ) __5921__ (
    .I4(__917__),
    .I3(__353__),
    .I2(__972__),
    .I1(__1444__),
    .I0(__1443__),
    .O(__2541__)
  );
  LUT5 #(
    .INIT(32'hffa0cfc0)
  ) __5922__ (
    .I4(__1643__),
    .I3(__958__),
    .I2(g35),
    .I1(__1208__),
    .I0(__2541__),
    .O(__2542__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5923__ (
    .I1(__874__),
    .I0(__1264__),
    .O(__2543__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5924__ (
    .I5(g35),
    .I4(__2543__),
    .I3(__2158__),
    .I2(__1120__),
    .I1(__165__),
    .I0(__1391__),
    .O(__2544__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5925__ (
    .I5(g35),
    .I4(__1692__),
    .I3(__2263__),
    .I2(__533__),
    .I1(__1132__),
    .I0(__1391__),
    .O(__2545__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5926__ (
    .I1(__267__),
    .I0(__425__),
    .O(__2546__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5927__ (
    .I5(g35),
    .I4(__2266__),
    .I3(__2546__),
    .I2(__57__),
    .I1(__444__),
    .I0(__1391__),
    .O(__2547__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5928__ (
    .I1(__1173__),
    .I0(__418__),
    .O(__2548__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5929__ (
    .I5(g35),
    .I4(__2548__),
    .I3(__1874__),
    .I2(__513__),
    .I1(__601__),
    .I0(__1391__),
    .O(__2549__)
  );
  LUT5 #(
    .INIT(32'h80000000)
  ) __5930__ (
    .I4(__217__),
    .I3(__395__),
    .I2(__1180__),
    .I1(__691__),
    .I0(__1438__),
    .O(__2550__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5931__ (
    .I1(__691__),
    .I0(__1180__),
    .O(__2551__)
  );
  LUT6 #(
    .INIT(64'h0fffffffffff7777)
  ) __5932__ (
    .I5(__1180__),
    .I4(__691__),
    .I3(__635__),
    .I2(__138__),
    .I1(__56__),
    .I0(__593__),
    .O(__2552__)
  );
  LUT6 #(
    .INIT(64'h7f00000000007f00)
  ) __5933__ (
    .I5(__395__),
    .I4(__1276__),
    .I3(__2552__),
    .I2(__2551__),
    .I1(__30__),
    .I0(__488__),
    .O(__2553__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5934__ (
    .I1(__1180__),
    .I0(__691__),
    .O(__2554__)
  );
  LUT6 #(
    .INIT(64'hffff0fffffff7777)
  ) __5935__ (
    .I5(__691__),
    .I4(__1180__),
    .I3(__1056__),
    .I2(__56__),
    .I1(__165__),
    .I0(__30__),
    .O(__2555__)
  );
  LUT6 #(
    .INIT(64'h00007f007f000000)
  ) __5936__ (
    .I5(__395__),
    .I4(__1276__),
    .I3(__2555__),
    .I2(__2554__),
    .I1(__1120__),
    .I0(__635__),
    .O(__2556__)
  );
  LUT4 #(
    .INIT(16'h8000)
  ) __5937__ (
    .I3(__217__),
    .I2(__395__),
    .I1(__1180__),
    .I0(__691__),
    .O(__2557__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5938__ (
    .I1(__520__),
    .I0(__326__),
    .O(__2558__)
  );
  LUT6 #(
    .INIT(64'h007f7f7f00000000)
  ) __5939__ (
    .I5(__395__),
    .I4(__2551__),
    .I3(__2558__),
    .I2(__1576__),
    .I1(__1169__),
    .I0(__268__),
    .O(__2559__)
  );
  LUT6 #(
    .INIT(64'h000000f800000088)
  ) __5940__ (
    .I5(__573__),
    .I4(__1180__),
    .I3(__691__),
    .I2(__558__),
    .I1(__59__),
    .I0(__164__),
    .O(__2560__)
  );
  LUT6 #(
    .INIT(64'h000007770000ffff)
  ) __5941__ (
    .I5(__2554__),
    .I4(__2560__),
    .I3(__1276__),
    .I2(__827__),
    .I1(__450__),
    .I0(__879__),
    .O(__2561__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __5942__ (
    .I1(__1180__),
    .I0(__691__),
    .O(__2562__)
  );
  LUT6 #(
    .INIT(64'h0000f88800000000)
  ) __5943__ (
    .I5(__691__),
    .I4(__1180__),
    .I3(__573__),
    .I2(__1132__),
    .I1(__59__),
    .I0(__37__),
    .O(__2563__)
  );
  LUT6 #(
    .INIT(64'h0000f88800000000)
  ) __5944__ (
    .I5(__1180__),
    .I4(__691__),
    .I3(__217__),
    .I2(__715__),
    .I1(__1169__),
    .I0(__144__),
    .O(__2564__)
  );
  LUT6 #(
    .INIT(64'h000007770000ffff)
  ) __5945__ (
    .I5(__1576__),
    .I4(__2564__),
    .I3(__1276__),
    .I2(__172__),
    .I1(__450__),
    .I0(__533__),
    .O(__2565__)
  );
  LUT6 #(
    .INIT(64'h0000007f00000000)
  ) __5946__ (
    .I5(__2565__),
    .I4(__395__),
    .I3(__2563__),
    .I2(__2562__),
    .I1(__948__),
    .I0(__520__),
    .O(__2566__)
  );
  LUT3 #(
    .INIT(8'h07)
  ) __5947__ (
    .I2(__2566__),
    .I1(__2561__),
    .I0(__2559__),
    .O(__2567__)
  );
  LUT6 #(
    .INIT(64'hfffff11100000000)
  ) __5948__ (
    .I5(__1438__),
    .I4(__2567__),
    .I3(__2557__),
    .I2(__1219__),
    .I1(__2556__),
    .I0(__2553__),
    .O(__2568__)
  );
  LUT5 #(
    .INIT(32'hcf30aaaa)
  ) __5949__ (
    .I4(g35),
    .I3(__2568__),
    .I2(__902__),
    .I1(__2550__),
    .I0(__1020__),
    .O(__2569__)
  );
  LUT6 #(
    .INIT(64'hcf03cf03cf038b8b)
  ) __5950__ (
    .I5(g113),
    .I4(__1283__),
    .I3(__607__),
    .I2(__821__),
    .I1(__1750__),
    .I0(__999__),
    .O(__2570__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __5951__ (
    .I2(g35),
    .I1(__2570__),
    .I0(__101__),
    .O(__2571__)
  );
  LUT6 #(
    .INIT(64'h6c206c6cf0f0f0f0)
  ) __5952__ (
    .I5(g35),
    .I4(__973__),
    .I3(__279__),
    .I2(__252__),
    .I1(__790__),
    .I0(__1818__),
    .O(__2572__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5953__ (
    .I5(g35),
    .I4(__2158__),
    .I3(__1761__),
    .I2(__138__),
    .I1(__488__),
    .I0(__1391__),
    .O(__2573__)
  );
  LUT5 #(
    .INIT(32'hccaa0f0f)
  ) __5954__ (
    .I4(__2019__),
    .I3(__1503__),
    .I2(__1158__),
    .I1(__999__),
    .I0(__1101__),
    .O(__2574__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __5955__ (
    .I2(g35),
    .I1(__2574__),
    .I0(__821__),
    .O(__2575__)
  );
  LUT6 #(
    .INIT(64'h3fc0ff00aaaaaaaa)
  ) __5956__ (
    .I5(g35),
    .I4(__784__),
    .I3(__743__),
    .I2(__462__),
    .I1(__1446__),
    .I0(__322__),
    .O(__2576__)
  );
  LUT6 #(
    .INIT(64'hff00df10ffff0000)
  ) __5957__ (
    .I5(g35),
    .I4(__962__),
    .I3(__1053__),
    .I2(__1393__),
    .I1(__1034__),
    .I0(__1391__),
    .O(__2577__)
  );
  LUT4 #(
    .INIT(16'h7f00)
  ) __5958__ (
    .I3(__261__),
    .I2(g35),
    .I1(__897__),
    .I0(__2040__),
    .O(__2578__)
  );
  LUT6 #(
    .INIT(64'h00005af0aaaaaaaa)
  ) __5959__ (
    .I5(g35),
    .I4(__1441__),
    .I3(__151__),
    .I2(__926__),
    .I1(__995__),
    .I0(__1192__),
    .O(__2579__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __5960__ (
    .I2(g35),
    .I1(__847__),
    .I0(__959__),
    .O(__2580__)
  );
  LUT6 #(
    .INIT(64'h0fff7f0070ff0000)
  ) __5961__ (
    .I5(__46__),
    .I4(__1211__),
    .I3(g35),
    .I2(__1678__),
    .I1(__1338__),
    .I0(__1677__),
    .O(__2581__)
  );
  LUT6 #(
    .INIT(64'hefffffff00000000)
  ) __5962__ (
    .I5(g35),
    .I4(__1110__),
    .I3(__762__),
    .I2(__1251__),
    .I1(__1043__),
    .I0(__1476__),
    .O(__2582__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __5963__ (
    .I2(__2582__),
    .I1(__579__),
    .I0(__77__),
    .O(__2583__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5964__ (
    .I1(__540__),
    .I0(__112__),
    .O(__2584__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5965__ (
    .I1(__23__),
    .I0(__142__),
    .O(__2585__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __5966__ (
    .I5(g35),
    .I4(__1430__),
    .I3(__2585__),
    .I2(__1080__),
    .I1(__8__),
    .I0(__2584__),
    .O(__2586__)
  );
  LUT5 #(
    .INIT(32'h80000000)
  ) __5967__ (
    .I4(__1004__),
    .I3(__1147__),
    .I2(__637__),
    .I1(__914__),
    .I0(__342__),
    .O(__2587__)
  );
  LUT5 #(
    .INIT(32'h0af0cccc)
  ) __5968__ (
    .I4(g35),
    .I3(__564__),
    .I2(__2587__),
    .I1(__637__),
    .I0(__1147__),
    .O(__2588__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5969__ (
    .I1(g35),
    .I0(__561__),
    .O(__2589__)
  );
  LUT3 #(
    .INIT(8'h04)
  ) __5970__ (
    .I2(__1538__),
    .I1(g35),
    .I0(__1535__),
    .O(__2590__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __5971__ (
    .I2(__1126__),
    .I1(__1261__),
    .I0(__1044__),
    .O(__2591__)
  );
  LUT5 #(
    .INIT(32'h00000008)
  ) __5972__ (
    .I4(__282__),
    .I3(__132__),
    .I2(__452__),
    .I1(__32__),
    .I0(__347__),
    .O(__2592__)
  );
  LUT6 #(
    .INIT(64'hebaa00aa00000000)
  ) __5973__ (
    .I5(g35),
    .I4(__2592__),
    .I3(__2301__),
    .I2(__1154__),
    .I1(__2591__),
    .I0(__906__),
    .O(__2593__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __5974__ (
    .I1(__833__),
    .I0(__1216__),
    .O(__2594__)
  );
  LUT6 #(
    .INIT(64'h0a03000000000000)
  ) __5975__ (
    .I5(g35),
    .I4(__2594__),
    .I3(__1199__),
    .I2(__187__),
    .I1(__103__),
    .I0(__823__),
    .O(__2595__)
  );
  LUT6 #(
    .INIT(64'hefefff00ff00ff00)
  ) __5976__ (
    .I5(g35),
    .I4(__341__),
    .I3(__266__),
    .I2(g72),
    .I1(g73),
    .I0(__1280__),
    .O(__2596__)
  );
  LUT6 #(
    .INIT(64'hfffc0003aaaaaaaa)
  ) __5977__ (
    .I5(g35),
    .I4(__969__),
    .I3(__728__),
    .I2(__1348__),
    .I1(__801__),
    .I0(__602__),
    .O(__2597__)
  );
  LUT6 #(
    .INIT(64'haaaaaaaccccccccc)
  ) __5978__ (
    .I5(g35),
    .I4(__595__),
    .I3(__112__),
    .I2(__1521__),
    .I1(__491__),
    .I0(__17__),
    .O(__2598__)
  );
  LUT6 #(
    .INIT(64'hcfcccfcc4544cfcc)
  ) __5979__ (
    .I5(__972__),
    .I4(__1444__),
    .I3(__1208__),
    .I2(__958__),
    .I1(__191__),
    .I0(__1953__),
    .O(__2599__)
  );
  LUT5 #(
    .INIT(32'h33aaf0f0)
  ) __5980__ (
    .I4(g35),
    .I3(__1643__),
    .I2(__41__),
    .I1(__2599__),
    .I0(__958__),
    .O(__2600__)
  );
  LUT5 #(
    .INIT(32'h00000008)
  ) __5981__ (
    .I4(g113),
    .I3(__1283__),
    .I2(__779__),
    .I1(__1060__),
    .I0(__1411__),
    .O(__2601__)
  );
  LUT5 #(
    .INIT(32'haaf030f0)
  ) __5982__ (
    .I4(__1555__),
    .I3(g35),
    .I2(__352__),
    .I1(__2601__),
    .I0(__746__),
    .O(__2602__)
  );
  LUT5 #(
    .INIT(32'h00cef0f0)
  ) __5983__ (
    .I4(g35),
    .I3(__74__),
    .I2(__464__),
    .I1(__227__),
    .I0(__193__),
    .O(__2603__)
  );
  LUT5 #(
    .INIT(32'hccaa0f0f)
  ) __5984__ (
    .I4(__2257__),
    .I3(__1503__),
    .I2(__9__),
    .I1(__999__),
    .I0(__933__),
    .O(__2604__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __5985__ (
    .I2(g35),
    .I1(__2604__),
    .I0(__1158__),
    .O(__2605__)
  );
  LUT4 #(
    .INIT(16'heef0)
  ) __5986__ (
    .I3(g35),
    .I2(__772__),
    .I1(__1273__),
    .I0(__755__),
    .O(__2606__)
  );
  LUT6 #(
    .INIT(64'hff00df10ffff0000)
  ) __5987__ (
    .I5(g35),
    .I4(__253__),
    .I3(__405__),
    .I2(__2516__),
    .I1(__689__),
    .I0(__1391__),
    .O(__2607__)
  );
  LUT5 #(
    .INIT(32'h143ccccc)
  ) __5988__ (
    .I4(g35),
    .I3(__1696__),
    .I2(__203__),
    .I1(__706__),
    .I0(__1396__),
    .O(__2608__)
  );
  LUT6 #(
    .INIT(64'h7f33b3b3cc000000)
  ) __5989__ (
    .I5(__211__),
    .I4(__687__),
    .I3(__214__),
    .I2(__197__),
    .I1(g35),
    .I0(__2351__),
    .O(__2609__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __5990__ (
    .I2(__1766__),
    .I1(__783__),
    .I0(__97__),
    .O(__2610__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5991__ (
    .I1(__1114__),
    .I0(__964__),
    .O(__2611__)
  );
  LUT6 #(
    .INIT(64'h3caaaaaaf0f0f0f0)
  ) __5992__ (
    .I5(g35),
    .I4(__1383__),
    .I3(__2611__),
    .I2(__1016__),
    .I1(__225__),
    .I0(__844__),
    .O(__2612__)
  );
  LUT3 #(
    .INIT(8'h08)
  ) __5993__ (
    .I2(__794__),
    .I1(g35),
    .I0(__1432__),
    .O(__2613__)
  );
  LUT6 #(
    .INIT(64'h000100ff00000000)
  ) __5994__ (
    .I5(__1423__),
    .I4(g35),
    .I3(__1421__),
    .I2(__20__),
    .I1(__750__),
    .I0(__1265__),
    .O(__2614__)
  );
  LUT4 #(
    .INIT(16'hbbf0)
  ) __5995__ (
    .I3(g35),
    .I2(__1061__),
    .I1(__2614__),
    .I0(__429__),
    .O(__2615__)
  );
  LUT3 #(
    .INIT(8'h2c)
  ) __5996__ (
    .I2(__396__),
    .I1(__544__),
    .I0(__646__),
    .O(__2616__)
  );
  LUT5 #(
    .INIT(32'h5df080f0)
  ) __5997__ (
    .I4(__594__),
    .I3(g35),
    .I2(__331__),
    .I1(__1207__),
    .I0(__2616__),
    .O(__2617__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __5998__ (
    .I2(g35),
    .I1(__415__),
    .I0(__104__),
    .O(__2618__)
  );
  LUT6 #(
    .INIT(64'h3bcc3bcc00000000)
  ) __5999__ (
    .I5(g35),
    .I4(__881__),
    .I3(__660__),
    .I2(__1115__),
    .I1(__170__),
    .I0(__1401__),
    .O(__2619__)
  );
  LUT5 #(
    .INIT(32'h80000000)
  ) __6000__ (
    .I4(__1063__),
    .I3(__376__),
    .I2(__527__),
    .I1(__254__),
    .I0(__1630__),
    .O(__2620__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __6001__ (
    .I1(__527__),
    .I0(__254__),
    .O(__2621__)
  );
  LUT6 #(
    .INIT(64'h0fffffffffff7777)
  ) __6002__ (
    .I5(__527__),
    .I4(__254__),
    .I3(__1074__),
    .I2(__531__),
    .I1(__1123__),
    .I0(__89__),
    .O(__2622__)
  );
  LUT6 #(
    .INIT(64'h7f00000000007f00)
  ) __6003__ (
    .I5(__376__),
    .I4(__1040__),
    .I3(__2622__),
    .I2(__286__),
    .I1(__351__),
    .I0(__2621__),
    .O(__2623__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __6004__ (
    .I1(__254__),
    .I0(__527__),
    .O(__2624__)
  );
  LUT6 #(
    .INIT(64'hffff0fffffff7777)
  ) __6005__ (
    .I5(__527__),
    .I4(__254__),
    .I3(__1123__),
    .I2(__797__),
    .I1(__351__),
    .I0(__703__),
    .O(__2625__)
  );
  LUT6 #(
    .INIT(64'h00007f007f000000)
  ) __6006__ (
    .I5(__376__),
    .I4(__1040__),
    .I3(__2625__),
    .I2(__1074__),
    .I1(__2624__),
    .I0(__856__),
    .O(__2626__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6007__ (
    .I1(__887__),
    .I0(__67__),
    .O(__2627__)
  );
  LUT6 #(
    .INIT(64'h007f7f7f00000000)
  ) __6008__ (
    .I5(__376__),
    .I4(__2621__),
    .I3(__2627__),
    .I2(__1570__),
    .I1(__72__),
    .I0(__852__),
    .O(__2628__)
  );
  LUT6 #(
    .INIT(64'h000000f800000088)
  ) __6009__ (
    .I5(__684__),
    .I4(__527__),
    .I3(__254__),
    .I2(__1053__),
    .I1(__920__),
    .I0(__634__),
    .O(__2629__)
  );
  LUT6 #(
    .INIT(64'h000007770000ffff)
  ) __6010__ (
    .I5(__2624__),
    .I4(__2629__),
    .I3(__929__),
    .I2(__1040__),
    .I1(__150__),
    .I0(__263__),
    .O(__2630__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __6011__ (
    .I1(__527__),
    .I0(__254__),
    .O(__2631__)
  );
  LUT6 #(
    .INIT(64'h0000f88800000000)
  ) __6012__ (
    .I5(__527__),
    .I4(__254__),
    .I3(__684__),
    .I2(__574__),
    .I1(__920__),
    .I0(__921__),
    .O(__2632__)
  );
  LUT6 #(
    .INIT(64'h0000f88800000000)
  ) __6013__ (
    .I5(__254__),
    .I4(__527__),
    .I3(__1063__),
    .I2(__1054__),
    .I1(__72__),
    .I0(__86__),
    .O(__2633__)
  );
  LUT6 #(
    .INIT(64'h000007770000ffff)
  ) __6014__ (
    .I5(__1570__),
    .I4(__2633__),
    .I3(__1040__),
    .I2(__1049__),
    .I1(__263__),
    .I0(__1163__),
    .O(__2634__)
  );
  LUT6 #(
    .INIT(64'h0000007f00000000)
  ) __6015__ (
    .I5(__2634__),
    .I4(__376__),
    .I3(__2632__),
    .I2(__2631__),
    .I1(__1007__),
    .I0(__887__),
    .O(__2635__)
  );
  LUT3 #(
    .INIT(8'h07)
  ) __6016__ (
    .I2(__2635__),
    .I1(__2630__),
    .I0(__2628__),
    .O(__2636__)
  );
  LUT6 #(
    .INIT(64'hfffff11100000000)
  ) __6017__ (
    .I5(__1630__),
    .I4(__2636__),
    .I3(__1847__),
    .I2(__1212__),
    .I1(__2626__),
    .I0(__2623__),
    .O(__2637__)
  );
  LUT5 #(
    .INIT(32'hcf30aaaa)
  ) __6018__ (
    .I4(g35),
    .I3(__2637__),
    .I2(__656__),
    .I1(__2620__),
    .I0(__951__),
    .O(__2638__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6019__ (
    .I5(g35),
    .I4(__2382__),
    .I3(__1793__),
    .I2(__807__),
    .I1(__234__),
    .I0(__1391__),
    .O(__2639__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6020__ (
    .I2(g35),
    .I1(__493__),
    .I0(__895__),
    .O(__2640__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __6021__ (
    .I1(__352__),
    .I0(__1555__),
    .O(__2641__)
  );
  LUT6 #(
    .INIT(64'hf055f0f0cccccccc)
  ) __6022__ (
    .I5(g35),
    .I4(__2641__),
    .I3(__793__),
    .I2(__402__),
    .I1(__1241__),
    .I0(__1552__),
    .O(__2642__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __6023__ (
    .I1(__1111__),
    .I0(__1782__),
    .O(__2643__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6024__ (
    .I5(g35),
    .I4(__860__),
    .I3(__2643__),
    .I2(__233__),
    .I1(__690__),
    .I0(__2034__),
    .O(__2644__)
  );
  LUT6 #(
    .INIT(64'hfefeff00ff00ff00)
  ) __6025__ (
    .I5(g35),
    .I4(__341__),
    .I3(__553__),
    .I2(g72),
    .I1(g73),
    .I0(__390__),
    .O(__2645__)
  );
  LUT6 #(
    .INIT(64'haaaaaaaccccccccc)
  ) __6026__ (
    .I5(g35),
    .I4(__1269__),
    .I3(__1638__),
    .I2(__318__),
    .I1(__355__),
    .I0(__978__),
    .O(__2646__)
  );
  LUT6 #(
    .INIT(64'h000000000000bf00)
  ) __6027__ (
    .I5(__425__),
    .I4(__157__),
    .I3(g35),
    .I2(__1773__),
    .I1(__1303__),
    .I0(__810__),
    .O(__2647__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6028__ (
    .I5(g35),
    .I4(__2546__),
    .I3(__1790__),
    .I2(__420__),
    .I1(__324__),
    .I0(__1391__),
    .O(__2648__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6029__ (
    .I5(g35),
    .I4(__1946__),
    .I3(__2516__),
    .I2(__628__),
    .I1(__858__),
    .I0(__1391__),
    .O(__2649__)
  );
  LUT3 #(
    .INIT(8'h35)
  ) __6030__ (
    .I2(__1142__),
    .I1(__384__),
    .I0(__448__),
    .O(__2650__)
  );
  LUT5 #(
    .INIT(32'h4040ff00)
  ) __6031__ (
    .I4(g35),
    .I3(__218__),
    .I2(__1033__),
    .I1(__2650__),
    .I0(__303__),
    .O(__2651__)
  );
  LUT6 #(
    .INIT(64'haaaaaaaccccccccc)
  ) __6032__ (
    .I5(g35),
    .I4(__746__),
    .I3(__793__),
    .I2(__1555__),
    .I1(__855__),
    .I0(__332__),
    .O(__2652__)
  );
  LUT5 #(
    .INIT(32'h7fff0000)
  ) __6033__ (
    .I4(__678__),
    .I3(g35),
    .I2(__1503__),
    .I1(__1440__),
    .I0(__15__),
    .O(__2653__)
  );
  LUT5 #(
    .INIT(32'hbf80aaaa)
  ) __6034__ (
    .I4(g35),
    .I3(__765__),
    .I2(__1896__),
    .I1(__1904__),
    .I0(__1232__),
    .O(__2654__)
  );
  LUT5 #(
    .INIT(32'hccaaf0f0)
  ) __6035__ (
    .I4(g35),
    .I3(__1864__),
    .I2(__439__),
    .I1(__994__),
    .I0(__22__),
    .O(__2655__)
  );
  LUT6 #(
    .INIT(64'h4444f0f0ff00ff00)
  ) __6036__ (
    .I5(g35),
    .I4(__1451__),
    .I3(__184__),
    .I2(__949__),
    .I1(__480__),
    .I0(__758__),
    .O(__2656__)
  );
  LUT6 #(
    .INIT(64'hefefff00ff00ff00)
  ) __6037__ (
    .I5(g35),
    .I4(__341__),
    .I3(__919__),
    .I2(g73),
    .I1(g72),
    .I0(__25__),
    .O(__2657__)
  );
  LUT5 #(
    .INIT(32'haaf030f0)
  ) __6038__ (
    .I4(__1521__),
    .I3(g35),
    .I2(__540__),
    .I1(__1523__),
    .I0(__595__),
    .O(__2658__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __6039__ (
    .I1(__190__),
    .I0(__1028__),
    .O(__2659__)
  );
  LUT6 #(
    .INIT(64'hf055f0f0cccccccc)
  ) __6040__ (
    .I5(g35),
    .I4(__2659__),
    .I3(__1489__),
    .I2(__922__),
    .I1(__411__),
    .I0(__1980__),
    .O(__2660__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6041__ (
    .I1(__506__),
    .I0(__934__),
    .O(__2661__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __6042__ (
    .I1(__78__),
    .I0(__934__),
    .O(__2662__)
  );
  LUT6 #(
    .INIT(64'hffccff00f0f0fafa)
  ) __6043__ (
    .I5(__653__),
    .I4(__1237__),
    .I3(__2662__),
    .I2(__2661__),
    .I1(__1131__),
    .I0(__675__),
    .O(__2663__)
  );
  LUT5 #(
    .INIT(32'h0f05030f)
  ) __6044__ (
    .I4(__1237__),
    .I3(__934__),
    .I2(__2663__),
    .I1(__1023__),
    .I0(__763__),
    .O(__2664__)
  );
  LUT5 #(
    .INIT(32'h33aaf0f0)
  ) __6045__ (
    .I4(g35),
    .I3(__1708__),
    .I2(__1237__),
    .I1(__2664__),
    .I0(__1048__),
    .O(__2665__)
  );
  LUT4 #(
    .INIT(16'h3caa)
  ) __6046__ (
    .I3(g35),
    .I2(__2550__),
    .I1(__630__),
    .I0(__201__),
    .O(__2666__)
  );
  LUT4 #(
    .INIT(16'h1f30)
  ) __6047__ (
    .I3(__1187__),
    .I2(g35),
    .I1(__31__),
    .I0(__1885__),
    .O(__2667__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6048__ (
    .I5(g35),
    .I4(__2450__),
    .I3(__1632__),
    .I2(__909__),
    .I1(__826__),
    .I0(__1391__),
    .O(__2668__)
  );
  LUT6 #(
    .INIT(64'h03300ff0aaaaaaaa)
  ) __6049__ (
    .I5(g35),
    .I4(__1696__),
    .I3(__1698__),
    .I2(__32__),
    .I1(__1396__),
    .I0(__1069__),
    .O(__2669__)
  );
  LUT6 #(
    .INIT(64'h7fd55555aa000000)
  ) __6050__ (
    .I5(__810__),
    .I4(__752__),
    .I3(__757__),
    .I2(__445__),
    .I1(__2005__),
    .I0(g35),
    .O(__2670__)
  );
  LUT5 #(
    .INIT(32'h00cef0f0)
  ) __6051__ (
    .I4(g35),
    .I3(__1270__),
    .I2(__848__),
    .I1(__1167__),
    .I0(__624__),
    .O(__2671__)
  );
  LUT5 #(
    .INIT(32'h7d55a000)
  ) __6052__ (
    .I4(__795__),
    .I3(__650__),
    .I2(__465__),
    .I1(__718__),
    .I0(g35),
    .O(__2672__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6053__ (
    .I2(g35),
    .I1(__297__),
    .I0(__1057__),
    .O(__2673__)
  );
  LUT6 #(
    .INIT(64'hb3bb8088aaaaaaaa)
  ) __6054__ (
    .I5(g35),
    .I4(__596__),
    .I3(__599__),
    .I2(__461__),
    .I1(__1586__),
    .I0(__779__),
    .O(__2674__)
  );
  LUT6 #(
    .INIT(64'heaaa2aaaffff0000)
  ) __6055__ (
    .I5(g35),
    .I4(__110__),
    .I3(__457__),
    .I2(__874__),
    .I1(__1264__),
    .I0(__1020__),
    .O(__2675__)
  );
  LUT6 #(
    .INIT(64'h7f5f8f0ff0500000)
  ) __6056__ (
    .I5(__289__),
    .I4(__116__),
    .I3(__1832__),
    .I2(g35),
    .I1(__413__),
    .I0(__2172__),
    .O(__2676__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6057__ (
    .I1(g35),
    .I0(__874__),
    .O(__2677__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __6058__ (
    .I1(__760__),
    .I0(__541__),
    .O(__2678__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6059__ (
    .I5(g35),
    .I4(__1299__),
    .I3(__2678__),
    .I2(__453__),
    .I1(__1050__),
    .I0(__2659__),
    .O(__2679__)
  );
  LUT6 #(
    .INIT(64'h5adaaa2affff0000)
  ) __6060__ (
    .I5(g35),
    .I4(__552__),
    .I3(__769__),
    .I2(__1286__),
    .I1(__819__),
    .I0(__1194__),
    .O(__2680__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6061__ (
    .I5(g35),
    .I4(__1712__),
    .I3(__1805__),
    .I2(__568__),
    .I1(__1259__),
    .I0(__1391__),
    .O(__2681__)
  );
  LUT5 #(
    .INIT(32'h7d55a000)
  ) __6062__ (
    .I4(__1190__),
    .I3(__752__),
    .I2(__1224__),
    .I1(__614__),
    .I0(g35),
    .O(__2682__)
  );
  LUT6 #(
    .INIT(64'h0000000000008000)
  ) __6063__ (
    .I5(__917__),
    .I4(__353__),
    .I3(__972__),
    .I2(__1503__),
    .I1(__1443__),
    .I0(__1708__),
    .O(__2683__)
  );
  LUT6 #(
    .INIT(64'hf30caaaaf0f0f0f0)
  ) __6064__ (
    .I5(g35),
    .I4(__2683__),
    .I3(__749__),
    .I2(__934__),
    .I1(__1237__),
    .I0(__174__),
    .O(__2684__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6065__ (
    .I5(g35),
    .I4(__2046__),
    .I3(__2382__),
    .I2(__1064__),
    .I1(__1191__),
    .I0(__1391__),
    .O(__2685__)
  );
  LUT3 #(
    .INIT(8'he0)
  ) __6066__ (
    .I2(__1041__),
    .I1(__1207__),
    .I0(__936__),
    .O(__2686__)
  );
  LUT6 #(
    .INIT(64'hefffefffffff0000)
  ) __6067__ (
    .I5(g35),
    .I4(__40__),
    .I3(__1115__),
    .I2(__2686__),
    .I1(__1399__),
    .I0(__345__),
    .O(__2687__)
  );
  LUT6 #(
    .INIT(64'h3f3f002affff00aa)
  ) __6068__ (
    .I5(__972__),
    .I4(__13__),
    .I3(__711__),
    .I2(__1444__),
    .I1(__1298__),
    .I0(__91__),
    .O(__2688__)
  );
  LUT5 #(
    .INIT(32'h33aaf0f0)
  ) __6069__ (
    .I4(g35),
    .I3(__1718__),
    .I2(__737__),
    .I1(__2688__),
    .I0(__711__),
    .O(__2689__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6070__ (
    .I1(__798__),
    .I0(__386__),
    .O(__2690__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6071__ (
    .I5(g35),
    .I4(__2690__),
    .I3(__1715__),
    .I2(__797__),
    .I1(__856__),
    .I0(__1391__),
    .O(__2691__)
  );
  LUT5 #(
    .INIT(32'h40ff0000)
  ) __6072__ (
    .I4(__582__),
    .I3(g35),
    .I2(__482__),
    .I1(__1432__),
    .I0(__794__),
    .O(__2692__)
  );
  LUT5 #(
    .INIT(32'h10ff0000)
  ) __6073__ (
    .I4(g35),
    .I3(__2199__),
    .I2(__2196__),
    .I1(__151__),
    .I0(__2195__),
    .O(__2693__)
  );
  LUT5 #(
    .INIT(32'hf3ff8ccc)
  ) __6074__ (
    .I4(__269__),
    .I3(__321__),
    .I2(__1147__),
    .I1(g35),
    .I0(__776__),
    .O(__2694__)
  );
  LUT5 #(
    .INIT(32'h00000080)
  ) __6075__ (
    .I4(__132__),
    .I3(__452__),
    .I2(__282__),
    .I1(__32__),
    .I0(__347__),
    .O(__2695__)
  );
  LUT6 #(
    .INIT(64'hccccf0aaf0f0f0f0)
  ) __6076__ (
    .I5(g35),
    .I4(__1609__),
    .I3(__2695__),
    .I2(__679__),
    .I1(__515__),
    .I0(__125__),
    .O(__2696__)
  );
  LUT4 #(
    .INIT(16'h0080)
  ) __6077__ (
    .I3(__1240__),
    .I2(__1567__),
    .I1(__1052__),
    .I0(__1236__),
    .O(__2697__)
  );
  LUT6 #(
    .INIT(64'h0fff7f0070ff0000)
  ) __6078__ (
    .I5(__830__),
    .I4(__726__),
    .I3(g35),
    .I2(__2254__),
    .I1(__1338__),
    .I0(__2697__),
    .O(__2698__)
  );
  LUT5 #(
    .INIT(32'hefefff00)
  ) __6079__ (
    .I4(g35),
    .I3(__345__),
    .I2(g44),
    .I1(__388__),
    .I0(__478__),
    .O(__2699__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6080__ (
    .I1(g35),
    .I0(__892__),
    .O(__2700__)
  );
  LUT4 #(
    .INIT(16'h3caa)
  ) __6081__ (
    .I3(g35),
    .I2(__1110__),
    .I1(__762__),
    .I0(__1043__),
    .O(__2701__)
  );
  LUT6 #(
    .INIT(64'h5adaaa2affff0000)
  ) __6082__ (
    .I5(g35),
    .I4(__369__),
    .I3(__462__),
    .I2(__1446__),
    .I1(__469__),
    .I0(__108__),
    .O(__2702__)
  );
  LUT5 #(
    .INIT(32'hffa0cfc0)
  ) __6083__ (
    .I4(__1430__),
    .I3(__243__),
    .I2(g35),
    .I1(__23__),
    .I0(__1466__),
    .O(__2703__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __6084__ (
    .I1(__1028__),
    .I0(__1489__),
    .O(__2704__)
  );
  LUT6 #(
    .INIT(64'hf055f0f0cccccccc)
  ) __6085__ (
    .I5(g35),
    .I4(__2704__),
    .I3(__190__),
    .I2(__431__),
    .I1(__800__),
    .I0(__1980__),
    .O(__2705__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6086__ (
    .I1(__142__),
    .I0(__243__),
    .O(__2706__)
  );
  LUT6 #(
    .INIT(64'hc3aaaaaaf0f0f0f0)
  ) __6087__ (
    .I5(g35),
    .I4(__1430__),
    .I3(__2706__),
    .I2(__1231__),
    .I1(__1062__),
    .I0(__534__),
    .O(__2707__)
  );
  LUT4 #(
    .INIT(16'hefa0)
  ) __6088__ (
    .I3(__756__),
    .I2(g35),
    .I1(__2402__),
    .I0(__192__),
    .O(__2708__)
  );
  LUT6 #(
    .INIT(64'h06666666aaaaaaaa)
  ) __6089__ (
    .I5(g35),
    .I4(__1303__),
    .I3(__810__),
    .I2(__1302__),
    .I1(__900__),
    .I0(__412__),
    .O(__2709__)
  );
  LUT4 #(
    .INIT(16'h8f00)
  ) __6090__ (
    .I3(__1251__),
    .I2(g35),
    .I1(__1110__),
    .I0(__547__),
    .O(__2710__)
  );
  LUT6 #(
    .INIT(64'h0000ff000000efef)
  ) __6091__ (
    .I5(__1469__),
    .I4(__1473__),
    .I3(__804__),
    .I2(__1248__),
    .I1(__1342__),
    .I0(__1472__),
    .O(__2711__)
  );
  LUT6 #(
    .INIT(64'h6666666affff0000)
  ) __6092__ (
    .I5(g35),
    .I4(__645__),
    .I3(__950__),
    .I2(__1473__),
    .I1(__632__),
    .I0(__2711__),
    .O(__2712__)
  );
  LUT6 #(
    .INIT(64'hfffc0003aaaaaaaa)
  ) __6093__ (
    .I5(g35),
    .I4(__578__),
    .I3(__950__),
    .I2(__645__),
    .I1(__1473__),
    .I0(__1149__),
    .O(__2713__)
  );
  LUT6 #(
    .INIT(64'haaaaaaaccccccccc)
  ) __6094__ (
    .I5(g35),
    .I4(__746__),
    .I3(__793__),
    .I2(__1555__),
    .I1(__1230__),
    .I0(__82__),
    .O(__2714__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6095__ (
    .I1(__1208__),
    .I0(__589__),
    .O(__2715__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __6096__ (
    .I1(__834__),
    .I0(__1208__),
    .O(__2716__)
  );
  LUT6 #(
    .INIT(64'hffccff00f0f0fafa)
  ) __6097__ (
    .I5(__958__),
    .I4(__191__),
    .I3(__2716__),
    .I2(__2715__),
    .I1(__532__),
    .I0(__1059__),
    .O(__2717__)
  );
  LUT5 #(
    .INIT(32'h0f05030f)
  ) __6098__ (
    .I4(__191__),
    .I3(__1208__),
    .I2(__2717__),
    .I1(__828__),
    .I0(__63__),
    .O(__2718__)
  );
  LUT5 #(
    .INIT(32'h33aaf0f0)
  ) __6099__ (
    .I4(g35),
    .I3(__1643__),
    .I2(__191__),
    .I1(__2718__),
    .I0(__963__),
    .O(__2719__)
  );
  LUT3 #(
    .INIT(8'h78)
  ) __6100__ (
    .I2(__707__),
    .I1(g35),
    .I0(__117__),
    .O(__2720__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6101__ (
    .I2(g35),
    .I1(__638__),
    .I0(__888__),
    .O(__2721__)
  );
  LUT6 #(
    .INIT(64'haaaaaaaccccccccc)
  ) __6102__ (
    .I5(g35),
    .I4(__196__),
    .I3(__1028__),
    .I2(__1489__),
    .I1(__1002__),
    .I0(__372__),
    .O(__2722__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6103__ (
    .I2(g35),
    .I1(__104__),
    .I0(__494__),
    .O(__2723__)
  );
  LUT5 #(
    .INIT(32'h10ff0000)
  ) __6104__ (
    .I4(__832__),
    .I3(g35),
    .I2(__791__),
    .I1(__898__),
    .I0(__1835__),
    .O(__2724__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __6105__ (
    .I1(__950__),
    .I0(__1473__),
    .O(__2725__)
  );
  LUT6 #(
    .INIT(64'hf055f0f0cccccccc)
  ) __6106__ (
    .I5(g35),
    .I4(__2725__),
    .I3(__1014__),
    .I2(__589__),
    .I1(__532__),
    .I0(__1470__),
    .O(__2726__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6107__ (
    .I5(g35),
    .I4(__1866__),
    .I3(__1633__),
    .I2(__377__),
    .I1(__370__),
    .I0(__1391__),
    .O(__2727__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __6108__ (
    .I1(__1242__),
    .I0(g35),
    .O(__2728__)
  );
  LUT6 #(
    .INIT(64'h8000000000000000)
  ) __6109__ (
    .I5(__1043__),
    .I4(__1110__),
    .I3(__762__),
    .I2(__1251__),
    .I1(__265__),
    .I0(__695__),
    .O(__2729__)
  );
  LUT6 #(
    .INIT(64'h7fffd50055005500)
  ) __6110__ (
    .I5(__1549__),
    .I4(__1125__),
    .I3(__414__),
    .I2(__403__),
    .I1(__2729__),
    .I0(g35),
    .O(__2730__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6111__ (
    .I5(g35),
    .I4(__112__),
    .I3(__1828__),
    .I2(__8__),
    .I1(__608__),
    .I0(__1827__),
    .O(__2731__)
  );
  LUT5 #(
    .INIT(32'hffa0cfc0)
  ) __6112__ (
    .I4(__1718__),
    .I3(__711__),
    .I2(g35),
    .I1(__91__),
    .I0(__1717__),
    .O(__2732__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6113__ (
    .I5(g35),
    .I4(__306__),
    .I3(__1660__),
    .I2(__458__),
    .I1(__1185__),
    .I0(__1391__),
    .O(__2733__)
  );
  LUT5 #(
    .INIT(32'hd2dd0000)
  ) __6114__ (
    .I4(g35),
    .I3(__1248__),
    .I2(__1245__),
    .I1(__1528__),
    .I0(__1024__),
    .O(__2734__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6115__ (
    .I2(g35),
    .I1(__291__),
    .I0(__1035__),
    .O(__2735__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6116__ (
    .I1(__469__),
    .I0(__336__),
    .O(__2736__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __6117__ (
    .I1(__690__),
    .I0(__469__),
    .O(__2737__)
  );
  LUT6 #(
    .INIT(64'hffccff00f0f0fafa)
  ) __6118__ (
    .I5(__462__),
    .I4(__784__),
    .I3(__2737__),
    .I2(__2736__),
    .I1(__7__),
    .I0(__233__),
    .O(__2738__)
  );
  LUT5 #(
    .INIT(32'h0f05030f)
  ) __6119__ (
    .I4(__784__),
    .I3(__469__),
    .I2(__2738__),
    .I1(__111__),
    .I0(__1122__),
    .O(__2739__)
  );
  LUT5 #(
    .INIT(32'h33aaf0f0)
  ) __6120__ (
    .I4(g35),
    .I3(__1446__),
    .I2(__784__),
    .I1(__2739__),
    .I0(__369__),
    .O(__2740__)
  );
  LUT5 #(
    .INIT(32'h3caaf0f0)
  ) __6121__ (
    .I4(g35),
    .I3(__2620__),
    .I2(__656__),
    .I1(__951__),
    .I0(__298__),
    .O(__2741__)
  );
  LUT6 #(
    .INIT(64'hee22eeeef0f0f0f0)
  ) __6122__ (
    .I5(g35),
    .I4(__1248__),
    .I3(__1245__),
    .I2(__354__),
    .I1(__1584__),
    .I0(__173__),
    .O(__2742__)
  );
  LUT6 #(
    .INIT(64'heaaa2aaaffff0000)
  ) __6123__ (
    .I5(g35),
    .I4(__915__),
    .I3(__253__),
    .I2(__689__),
    .I1(__623__),
    .I0(__676__),
    .O(__2743__)
  );
  LUT6 #(
    .INIT(64'h0000000080000000)
  ) __6124__ (
    .I5(__596__),
    .I4(__639__),
    .I3(__163__),
    .I2(__2372__),
    .I1(__955__),
    .I0(__1203__),
    .O(__2744__)
  );
  LUT5 #(
    .INIT(32'h73bbc000)
  ) __6125__ (
    .I4(__641__),
    .I3(__277__),
    .I2(__2372__),
    .I1(g35),
    .I0(__2744__),
    .O(__2745__)
  );
  LUT5 #(
    .INIT(32'h08880808)
  ) __6126__ (
    .I4(__881__),
    .I3(__660__),
    .I2(__1115__),
    .I1(__170__),
    .I0(__1401__),
    .O(__2746__)
  );
  LUT5 #(
    .INIT(32'h575d0a00)
  ) __6127__ (
    .I4(__134__),
    .I3(__148__),
    .I2(__2746__),
    .I1(__1973__),
    .I0(g35),
    .O(__2747__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6128__ (
    .I5(g35),
    .I4(__1791__),
    .I3(__2266__),
    .I2(__444__),
    .I1(__95__),
    .I0(__1391__),
    .O(__2748__)
  );
  LUT6 #(
    .INIT(64'hf0f04444ff00ff00)
  ) __6129__ (
    .I5(g35),
    .I4(__1555__),
    .I3(__422__),
    .I2(__352__),
    .I1(__793__),
    .I0(__2601__),
    .O(__2749__)
  );
  LUT6 #(
    .INIT(64'hff3030bfffff0000)
  ) __6130__ (
    .I5(g35),
    .I4(__576__),
    .I3(__734__),
    .I2(__588__),
    .I1(__1003__),
    .I0(__1011__),
    .O(__2750__)
  );
  LUT6 #(
    .INIT(64'h557f55d500aa0000)
  ) __6131__ (
    .I5(__132__),
    .I4(__282__),
    .I3(__1697__),
    .I2(__347__),
    .I1(__1859__),
    .I0(g35),
    .O(__2751__)
  );
  LUT6 #(
    .INIT(64'h3fffc000aaaaaaaa)
  ) __6132__ (
    .I5(g35),
    .I4(__658__),
    .I3(__253__),
    .I2(__689__),
    .I1(__623__),
    .I0(__918__),
    .O(__2752__)
  );
  LUT6 #(
    .INIT(64'h5adaaa2affff0000)
  ) __6133__ (
    .I5(g35),
    .I4(__537__),
    .I3(__243__),
    .I2(__1430__),
    .I1(__23__),
    .I0(__373__),
    .O(__2753__)
  );
  LUT5 #(
    .INIT(32'haaf030f0)
  ) __6134__ (
    .I4(__1473__),
    .I3(g35),
    .I2(__1014__),
    .I1(__2215__),
    .I0(__645__),
    .O(__2754__)
  );
  LUT3 #(
    .INIT(8'h08)
  ) __6135__ (
    .I2(__507__),
    .I1(__1032__),
    .I0(__709__),
    .O(__2755__)
  );
  LUT6 #(
    .INIT(64'hdfff7555aaaa0000)
  ) __6136__ (
    .I5(__767__),
    .I4(__334__),
    .I3(__88__),
    .I2(__2755__),
    .I1(__835__),
    .I0(g35),
    .O(__2756__)
  );
  LUT5 #(
    .INIT(32'hc3aaf0f0)
  ) __6137__ (
    .I4(g35),
    .I3(__2459__),
    .I2(__360__),
    .I1(__1119__),
    .I0(__602__),
    .O(__2757__)
  );
  LUT4 #(
    .INIT(16'h0008)
  ) __6138__ (
    .I3(__1240__),
    .I2(__1052__),
    .I1(__1567__),
    .I0(__1236__),
    .O(__2758__)
  );
  LUT6 #(
    .INIT(64'h0077ff00f0f0f0f0)
  ) __6139__ (
    .I5(g35),
    .I4(__1673__),
    .I3(__511__),
    .I2(__31__),
    .I1(__1338__),
    .I0(__2758__),
    .O(__2759__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6140__ (
    .I5(g35),
    .I4(__1660__),
    .I3(__2363__),
    .I2(__1015__),
    .I1(__1214__),
    .I0(__1391__),
    .O(__2760__)
  );
  LUT4 #(
    .INIT(16'h3caa)
  ) __6141__ (
    .I3(g35),
    .I2(__2343__),
    .I1(__915__),
    .I0(__971__),
    .O(__2761__)
  );
  LUT5 #(
    .INIT(32'h01ff0000)
  ) __6142__ (
    .I4(g35),
    .I3(__473__),
    .I2(__1503__),
    .I1(g72),
    .I0(g73),
    .O(__2762__)
  );
  LUT6 #(
    .INIT(64'h7fffffff00000000)
  ) __6143__ (
    .I5(__2762__),
    .I4(__738__),
    .I3(__976__),
    .I2(__1775__),
    .I1(__871__),
    .I0(__301__),
    .O(__2763__)
  );
  LUT6 #(
    .INIT(64'h7fffd50055005500)
  ) __6144__ (
    .I5(__2763__),
    .I4(__92__),
    .I3(__114__),
    .I2(__343__),
    .I1(__1871__),
    .I0(g35),
    .O(__2764__)
  );
  LUT6 #(
    .INIT(64'h00007fff7fff7fff)
  ) __6145__ (
    .I5(__1696__),
    .I4(__1396__),
    .I3(__1235__),
    .I2(__203__),
    .I1(__153__),
    .I0(__706__),
    .O(__2765__)
  );
  LUT6 #(
    .INIT(64'h48888888ffff0000)
  ) __6146__ (
    .I5(g35),
    .I4(__1235__),
    .I3(__203__),
    .I2(__706__),
    .I1(__2765__),
    .I0(__447__),
    .O(__2766__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6147__ (
    .I5(g35),
    .I4(__989__),
    .I3(__1793__),
    .I2(__883__),
    .I1(__570__),
    .I0(__1391__),
    .O(__2767__)
  );
  LUT6 #(
    .INIT(64'h7fd55555aa000000)
  ) __6148__ (
    .I5(__719__),
    .I4(__214__),
    .I3(__1117__),
    .I2(__606__),
    .I1(__546__),
    .I0(g35),
    .O(__2768__)
  );
  LUT6 #(
    .INIT(64'hfffc0003aaaaaaaa)
  ) __6149__ (
    .I5(g35),
    .I4(__308__),
    .I3(__944__),
    .I2(__296__),
    .I1(__1600__),
    .I0(__183__),
    .O(__2769__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __6150__ (
    .I2(__1224__),
    .I1(__1190__),
    .I0(__614__),
    .O(__2770__)
  );
  LUT5 #(
    .INIT(32'h78ccffcc)
  ) __6151__ (
    .I4(__752__),
    .I3(g35),
    .I2(__445__),
    .I1(__519__),
    .I0(__2770__),
    .O(__2771__)
  );
  LUT6 #(
    .INIT(64'h22882c8cff00ff00)
  ) __6152__ (
    .I5(g35),
    .I4(__544__),
    .I3(__1036__),
    .I2(__646__),
    .I1(__775__),
    .I0(__1813__),
    .O(__2772__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __6153__ (
    .I1(__318__),
    .I0(__1638__),
    .O(__2773__)
  );
  LUT6 #(
    .INIT(64'hf055f0f0cccccccc)
  ) __6154__ (
    .I5(g35),
    .I4(__2773__),
    .I3(__617__),
    .I2(__307__),
    .I1(__839__),
    .I0(__1733__),
    .O(__2774__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6155__ (
    .I2(g35),
    .I1(__884__),
    .I0(__1220__),
    .O(__2775__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6156__ (
    .I1(g35),
    .I0(__1118__),
    .O(__2776__)
  );
  LUT6 #(
    .INIT(64'heaaa2aaaffff0000)
  ) __6157__ (
    .I5(g35),
    .I4(__1089__),
    .I3(__313__),
    .I2(__569__),
    .I1(__989__),
    .I0(__1256__),
    .O(__2777__)
  );
  LUT5 #(
    .INIT(32'hbfbfff00)
  ) __6158__ (
    .I4(g35),
    .I3(__694__),
    .I2(__99__),
    .I1(__1018__),
    .I0(__209__),
    .O(__2778__)
  );
  LUT6 #(
    .INIT(64'h4ccccccc00000000)
  ) __6159__ (
    .I5(__706__),
    .I4(__282__),
    .I3(__132__),
    .I2(__1672__),
    .I1(__2255__),
    .I0(__125__),
    .O(__2779__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __6160__ (
    .I1(__830__),
    .I0(__726__),
    .O(__2780__)
  );
  LUT6 #(
    .INIT(64'h0fffffffffff7777)
  ) __6161__ (
    .I5(__726__),
    .I4(__830__),
    .I3(__518__),
    .I2(__309__),
    .I1(__723__),
    .I0(__1176__),
    .O(__2781__)
  );
  LUT6 #(
    .INIT(64'h7f00000000007f00)
  ) __6162__ (
    .I5(__68__),
    .I4(__816__),
    .I3(__2781__),
    .I2(__901__),
    .I1(__522__),
    .I0(__2780__),
    .O(__2782__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __6163__ (
    .I1(__726__),
    .I0(__830__),
    .O(__2783__)
  );
  LUT6 #(
    .INIT(64'hffff0fffffff7777)
  ) __6164__ (
    .I5(__830__),
    .I4(__726__),
    .I3(__723__),
    .I2(__354__),
    .I1(__901__),
    .I0(__136__),
    .O(__2784__)
  );
  LUT6 #(
    .INIT(64'h00007f007f000000)
  ) __6165__ (
    .I5(__68__),
    .I4(__816__),
    .I3(__2784__),
    .I2(__518__),
    .I1(__212__),
    .I0(__2783__),
    .O(__2785__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6166__ (
    .I1(__726__),
    .I0(__830__),
    .O(__2786__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6167__ (
    .I1(__98__),
    .I0(__556__),
    .O(__2787__)
  );
  LUT6 #(
    .INIT(64'h007f7f7f00000000)
  ) __6168__ (
    .I5(__816__),
    .I4(__2780__),
    .I3(__2787__),
    .I2(__2786__),
    .I1(__312__),
    .I0(__1229__),
    .O(__2788__)
  );
  LUT6 #(
    .INIT(64'h000000f800000088)
  ) __6169__ (
    .I5(__1006__),
    .I4(__726__),
    .I3(__830__),
    .I2(__826__),
    .I1(__416__),
    .I0(__311__),
    .O(__2789__)
  );
  LUT6 #(
    .INIT(64'h000007770000ffff)
  ) __6170__ (
    .I5(__2783__),
    .I4(__2789__),
    .I3(__68__),
    .I2(__545__),
    .I1(__398__),
    .I0(__909__),
    .O(__2790__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __6171__ (
    .I1(__726__),
    .I0(__830__),
    .O(__2791__)
  );
  LUT6 #(
    .INIT(64'h0000f88800000000)
  ) __6172__ (
    .I5(__830__),
    .I4(__726__),
    .I3(__1006__),
    .I2(__677__),
    .I1(__416__),
    .I0(__194__),
    .O(__2792__)
  );
  LUT6 #(
    .INIT(64'h0000f88800000000)
  ) __6173__ (
    .I5(__726__),
    .I4(__830__),
    .I3(__644__),
    .I2(__699__),
    .I1(__1010__),
    .I0(__312__),
    .O(__2793__)
  );
  LUT6 #(
    .INIT(64'h000007770000ffff)
  ) __6174__ (
    .I5(__2786__),
    .I4(__2793__),
    .I3(__68__),
    .I2(__281__),
    .I1(__370__),
    .I0(__398__),
    .O(__2794__)
  );
  LUT6 #(
    .INIT(64'h0000007f00000000)
  ) __6175__ (
    .I5(__2794__),
    .I4(__816__),
    .I3(__2792__),
    .I2(__377__),
    .I1(__2791__),
    .I0(__98__),
    .O(__2795__)
  );
  LUT3 #(
    .INIT(8'h07)
  ) __6176__ (
    .I2(__2795__),
    .I1(__2790__),
    .I0(__2788__),
    .O(__2796__)
  );
  LUT6 #(
    .INIT(64'hfffff11100000000)
  ) __6177__ (
    .I5(__2254__),
    .I4(__2796__),
    .I3(__2255__),
    .I2(__173__),
    .I1(__2785__),
    .I0(__2782__),
    .O(__2797__)
  );
  LUT5 #(
    .INIT(32'hcf30aaaa)
  ) __6178__ (
    .I4(g35),
    .I3(__2797__),
    .I2(__609__),
    .I1(__2779__),
    .I0(__195__),
    .O(__2798__)
  );
  LUT6 #(
    .INIT(64'hf0f04444ff00ff00)
  ) __6179__ (
    .I5(g35),
    .I4(__1348__),
    .I3(__812__),
    .I2(__179__),
    .I1(__801__),
    .I0(__1983__),
    .O(__2799__)
  );
  LUT4 #(
    .INIT(16'he0ee)
  ) __6180__ (
    .I3(__1813__),
    .I2(__1036__),
    .I1(__544__),
    .I0(__646__),
    .O(__2800__)
  );
  LUT6 #(
    .INIT(64'h7f5f8f0ff0500000)
  ) __6181__ (
    .I5(__1105__),
    .I4(__766__),
    .I3(__1813__),
    .I2(g35),
    .I1(__775__),
    .I0(__2800__),
    .O(__2801__)
  );
  LUT4 #(
    .INIT(16'h7f8a)
  ) __6182__ (
    .I3(__718__),
    .I2(__650__),
    .I1(__795__),
    .I0(g35),
    .O(__2802__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6183__ (
    .I1(g35),
    .I0(__590__),
    .O(__2803__)
  );
  LUT6 #(
    .INIT(64'h23238c8cff00ff00)
  ) __6184__ (
    .I5(g35),
    .I4(__587__),
    .I3(__497__),
    .I2(__973__),
    .I1(__1816__),
    .I0(__279__),
    .O(__2804__)
  );
  LUT5 #(
    .INIT(32'h0af0cccc)
  ) __6185__ (
    .I4(g35),
    .I3(__285__),
    .I2(__2065__),
    .I1(__1117__),
    .I0(__214__),
    .O(__2805__)
  );
  LUT3 #(
    .INIT(8'h01)
  ) __6186__ (
    .I2(__832__),
    .I1(__791__),
    .I0(__898__),
    .O(__2806__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6187__ (
    .I5(g35),
    .I4(__2806__),
    .I3(__2451__),
    .I2(__281__),
    .I1(__194__),
    .I0(__1391__),
    .O(__2807__)
  );
  LUT6 #(
    .INIT(64'hefefff00ff00ff00)
  ) __6188__ (
    .I5(g35),
    .I4(__341__),
    .I3(__391__),
    .I2(g72),
    .I1(g73),
    .I0(__25__),
    .O(__2808__)
  );
  LUT6 #(
    .INIT(64'h3fffc000aaaaaaaa)
  ) __6189__ (
    .I5(g35),
    .I4(__454__),
    .I3(__769__),
    .I2(__1286__),
    .I1(__982__),
    .I0(__16__),
    .O(__2809__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6190__ (
    .I1(g35),
    .I0(__785__),
    .O(__2810__)
  );
  LUT5 #(
    .INIT(32'hffa0cfc0)
  ) __6191__ (
    .I4(__1708__),
    .I3(__653__),
    .I2(g35),
    .I1(__934__),
    .I0(__1707__),
    .O(__2811__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6192__ (
    .I2(g35),
    .I1(__1204__),
    .I0(__1273__),
    .O(__2812__)
  );
  LUT6 #(
    .INIT(64'h45aa45aaffff0000)
  ) __6193__ (
    .I5(g35),
    .I4(__407__),
    .I3(__716__),
    .I2(__751__),
    .I1(__869__),
    .I0(__2441__),
    .O(__2813__)
  );
  LUT6 #(
    .INIT(64'h06666666aaaaaaaa)
  ) __6194__ (
    .I5(g35),
    .I4(__1773__),
    .I3(__1303__),
    .I2(__810__),
    .I1(__704__),
    .I0(__898__),
    .O(__2814__)
  );
  LUT5 #(
    .INIT(32'h73bbc000)
  ) __6195__ (
    .I4(__592__),
    .I3(__890__),
    .I2(__1147__),
    .I1(g35),
    .I0(__1662__),
    .O(__2815__)
  );
  LUT5 #(
    .INIT(32'h7d55a000)
  ) __6196__ (
    .I4(__914__),
    .I3(__1147__),
    .I2(__1004__),
    .I1(__342__),
    .I0(g35),
    .O(__2816__)
  );
  LUT6 #(
    .INIT(64'h00ff33330f0f5555)
  ) __6197__ (
    .I5(__465__),
    .I4(__842__),
    .I3(__101__),
    .I2(__821__),
    .I1(__1158__),
    .I0(__9__),
    .O(__2817__)
  );
  LUT5 #(
    .INIT(32'hff44f0f0)
  ) __6198__ (
    .I4(g35),
    .I3(__2237__),
    .I2(__899__),
    .I1(__247__),
    .I0(__1673__),
    .O(__2818__)
  );
  LUT4 #(
    .INIT(16'heef0)
  ) __6199__ (
    .I3(g35),
    .I2(__224__),
    .I1(__620__),
    .I0(__338__),
    .O(__2819__)
  );
  LUT5 #(
    .INIT(32'hffe0ffff)
  ) __6200__ (
    .I4(g35),
    .I3(__2350__),
    .I2(__1041__),
    .I1(__1207__),
    .I0(__936__),
    .O(__2820__)
  );
  LUT5 #(
    .INIT(32'hff44f0f0)
  ) __6201__ (
    .I4(g35),
    .I3(__2797__),
    .I2(__173__),
    .I1(__549__),
    .I0(__2254__),
    .O(__2821__)
  );
  LUT5 #(
    .INIT(32'hfff8ffff)
  ) __6202__ (
    .I4(g35),
    .I3(__84__),
    .I2(__1512__),
    .I1(__913__),
    .I0(__486__),
    .O(__2822__)
  );
  LUT4 #(
    .INIT(16'h7da0)
  ) __6203__ (
    .I3(__1233__),
    .I2(__770__),
    .I1(__385__),
    .I0(g35),
    .O(__2823__)
  );
  LUT6 #(
    .INIT(64'h5adaaa2affff0000)
  ) __6204__ (
    .I5(g35),
    .I4(__1048__),
    .I3(__653__),
    .I2(__1708__),
    .I1(__934__),
    .I0(__894__),
    .O(__2824__)
  );
  LUT5 #(
    .INIT(32'h3caaf0f0)
  ) __6205__ (
    .I4(g35),
    .I3(__2281__),
    .I2(__1234__),
    .I1(__178__),
    .I0(__1265__),
    .O(__2825__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6206__ (
    .I2(__254__),
    .I1(__729__),
    .I0(__1017__),
    .O(__2826__)
  );
  LUT6 #(
    .INIT(64'hebaa00aa00000000)
  ) __6207__ (
    .I5(g35),
    .I4(__2178__),
    .I3(__1630__),
    .I2(__527__),
    .I1(__2826__),
    .I0(__889__),
    .O(__2827__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6208__ (
    .I2(g35),
    .I1(__1153__),
    .I0(__1159__),
    .O(__2828__)
  );
  LUT3 #(
    .INIT(8'he0)
  ) __6209__ (
    .I2(g35),
    .I1(__1171__),
    .I0(__455__),
    .O(__2829__)
  );
  LUT3 #(
    .INIT(8'he0)
  ) __6210__ (
    .I2(g35),
    .I1(__201__),
    .I0(__292__),
    .O(__2830__)
  );
  LUT3 #(
    .INIT(8'he0)
  ) __6211__ (
    .I2(g35),
    .I1(__846__),
    .I0(__1133__),
    .O(__2831__)
  );
  LUT5 #(
    .INIT(32'hfffefee0)
  ) __6212__ (
    .I4(__2831__),
    .I3(__2830__),
    .I2(__2829__),
    .I1(__368__),
    .I0(__1155__),
    .O(__2832__)
  );
  LUT3 #(
    .INIT(8'he0)
  ) __6213__ (
    .I2(g35),
    .I1(__571__),
    .I0(__424__),
    .O(__2833__)
  );
  LUT5 #(
    .INIT(32'h01010157)
  ) __6214__ (
    .I4(__971__),
    .I3(__567__),
    .I2(__1076__),
    .I1(__167__),
    .I0(__2833__),
    .O(__2834__)
  );
  LUT6 #(
    .INIT(64'h000000000000001f)
  ) __6215__ (
    .I5(__2831__),
    .I4(__2830__),
    .I3(__2829__),
    .I2(g35),
    .I1(__368__),
    .I0(__1155__),
    .O(__2835__)
  );
  LUT3 #(
    .INIT(8'he0)
  ) __6216__ (
    .I2(g35),
    .I1(__903__),
    .I0(__512__),
    .O(__2836__)
  );
  LUT6 #(
    .INIT(64'h000000000001ffff)
  ) __6217__ (
    .I5(__2833__),
    .I4(g35),
    .I3(__971__),
    .I2(__1076__),
    .I1(__567__),
    .I0(__167__),
    .O(__2837__)
  );
  LUT5 #(
    .INIT(32'hc05500c0)
  ) __6218__ (
    .I4(__2837__),
    .I3(__2836__),
    .I2(__2835__),
    .I1(__2834__),
    .I0(__2832__),
    .O(__2838__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __6219__ (
    .I1(__900__),
    .I0(__817__),
    .O(__2839__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6220__ (
    .I5(g35),
    .I4(__2839__),
    .I3(__1417__),
    .I2(__1096__),
    .I1(__1239__),
    .I0(__1391__),
    .O(__2840__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6221__ (
    .I1(__555__),
    .I0(__713__),
    .O(__2841__)
  );
  LUT6 #(
    .INIT(64'hf0ff00ffffff7777)
  ) __6222__ (
    .I5(__437__),
    .I4(__1398__),
    .I3(__2346__),
    .I2(__1029__),
    .I1(__289__),
    .I0(__2841__),
    .O(__2842__)
  );
  LUT6 #(
    .INIT(64'hf57f554400000000)
  ) __6223__ (
    .I5(g35),
    .I4(__35__),
    .I3(__631__),
    .I2(__299__),
    .I1(__736__),
    .I0(__2842__),
    .O(__2843__)
  );
  LUT6 #(
    .INIT(64'hff00df10ffff0000)
  ) __6224__ (
    .I5(g35),
    .I4(__817__),
    .I3(__1239__),
    .I2(__1852__),
    .I1(__900__),
    .I0(__1391__),
    .O(__2844__)
  );
  LUT5 #(
    .INIT(32'h0af0cccc)
  ) __6225__ (
    .I4(g35),
    .I3(__575__),
    .I2(__2373__),
    .I1(__277__),
    .I0(__2372__),
    .O(__2845__)
  );
  LUT4 #(
    .INIT(16'h3caa)
  ) __6226__ (
    .I3(g35),
    .I2(__897__),
    .I1(__2040__),
    .I0(__346__),
    .O(__2846__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6227__ (
    .I5(g35),
    .I4(__2806__),
    .I3(__2304__),
    .I2(__545__),
    .I1(__311__),
    .I0(__1391__),
    .O(__2847__)
  );
  LUT4 #(
    .INIT(16'h070c)
  ) __6228__ (
    .I3(__282__),
    .I2(__452__),
    .I1(__132__),
    .I0(__356__),
    .O(__2848__)
  );
  LUT6 #(
    .INIT(64'h00ff33330f0f5555)
  ) __6229__ (
    .I5(__282__),
    .I4(__132__),
    .I3(__1039__),
    .I2(__1071__),
    .I1(__508__),
    .I0(__161__),
    .O(__2849__)
  );
  LUT6 #(
    .INIT(64'hcccccffc00ff5555)
  ) __6230__ (
    .I5(__347__),
    .I4(__32__),
    .I3(__1292__),
    .I2(__2849__),
    .I1(__452__),
    .I0(__2848__),
    .O(__2850__)
  );
  LUT3 #(
    .INIT(8'h01)
  ) __6231__ (
    .I2(__52__),
    .I1(__124__),
    .I0(__21__),
    .O(__2851__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __6232__ (
    .I1(__124__),
    .I0(__1083__),
    .O(__2852__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6233__ (
    .I1(__21__),
    .I0(__809__),
    .O(__2853__)
  );
  LUT6 #(
    .INIT(64'h0000000000005f13)
  ) __6234__ (
    .I5(__2853__),
    .I4(__2852__),
    .I3(__549__),
    .I2(__52__),
    .I1(__706__),
    .I0(__247__),
    .O(__2854__)
  );
  LUT5 #(
    .INIT(32'h10ff0000)
  ) __6235__ (
    .I4(g35),
    .I3(__2854__),
    .I2(__2851__),
    .I1(__706__),
    .I0(__2850__),
    .O(__2855__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6236__ (
    .I1(__91__),
    .I0(__358__),
    .O(__2856__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __6237__ (
    .I1(__402__),
    .I0(__91__),
    .O(__2857__)
  );
  LUT6 #(
    .INIT(64'hffccff00f0f0fafa)
  ) __6238__ (
    .I5(__711__),
    .I4(__13__),
    .I3(__2857__),
    .I2(__2856__),
    .I1(__668__),
    .I0(__669__),
    .O(__2858__)
  );
  LUT5 #(
    .INIT(32'h0f05030f)
  ) __6239__ (
    .I4(__13__),
    .I3(__91__),
    .I2(__2858__),
    .I1(__1241__),
    .I0(__988__),
    .O(__2859__)
  );
  LUT5 #(
    .INIT(32'h33aaf0f0)
  ) __6240__ (
    .I4(g35),
    .I3(__1718__),
    .I2(__13__),
    .I1(__2859__),
    .I0(__974__),
    .O(__2860__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __6241__ (
    .I1(__482__),
    .I0(__794__),
    .O(__2861__)
  );
  LUT6 #(
    .INIT(64'h000078f0aaaaaaaa)
  ) __6242__ (
    .I5(g35),
    .I4(__1776__),
    .I3(__1268__),
    .I2(__1052__),
    .I1(__2861__),
    .I0(__702__),
    .O(__2862__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __6243__ (
    .I1(__1217__),
    .I0(__1038__),
    .O(__2863__)
  );
  LUT6 #(
    .INIT(64'h0a03000000000000)
  ) __6244__ (
    .I5(g35),
    .I4(__2863__),
    .I3(__302__),
    .I2(__1162__),
    .I1(__935__),
    .I0(__451__),
    .O(__2864__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6245__ (
    .I5(g35),
    .I4(__2543__),
    .I3(__1704__),
    .I2(__1056__),
    .I1(__1120__),
    .I0(__1391__),
    .O(__2865__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __6246__ (
    .I1(__1681__),
    .I0(__1680__),
    .O(__2866__)
  );
  LUT6 #(
    .INIT(64'h0000000000000004)
  ) __6247__ (
    .I5(__143__),
    .I4(__1205__),
    .I3(__838__),
    .I2(__1070__),
    .I1(__492__),
    .I0(__392__),
    .O(__2867__)
  );
  LUT6 #(
    .INIT(64'h8000000000000000)
  ) __6248__ (
    .I5(__959__),
    .I4(__143__),
    .I3(__1205__),
    .I2(__838__),
    .I1(__1070__),
    .I0(__392__),
    .O(__2868__)
  );
  LUT6 #(
    .INIT(64'h000afff0cccccccc)
  ) __6249__ (
    .I5(g35),
    .I4(__1193__),
    .I3(__2868__),
    .I2(__2867__),
    .I1(__143__),
    .I0(__2866__),
    .O(__2869__)
  );
  LUT6 #(
    .INIT(64'h7fd55555aa000000)
  ) __6250__ (
    .I5(__400__),
    .I4(__875__),
    .I3(__177__),
    .I2(__1451__),
    .I1(__671__),
    .I0(g35),
    .O(__2870__)
  );
  LUT6 #(
    .INIT(64'h22882c8cff00ff00)
  ) __6251__ (
    .I5(g35),
    .I4(__631__),
    .I3(__555__),
    .I2(__736__),
    .I1(__413__),
    .I0(__1832__),
    .O(__2871__)
  );
  LUT5 #(
    .INIT(32'h575d0a00)
  ) __6252__ (
    .I4(__900__),
    .I3(__817__),
    .I2(__2182__),
    .I1(__412__),
    .I0(g35),
    .O(__2872__)
  );
  LUT5 #(
    .INIT(32'habff5400)
  ) __6253__ (
    .I4(__710__),
    .I3(__1115__),
    .I2(__35__),
    .I1(__437__),
    .I0(__667__),
    .O(__2873__)
  );
  LUT6 #(
    .INIT(64'hfa00f0f0cccccccc)
  ) __6254__ (
    .I5(g35),
    .I4(__2260__),
    .I3(__2873__),
    .I2(__1160__),
    .I1(__500__),
    .I0(__1497__),
    .O(__2874__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6255__ (
    .I5(g35),
    .I4(__1620__),
    .I3(__2363__),
    .I2(__272__),
    .I1(__317__),
    .I0(__1391__),
    .O(__2875__)
  );
  LUT5 #(
    .INIT(32'h33aaf0f0)
  ) __6256__ (
    .I4(g35),
    .I3(__1958__),
    .I2(__829__),
    .I1(__1827__),
    .I0(__1051__),
    .O(__2876__)
  );
  LUT6 #(
    .INIT(64'h0000000000000080)
  ) __6257__ (
    .I5(g113),
    .I4(__1283__),
    .I3(__757__),
    .I2(__1385__),
    .I1(__236__),
    .I0(__810__),
    .O(__2877__)
  );
  LUT5 #(
    .INIT(32'h575d0a00)
  ) __6258__ (
    .I4(__689__),
    .I3(__253__),
    .I2(__2877__),
    .I1(__623__),
    .I0(g35),
    .O(__2878__)
  );
  LUT5 #(
    .INIT(32'hff44f0f0)
  ) __6259__ (
    .I4(g35),
    .I3(__2537__),
    .I2(__1278__),
    .I1(__1083__),
    .I0(__2301__),
    .O(__2879__)
  );
  LUT5 #(
    .INIT(32'haaf030f0)
  ) __6260__ (
    .I4(__1600__),
    .I3(g35),
    .I2(__1027__),
    .I1(__2489__),
    .I0(__944__),
    .O(__2880__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __6261__ (
    .I2(g35),
    .I1(__940__),
    .I0(__1245__),
    .O(__2881__)
  );
  LUT6 #(
    .INIT(64'h337fb3b300cc0000)
  ) __6262__ (
    .I5(__1113__),
    .I4(__854__),
    .I3(__1788__),
    .I2(__207__),
    .I1(g35),
    .I0(__2270__),
    .O(__2882__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6263__ (
    .I1(g35),
    .I0(__961__),
    .O(__2883__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6264__ (
    .I2(__726__),
    .I1(__1066__),
    .I0(__12__),
    .O(__2884__)
  );
  LUT6 #(
    .INIT(64'hebaa00aa00000000)
  ) __6265__ (
    .I5(g35),
    .I4(__2695__),
    .I3(__2254__),
    .I2(__830__),
    .I1(__2884__),
    .I0(__679__),
    .O(__2885__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6266__ (
    .I5(g35),
    .I4(__2543__),
    .I3(__2263__),
    .I2(__165__),
    .I1(__172__),
    .I0(__1391__),
    .O(__2886__)
  );
  LUT6 #(
    .INIT(64'h337fb3b300cc0000)
  ) __6267__ (
    .I5(__226__),
    .I4(__799__),
    .I3(__1788__),
    .I2(__716__),
    .I1(g35),
    .I0(__2441__),
    .O(__2887__)
  );
  LUT5 #(
    .INIT(32'hc3aaf0f0)
  ) __6268__ (
    .I4(g35),
    .I3(__2057__),
    .I2(__676__),
    .I1(__915__),
    .I0(__567__),
    .O(__2888__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __6269__ (
    .I1(__343__),
    .I0(__92__),
    .O(__2889__)
  );
  LUT6 #(
    .INIT(64'h0000000000004000)
  ) __6270__ (
    .I5(__871__),
    .I4(__114__),
    .I3(__702__),
    .I2(__2308__),
    .I1(__2889__),
    .I0(__301__),
    .O(__2890__)
  );
  LUT3 #(
    .INIT(8'h01)
  ) __6271__ (
    .I2(__1240__),
    .I1(__738__),
    .I0(__976__),
    .O(__2891__)
  );
  LUT6 #(
    .INIT(64'h80008000ffff0000)
  ) __6272__ (
    .I5(g35),
    .I4(__1236__),
    .I3(__2861__),
    .I2(__2891__),
    .I1(__582__),
    .I0(__2890__),
    .O(__2892__)
  );
  LUT6 #(
    .INIT(64'heaaa2aaaffff0000)
  ) __6273__ (
    .I5(g35),
    .I4(__154__),
    .I3(__412__),
    .I2(__900__),
    .I1(__817__),
    .I0(__178__),
    .O(__2893__)
  );
  LUT6 #(
    .INIT(64'h6c206c6cf0f0f0f0)
  ) __6274__ (
    .I5(g35),
    .I4(__751__),
    .I3(__869__),
    .I2(__981__),
    .I1(__33__),
    .I0(__1455__),
    .O(__2894__)
  );
  LUT5 #(
    .INIT(32'h5df080f0)
  ) __6275__ (
    .I4(__1029__),
    .I3(g35),
    .I2(__319__),
    .I1(__437__),
    .I0(__2029__),
    .O(__2895__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6276__ (
    .I5(g35),
    .I4(__1866__),
    .I3(__2450__),
    .I2(__370__),
    .I1(__677__),
    .I0(__1391__),
    .O(__2896__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6277__ (
    .I2(__2582__),
    .I1(__77__),
    .I0(__584__),
    .O(__2897__)
  );
  LUT4 #(
    .INIT(16'h77f0)
  ) __6278__ (
    .I3(g35),
    .I2(__551__),
    .I1(__718__),
    .I0(__650__),
    .O(__2898__)
  );
  LUT5 #(
    .INIT(32'h7df05500)
  ) __6279__ (
    .I4(__1549__),
    .I3(__403__),
    .I2(__414__),
    .I1(__2729__),
    .I0(g35),
    .O(__2899__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6280__ (
    .I1(g35),
    .I0(__817__),
    .O(__2900__)
  );
  LUT6 #(
    .INIT(64'h3fffc000aaaaaaaa)
  ) __6281__ (
    .I5(g35),
    .I4(__1119__),
    .I3(__653__),
    .I2(__1237__),
    .I1(__1708__),
    .I0(__947__),
    .O(__2901__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6282__ (
    .I5(g35),
    .I4(__1964__),
    .I3(__2548__),
    .I2(__986__),
    .I1(__47__),
    .I0(__1391__),
    .O(__2902__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6283__ (
    .I2(g35),
    .I1(__840__),
    .I0(__730__),
    .O(__2903__)
  );
  LUT6 #(
    .INIT(64'hf0f04444ff00ff00)
  ) __6284__ (
    .I5(g35),
    .I4(__1638__),
    .I3(__651__),
    .I2(__617__),
    .I1(__1269__),
    .I0(__2461__),
    .O(__2904__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6285__ (
    .I5(g35),
    .I4(__950__),
    .I3(__1474__),
    .I2(__1059__),
    .I1(__834__),
    .I0(__1470__),
    .O(__2905__)
  );
  LUT5 #(
    .INIT(32'hfffe0000)
  ) __6286__ (
    .I4(g35),
    .I3(__322__),
    .I2(__470__),
    .I1(__260__),
    .I0(__16__),
    .O(__2906__)
  );
  LUT6 #(
    .INIT(64'h000000000001ffff)
  ) __6287__ (
    .I5(__2906__),
    .I4(g35),
    .I3(__844__),
    .I2(__947__),
    .I1(__1094__),
    .I0(__745__),
    .O(__2907__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __6288__ (
    .I1(__1722__),
    .I0(__1724__),
    .O(__2908__)
  );
  LUT5 #(
    .INIT(32'h0040c0c0)
  ) __6289__ (
    .I4(g35),
    .I3(__903__),
    .I2(__2837__),
    .I1(__2835__),
    .I0(__512__),
    .O(__2909__)
  );
  LUT6 #(
    .INIT(64'h0000000000008000)
  ) __6290__ (
    .I5(__264__),
    .I4(__249__),
    .I3(__2909__),
    .I2(__2908__),
    .I1(__2614__),
    .I0(__2907__),
    .O(__2910__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __6291__ (
    .I2(g35),
    .I1(__2910__),
    .I0(__44__),
    .O(__2911__)
  );
  LUT5 #(
    .INIT(32'h0af0cccc)
  ) __6292__ (
    .I4(g35),
    .I3(__210__),
    .I2(__1539__),
    .I1(__129__),
    .I0(__1541__),
    .O(__2912__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6293__ (
    .I5(g35),
    .I4(__2304__),
    .I3(__2450__),
    .I2(__522__),
    .I1(__545__),
    .I0(__1391__),
    .O(__2913__)
  );
  LUT6 #(
    .INIT(64'hfffcffffaaaaaaaa)
  ) __6294__ (
    .I5(g35),
    .I4(__1249__),
    .I3(__304__),
    .I2(__529__),
    .I1(__40__),
    .I0(__1260__),
    .O(__2914__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6295__ (
    .I5(g35),
    .I4(__2026__),
    .I3(__2546__),
    .I2(__1129__),
    .I1(__408__),
    .I0(__1391__),
    .O(__2915__)
  );
  LUT4 #(
    .INIT(16'h1caa)
  ) __6296__ (
    .I3(g35),
    .I2(__1757__),
    .I1(__659__),
    .I0(__1144__),
    .O(__2916__)
  );
  LUT5 #(
    .INIT(32'h575d0a00)
  ) __6297__ (
    .I4(__509__),
    .I3(__705__),
    .I2(__2477__),
    .I1(__306__),
    .I0(g35),
    .O(__2917__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __6298__ (
    .I2(g35),
    .I1(__1680__),
    .I0(__11__),
    .O(__2918__)
  );
  LUT5 #(
    .INIT(32'hff44f0f0)
  ) __6299__ (
    .I4(g35),
    .I3(__1331__),
    .I2(__831__),
    .I1(__663__),
    .I0(__1311__),
    .O(__2919__)
  );
  LUT6 #(
    .INIT(64'h0fff7f0070ff0000)
  ) __6300__ (
    .I5(__820__),
    .I4(__511__),
    .I3(g35),
    .I2(__1673__),
    .I1(__1338__),
    .I0(__2758__),
    .O(__2920__)
  );
  LUT6 #(
    .INIT(64'h00dfdf00ffff0000)
  ) __6301__ (
    .I5(g35),
    .I4(__989__),
    .I3(__313__),
    .I2(__1303__),
    .I1(__810__),
    .I0(__1670__),
    .O(__2921__)
  );
  LUT6 #(
    .INIT(64'h0000000000000008)
  ) __6302__ (
    .I5(__917__),
    .I4(__972__),
    .I3(g113),
    .I2(__1283__),
    .I1(__1286__),
    .I0(__1282__),
    .O(__2922__)
  );
  LUT6 #(
    .INIT(64'hf30caaaaf0f0f0f0)
  ) __6303__ (
    .I5(g35),
    .I4(__2922__),
    .I3(__749__),
    .I2(__819__),
    .I1(__982__),
    .I0(__543__),
    .O(__2923__)
  );
  LUT6 #(
    .INIT(64'hefffefffffff0000)
  ) __6304__ (
    .I5(g35),
    .I4(__264__),
    .I3(g91),
    .I2(__1841__),
    .I1(__694__),
    .I0(__1843__),
    .O(__2924__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6305__ (
    .I5(g35),
    .I4(__457__),
    .I3(__2264__),
    .I2(__164__),
    .I1(__268__),
    .I0(__1391__),
    .O(__2925__)
  );
  LUT5 #(
    .INIT(32'hccaaf0f0)
  ) __6306__ (
    .I4(g35),
    .I3(__1451__),
    .I2(__159__),
    .I1(__34__),
    .I0(__97__),
    .O(__2926__)
  );
  LUT4 #(
    .INIT(16'heef0)
  ) __6307__ (
    .I3(g35),
    .I2(__221__),
    .I1(__280__),
    .I0(__113__),
    .O(__2927__)
  );
  LUT6 #(
    .INIT(64'h0077ff00f0f0f0f0)
  ) __6308__ (
    .I5(g35),
    .I4(__2254__),
    .I3(__726__),
    .I2(__1066__),
    .I1(__1338__),
    .I0(__2697__),
    .O(__2928__)
  );
  LUT6 #(
    .INIT(64'h06666666aaaaaaaa)
  ) __6309__ (
    .I5(g35),
    .I4(__1303__),
    .I3(__810__),
    .I2(__1670__),
    .I1(__689__),
    .I0(__623__),
    .O(__2929__)
  );
  LUT6 #(
    .INIT(64'hdfffffffcfffffff)
  ) __6310__ (
    .I5(__1370__),
    .I4(__2150__),
    .I3(__2149__),
    .I2(__680__),
    .I1(__2146__),
    .I0(__2142__),
    .O(__2930__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6311__ (
    .I2(g35),
    .I1(g6750),
    .I0(__389__),
    .O(__2931__)
  );
  LUT5 #(
    .INIT(32'hc3aaf0f0)
  ) __6312__ (
    .I4(g35),
    .I3(__1556__),
    .I2(__82__),
    .I1(__1230__),
    .I0(__965__),
    .O(__2932__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6313__ (
    .I5(g35),
    .I4(__1708__),
    .I3(__2499__),
    .I2(__732__),
    .I1(__675__),
    .I0(__1640__),
    .O(__2933__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6314__ (
    .I2(g35),
    .I1(__214__),
    .I0(__739__),
    .O(__2934__)
  );
  LUT3 #(
    .INIT(8'h01)
  ) __6315__ (
    .I2(__860__),
    .I1(__1111__),
    .I0(__1782__),
    .O(__2935__)
  );
  LUT5 #(
    .INIT(32'hc3aaf0f0)
  ) __6316__ (
    .I4(g35),
    .I3(__2935__),
    .I2(__562__),
    .I1(__743__),
    .I0(__861__),
    .O(__2936__)
  );
  LUT6 #(
    .INIT(64'hc3aaaaaaf0f0f0f0)
  ) __6317__ (
    .I5(g35),
    .I4(__2255__),
    .I3(__2254__),
    .I2(__61__),
    .I1(__434__),
    .I0(__424__),
    .O(__2937__)
  );
  LUT6 #(
    .INIT(64'h3f3f002affff00aa)
  ) __6318__ (
    .I5(__972__),
    .I4(__1164__),
    .I3(__964__),
    .I2(__1444__),
    .I1(__1465__),
    .I0(__1114__),
    .O(__2938__)
  );
  LUT5 #(
    .INIT(32'h33aaf0f0)
  ) __6319__ (
    .I4(g35),
    .I3(__1383__),
    .I2(__581__),
    .I1(__2938__),
    .I0(__964__),
    .O(__2939__)
  );
  LUT6 #(
    .INIT(64'h0000000000000008)
  ) __6320__ (
    .I5(g113),
    .I4(__1283__),
    .I3(__757__),
    .I2(__810__),
    .I1(__236__),
    .I0(__2054__),
    .O(__2940__)
  );
  LUT5 #(
    .INIT(32'h10ff0000)
  ) __6321__ (
    .I4(__386__),
    .I3(g35),
    .I2(__798__),
    .I1(__1145__),
    .I0(__2940__),
    .O(__2941__)
  );
  LUT4 #(
    .INIT(16'hbf00)
  ) __6322__ (
    .I3(g35),
    .I2(__84__),
    .I1(__486__),
    .I0(__1512__),
    .O(__2942__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6323__ (
    .I5(g35),
    .I4(__2548__),
    .I3(__1793__),
    .I2(__1090__),
    .I1(__807__),
    .I0(__1391__),
    .O(__2943__)
  );
  LUT3 #(
    .INIT(8'h78)
  ) __6324__ (
    .I2(__476__),
    .I1(g35),
    .I0(__1138__),
    .O(__2944__)
  );
  LUT4 #(
    .INIT(16'h8000)
  ) __6325__ (
    .I3(__972__),
    .I2(__1383__),
    .I1(__1503__),
    .I0(__1465__),
    .O(__2945__)
  );
  LUT6 #(
    .INIT(64'hf30caaaaf0f0f0f0)
  ) __6326__ (
    .I5(g35),
    .I4(__2945__),
    .I3(__749__),
    .I2(__1114__),
    .I1(__1164__),
    .I0(__984__),
    .O(__2946__)
  );
  LUT3 #(
    .INIT(8'hf4)
  ) __6327__ (
    .I2(__2416__),
    .I1(__9__),
    .I0(g35),
    .O(__2947__)
  );
  LUT6 #(
    .INIT(64'hbfffffff00000000)
  ) __6328__ (
    .I5(__21__),
    .I4(g35),
    .I3(__1503__),
    .I2(__1567__),
    .I1(__15__),
    .I0(__1240__),
    .O(__2948__)
  );
  LUT5 #(
    .INIT(32'hccaaf0f0)
  ) __6329__ (
    .I4(g35),
    .I3(__1864__),
    .I2(__501__),
    .I1(__371__),
    .I0(__410__),
    .O(__2949__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6330__ (
    .I5(g35),
    .I4(__2027__),
    .I3(__1790__),
    .I2(__905__),
    .I1(__735__),
    .I0(__1391__),
    .O(__2950__)
  );
  LUT6 #(
    .INIT(64'heeeef0f0ff00ff00)
  ) __6331__ (
    .I5(g35),
    .I4(__1299__),
    .I3(__925__),
    .I2(__541__),
    .I1(__760__),
    .I0(__1710__),
    .O(__2951__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __6332__ (
    .I1(__357__),
    .I0(__613__),
    .O(__2952__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6333__ (
    .I5(g35),
    .I4(__2952__),
    .I3(__1611__),
    .I2(__430__),
    .I1(__761__),
    .I0(__1391__),
    .O(__2953__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __6334__ (
    .I2(__530__),
    .I1(__882__),
    .I0(__389__),
    .O(__2954__)
  );
  LUT5 #(
    .INIT(32'hfefeff00)
  ) __6335__ (
    .I4(__341__),
    .I3(__1213__),
    .I2(g72),
    .I1(g73),
    .I0(__824__),
    .O(__2955__)
  );
  LUT6 #(
    .INIT(64'heeaaff00f0f0ff00)
  ) __6336__ (
    .I5(__1689__),
    .I4(g35),
    .I3(__378__),
    .I2(__2955__),
    .I1(__2954__),
    .I0(__796__),
    .O(__2956__)
  );
  LUT6 #(
    .INIT(64'hc0c0c0cd00000000)
  ) __6337__ (
    .I5(g35),
    .I4(__944__),
    .I3(__2489__),
    .I2(__1600__),
    .I1(__296__),
    .I0(__1027__),
    .O(__2957__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __6338__ (
    .I2(g35),
    .I1(__912__),
    .I0(__36__),
    .O(__2958__)
  );
  LUT5 #(
    .INIT(32'h575d0a00)
  ) __6339__ (
    .I4(__788__),
    .I3(__1077__),
    .I2(__1441__),
    .I1(__1857__),
    .I0(g35),
    .O(__2959__)
  );
  LUT4 #(
    .INIT(16'heef0)
  ) __6340__ (
    .I3(g35),
    .I2(__428__),
    .I1(__432__),
    .I0(__616__),
    .O(__2960__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6341__ (
    .I5(g35),
    .I4(__2046__),
    .I3(__2548__),
    .I2(__565__),
    .I1(__1064__),
    .I0(__1391__),
    .O(__2961__)
  );
  LUT6 #(
    .INIT(64'h00dfdf00ffff0000)
  ) __6342__ (
    .I5(g35),
    .I4(__157__),
    .I3(__863__),
    .I2(__1773__),
    .I1(__810__),
    .I0(__1303__),
    .O(__2962__)
  );
  LUT5 #(
    .INIT(32'h3caaf0f0)
  ) __6343__ (
    .I4(g35),
    .I3(__1897__),
    .I2(__1210__),
    .I1(__449__),
    .I0(__1008__),
    .O(__2963__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6344__ (
    .I1(g35),
    .I0(__895__),
    .O(__2964__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __6345__ (
    .I1(__540__),
    .I0(__1521__),
    .O(__2965__)
  );
  LUT6 #(
    .INIT(64'hf055f0f0cccccccc)
  ) __6346__ (
    .I5(g35),
    .I4(__2965__),
    .I3(__595__),
    .I2(__1277__),
    .I1(__837__),
    .I0(__1827__),
    .O(__2966__)
  );
  LUT5 #(
    .INIT(32'h00000080)
  ) __6347__ (
    .I4(__1077__),
    .I3(__721__),
    .I2(__69__),
    .I1(__288__),
    .I0(__788__),
    .O(__2967__)
  );
  LUT6 #(
    .INIT(64'hccccf0aaf0f0f0f0)
  ) __6348__ (
    .I5(g35),
    .I4(__2179__),
    .I3(__2967__),
    .I2(__572__),
    .I1(__1279__),
    .I0(__780__),
    .O(__2968__)
  );
  LUT6 #(
    .INIT(64'h3fffc000aaaaaaaa)
  ) __6349__ (
    .I5(g35),
    .I4(__1253__),
    .I3(__1299__),
    .I2(__541__),
    .I1(__1197__),
    .I0(__260__),
    .O(__2969__)
  );
  LUT4 #(
    .INIT(16'h11f0)
  ) __6350__ (
    .I3(g35),
    .I2(__84__),
    .I1(__913__),
    .I0(__486__),
    .O(__2970__)
  );
  LUT4 #(
    .INIT(16'h3caa)
  ) __6351__ (
    .I3(g35),
    .I2(__62__),
    .I1(__1306__),
    .I0(__536__),
    .O(__2971__)
  );
  LUT6 #(
    .INIT(64'hccccf0aaf0f0f0f0)
  ) __6352__ (
    .I5(g35),
    .I4(__2179__),
    .I3(__2318__),
    .I2(__229__),
    .I1(__1279__),
    .I0(__727__),
    .O(__2972__)
  );
  LUT6 #(
    .INIT(64'hf055f0f0cccccccc)
  ) __6353__ (
    .I5(g35),
    .I4(__2643__),
    .I3(__908__),
    .I2(__111__),
    .I1(__1122__),
    .I0(__2034__),
    .O(__2973__)
  );
  LUT5 #(
    .INIT(32'h00cef0f0)
  ) __6354__ (
    .I4(g35),
    .I3(__189__),
    .I2(__857__),
    .I1(__619__),
    .I0(__1184__),
    .O(__2974__)
  );
  LUT6 #(
    .INIT(64'h3fffc000aaaaaaaa)
  ) __6355__ (
    .I5(g35),
    .I4(__1206__),
    .I3(__412__),
    .I2(__900__),
    .I1(__817__),
    .I0(__1265__),
    .O(__2975__)
  );
  LUT6 #(
    .INIT(64'h3fffc000aaaaaaaa)
  ) __6356__ (
    .I5(g35),
    .I4(__872__),
    .I3(__457__),
    .I2(__874__),
    .I1(__1264__),
    .I0(__750__),
    .O(__2976__)
  );
  LUT6 #(
    .INIT(64'heeeef0f0ff00ff00)
  ) __6357__ (
    .I5(g35),
    .I4(__1286__),
    .I3(__543__),
    .I2(__982__),
    .I1(__819__),
    .I0(__1284__),
    .O(__2977__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6358__ (
    .I2(g35),
    .I1(__1260__),
    .I0(__291__),
    .O(__2978__)
  );
  LUT5 #(
    .INIT(32'hccaaf0f0)
  ) __6359__ (
    .I4(g35),
    .I3(__1864__),
    .I2(__538__),
    .I1(__419__),
    .I0(__149__),
    .O(__2979__)
  );
  LUT6 #(
    .INIT(64'heaaa2aaaffff0000)
  ) __6360__ (
    .I5(g35),
    .I4(__850__),
    .I3(__1299__),
    .I2(__541__),
    .I1(__1197__),
    .I0(__893__),
    .O(__2980__)
  );
  LUT5 #(
    .INIT(32'h7d55a000)
  ) __6361__ (
    .I4(__955__),
    .I3(__2372__),
    .I2(__1203__),
    .I1(__2371__),
    .I0(g35),
    .O(__2981__)
  );
  LUT6 #(
    .INIT(64'h0f0f4f4fff00ff00)
  ) __6362__ (
    .I5(g35),
    .I4(__706__),
    .I3(__1280__),
    .I2(__2854__),
    .I1(__2851__),
    .I0(__2850__),
    .O(__2982__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __6363__ (
    .I1(__793__),
    .I0(__1555__),
    .O(__2983__)
  );
  LUT6 #(
    .INIT(64'hf055f0f0cccccccc)
  ) __6364__ (
    .I5(g35),
    .I4(__2983__),
    .I3(__352__),
    .I2(__358__),
    .I1(__668__),
    .I0(__1552__),
    .O(__2984__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6365__ (
    .I2(g35),
    .I1(__897__),
    .I0(__158__),
    .O(__2985__)
  );
  LUT5 #(
    .INIT(32'hccaaf0f0)
  ) __6366__ (
    .I4(g35),
    .I3(__170__),
    .I2(__99__),
    .I1(__204__),
    .I0(__717__),
    .O(__2986__)
  );
  LUT6 #(
    .INIT(64'h000014f0cccccccc)
  ) __6367__ (
    .I5(g35),
    .I4(__1776__),
    .I3(__1871__),
    .I2(__114__),
    .I1(__343__),
    .I0(__301__),
    .O(__2987__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6368__ (
    .I5(g35),
    .I4(__2361__),
    .I3(__2516__),
    .I2(__51__),
    .I1(__202__),
    .I0(__1391__),
    .O(__2988__)
  );
  LUT4 #(
    .INIT(16'h3caa)
  ) __6369__ (
    .I3(g35),
    .I2(__2620__),
    .I1(__1150__),
    .I0(__903__),
    .O(__2989__)
  );
  LUT6 #(
    .INIT(64'haaaaaaaccccccccc)
  ) __6370__ (
    .I5(g35),
    .I4(__860__),
    .I3(__1111__),
    .I2(__1782__),
    .I1(__621__),
    .I0(__273__),
    .O(__2990__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6371__ (
    .I5(g35),
    .I4(__1269__),
    .I3(__2773__),
    .I2(__742__),
    .I1(__145__),
    .I0(__1733__),
    .O(__2991__)
  );
  LUT6 #(
    .INIT(64'heaaa2aaaffff0000)
  ) __6372__ (
    .I5(g35),
    .I4(__1062__),
    .I3(__1430__),
    .I2(__142__),
    .I1(__243__),
    .I0(__1231__),
    .O(__2992__)
  );
  LUT4 #(
    .INIT(16'hbbf0)
  ) __6373__ (
    .I3(g35),
    .I2(__1170__),
    .I1(__2907__),
    .I0(__130__),
    .O(__2993__)
  );
  LUT6 #(
    .INIT(64'h7fffffff00000000)
  ) __6374__ (
    .I5(__1017__),
    .I4(g35),
    .I3(__376__),
    .I2(__1123__),
    .I1(__1627__),
    .I0(__1074__),
    .O(__2994__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6375__ (
    .I5(g35),
    .I4(__1946__),
    .I3(__1612__),
    .I2(__477__),
    .I1(__274__),
    .I0(__1391__),
    .O(__2995__)
  );
  LUT6 #(
    .INIT(64'h0f00afaacccccccc)
  ) __6376__ (
    .I5(g35),
    .I4(__659__),
    .I3(__427__),
    .I2(__479__),
    .I1(__320__),
    .I0(__1757__),
    .O(__2996__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6377__ (
    .I2(g35),
    .I1(__1143__),
    .I0(__961__),
    .O(__2997__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6378__ (
    .I5(g35),
    .I4(__2382__),
    .I3(__1964__),
    .I2(__47__),
    .I1(__808__),
    .I0(__1391__),
    .O(__2998__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6379__ (
    .I5(g35),
    .I4(__2263__),
    .I3(__1761__),
    .I2(__488__),
    .I1(__827__),
    .I0(__1391__),
    .O(__2999__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6380__ (
    .I5(g35),
    .I4(__1633__),
    .I3(__2304__),
    .I2(__309__),
    .I1(__522__),
    .I0(__1391__),
    .O(__3000__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6381__ (
    .I2(g35),
    .I1(__316__),
    .I0(__297__),
    .O(__3001__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __6382__ (
    .I2(__226__),
    .I1(__716__),
    .I0(__2441__),
    .O(__3002__)
  );
  LUT6 #(
    .INIT(64'h6c206c6cf0f0f0f0)
  ) __6383__ (
    .I5(g35),
    .I4(__751__),
    .I3(__869__),
    .I2(__799__),
    .I1(__123__),
    .I0(__3002__),
    .O(__3003__)
  );
  LUT6 #(
    .INIT(64'hc3aaaaaaf0f0f0f0)
  ) __6384__ (
    .I5(g35),
    .I4(__2288__),
    .I3(__1678__),
    .I2(__1221__),
    .I1(__1206__),
    .I0(__1171__),
    .O(__3004__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6385__ (
    .I5(g35),
    .I4(__306__),
    .I3(__2000__),
    .I2(__1137__),
    .I1(__475__),
    .I0(__1391__),
    .O(__3005__)
  );
  LUT4 #(
    .INIT(16'heef0)
  ) __6386__ (
    .I3(g35),
    .I2(__778__),
    .I1(__448__),
    .I0(__384__),
    .O(__3006__)
  );
  LUT5 #(
    .INIT(32'h33aaf0f0)
  ) __6387__ (
    .I4(g35),
    .I3(__2484__),
    .I2(__1139__),
    .I1(__1470__),
    .I0(__532__),
    .O(__3007__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6388__ (
    .I5(g35),
    .I4(__2448__),
    .I3(__2546__),
    .I2(__335__),
    .I1(__977__),
    .I0(__1391__),
    .O(__3008__)
  );
  LUT4 #(
    .INIT(16'h1f30)
  ) __6389__ (
    .I3(__840__),
    .I2(g35),
    .I1(__471__),
    .I0(__2012__),
    .O(__3009__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6390__ (
    .I5(g35),
    .I4(__2361__),
    .I3(__623__),
    .I2(__27__),
    .I1(__162__),
    .I0(__1391__),
    .O(__3010__)
  );
  LUT2 #(
    .INIT(4'hb)
  ) __6391__ (
    .I1(__680__),
    .I0(__2082__),
    .O(__3011__)
  );
  LUT5 #(
    .INIT(32'h00cef0f0)
  ) __6392__ (
    .I4(g35),
    .I3(__559__),
    .I2(__93__),
    .I1(__959__),
    .I0(__401__),
    .O(__3012__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __6393__ (
    .I1(__352__),
    .I0(__793__),
    .O(__3013__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __6394__ (
    .I1(__91__),
    .I0(__13__),
    .O(__3014__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6395__ (
    .I5(g35),
    .I4(__1718__),
    .I3(__3014__),
    .I2(__737__),
    .I1(__669__),
    .I0(__3013__),
    .O(__3015__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6396__ (
    .I5(g35),
    .I4(__2363__),
    .I3(__1742__),
    .I2(__670__),
    .I1(__421__),
    .I0(__1391__),
    .O(__3016__)
  );
  LUT3 #(
    .INIT(8'hc5)
  ) __6397__ (
    .I2(__54__),
    .I1(g116),
    .I0(g115),
    .O(__3017__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6398__ (
    .I2(__54__),
    .I1(g116),
    .I0(g114),
    .O(__3018__)
  );
  LUT5 #(
    .INIT(32'h90999990)
  ) __6399__ (
    .I4(g126),
    .I3(g120),
    .I2(__638__),
    .I1(__3018__),
    .I0(__3017__),
    .O(__3019__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __6400__ (
    .I2(g35),
    .I1(__3019__),
    .I0(__975__),
    .O(__3020__)
  );
  LUT3 #(
    .INIT(8'he0)
  ) __6401__ (
    .I2(g35),
    .I1(__304__),
    .I0(__426__),
    .O(__3021__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6402__ (
    .I1(g35),
    .I0(__468__),
    .O(__3022__)
  );
  LUT6 #(
    .INIT(64'h000000ff0000efef)
  ) __6403__ (
    .I5(__2033__),
    .I4(__1782__),
    .I3(__666__),
    .I2(__1248__),
    .I1(__1485__),
    .I0(__1781__),
    .O(__3023__)
  );
  LUT6 #(
    .INIT(64'h6666666affff0000)
  ) __6404__ (
    .I5(g35),
    .I4(__1111__),
    .I3(__860__),
    .I2(__1782__),
    .I1(__621__),
    .I0(__3023__),
    .O(__3024__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6405__ (
    .I1(__1067__),
    .I0(__2191__),
    .O(__3025__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6406__ (
    .I1(__364__),
    .I0(__2189__),
    .O(__3026__)
  );
  LUT6 #(
    .INIT(64'h7777f0f0ff00ff00)
  ) __6407__ (
    .I5(g35),
    .I4(__1041__),
    .I3(__293__),
    .I2(__3026__),
    .I1(__498__),
    .I0(__3025__),
    .O(__3027__)
  );
  LUT4 #(
    .INIT(16'h3acc)
  ) __6408__ (
    .I3(g35),
    .I2(__188__),
    .I1(__315__),
    .I0(__891__),
    .O(__3028__)
  );
  LUT5 #(
    .INIT(32'h5ffffff3)
  ) __6409__ (
    .I4(__1205__),
    .I3(__838__),
    .I2(__1070__),
    .I1(__492__),
    .I0(__959__),
    .O(__3029__)
  );
  LUT6 #(
    .INIT(64'h000a5555cccccccc)
  ) __6410__ (
    .I5(g35),
    .I4(__392__),
    .I3(__1681__),
    .I2(__1680__),
    .I1(__1070__),
    .I0(__3029__),
    .O(__3030__)
  );
  LUT2 #(
    .INIT(4'h2)
  ) __6411__ (
    .I1(__1280__),
    .I0(g73),
    .O(__3031__)
  );
  LUT6 #(
    .INIT(64'h7777f0f0ff00ff00)
  ) __6412__ (
    .I5(g35),
    .I4(__341__),
    .I3(__180__),
    .I2(__655__),
    .I1(g72),
    .I0(__3031__),
    .O(__3032__)
  );
  LUT5 #(
    .INIT(32'hc3aaf0f0)
  ) __6413__ (
    .I4(g35),
    .I3(__2051__),
    .I2(__1256__),
    .I1(__1089__),
    .I0(__1155__),
    .O(__3033__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6414__ (
    .I1(__203__),
    .I0(__706__),
    .O(__3034__)
  );
  LUT6 #(
    .INIT(64'hf8fff00000ff0000)
  ) __6415__ (
    .I5(__2765__),
    .I4(__447__),
    .I3(g35),
    .I2(__153__),
    .I1(__1235__),
    .I0(__3034__),
    .O(__3035__)
  );
  LUT6 #(
    .INIT(64'hff00df10ffff0000)
  ) __6416__ (
    .I5(g35),
    .I4(__874__),
    .I3(__558__),
    .I2(__2184__),
    .I1(__1264__),
    .I0(__1391__),
    .O(__3036__)
  );
  LUT5 #(
    .INIT(32'habff5400)
  ) __6417__ (
    .I4(__334__),
    .I3(__1041__),
    .I2(__1207__),
    .I1(__936__),
    .I0(__983__),
    .O(__3037__)
  );
  LUT6 #(
    .INIT(64'hcd00ccccf0f0f0f0)
  ) __6418__ (
    .I5(g35),
    .I4(__2755__),
    .I3(__3037__),
    .I2(__88__),
    .I1(__767__),
    .I0(__489__),
    .O(__3038__)
  );
  LUT5 #(
    .INIT(32'hcfdfffff)
  ) __6419__ (
    .I4(__680__),
    .I3(__2072__),
    .I2(__2095__),
    .I1(__2090__),
    .I0(__2086__),
    .O(__3039__)
  );
  LUT5 #(
    .INIT(32'hffa0cfc0)
  ) __6420__ (
    .I4(__383__),
    .I3(__440__),
    .I2(g35),
    .I1(__218__),
    .I0(__36__),
    .O(__3040__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6421__ (
    .I1(__1252__),
    .I0(__1114__),
    .O(__3041__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __6422__ (
    .I1(__145__),
    .I0(__1114__),
    .O(__3042__)
  );
  LUT6 #(
    .INIT(64'hffccff00f0f0fafa)
  ) __6423__ (
    .I5(__964__),
    .I4(__1164__),
    .I3(__3042__),
    .I2(__3041__),
    .I1(__649__),
    .I0(__742__),
    .O(__3043__)
  );
  LUT5 #(
    .INIT(32'h0f05030f)
  ) __6424__ (
    .I4(__1164__),
    .I3(__1114__),
    .I2(__3043__),
    .I1(__307__),
    .I0(__839__),
    .O(__3044__)
  );
  LUT5 #(
    .INIT(32'h33aaf0f0)
  ) __6425__ (
    .I4(g35),
    .I3(__1383__),
    .I2(__1164__),
    .I1(__3044__),
    .I0(__1178__),
    .O(__3045__)
  );
  LUT3 #(
    .INIT(8'h78)
  ) __6426__ (
    .I2(__940__),
    .I1(g35),
    .I0(__924__),
    .O(__3046__)
  );
  LUT6 #(
    .INIT(64'hfffc0003aaaaaaaa)
  ) __6427__ (
    .I5(g35),
    .I4(__460__),
    .I3(__746__),
    .I2(__793__),
    .I1(__1555__),
    .I0(__965__),
    .O(__3047__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6428__ (
    .I5(g35),
    .I4(__1743__),
    .I3(__1620__),
    .I2(__517__),
    .I1(__272__),
    .I0(__1391__),
    .O(__3048__)
  );
  LUT6 #(
    .INIT(64'h8000aaaa7fffffff)
  ) __6429__ (
    .I5(__1275__),
    .I4(__1813__),
    .I3(__1105__),
    .I2(__775__),
    .I1(__766__),
    .I0(__2800__),
    .O(__3049__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __6430__ (
    .I2(g35),
    .I1(__3049__),
    .I0(__766__),
    .O(__3050__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6431__ (
    .I5(g35),
    .I4(__1823__),
    .I3(__1660__),
    .I2(__1214__),
    .I1(__238__),
    .I0(__1391__),
    .O(__3051__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __6432__ (
    .I2(g35),
    .I1(__956__),
    .I0(__304__),
    .O(__3052__)
  );
  LUT6 #(
    .INIT(64'h0000000080000000)
  ) __6433__ (
    .I5(__757__),
    .I4(__605__),
    .I3(__445__),
    .I2(__810__),
    .I1(__2419__),
    .I0(__2420__),
    .O(__3053__)
  );
  LUT4 #(
    .INIT(16'h11f0)
  ) __6434__ (
    .I3(g35),
    .I2(__1082__),
    .I1(__752__),
    .I0(__3053__),
    .O(__3054__)
  );
  LUT3 #(
    .INIT(8'h08)
  ) __6435__ (
    .I2(__794__),
    .I1(__482__),
    .I0(__582__),
    .O(__3055__)
  );
  LUT6 #(
    .INIT(64'h7fffffff00000000)
  ) __6436__ (
    .I5(g35),
    .I4(__1052__),
    .I3(__1236__),
    .I2(__702__),
    .I1(__2307__),
    .I0(__3055__),
    .O(__3056__)
  );
  LUT6 #(
    .INIT(64'hf055f0f0cccccccc)
  ) __6437__ (
    .I5(g35),
    .I4(__2474__),
    .I3(__1638__),
    .I2(__145__),
    .I1(__307__),
    .I0(__1733__),
    .O(__3057__)
  );
  LUT6 #(
    .INIT(64'h00dfdf00ffff0000)
  ) __6438__ (
    .I5(g35),
    .I4(__425__),
    .I3(__267__),
    .I2(__1773__),
    .I1(__810__),
    .I0(__1303__),
    .O(__3058__)
  );
  LUT6 #(
    .INIT(64'h3caaaaaaf0f0f0f0)
  ) __6439__ (
    .I5(g35),
    .I4(__2557__),
    .I3(__1438__),
    .I2(__902__),
    .I1(__1020__),
    .I0(__750__),
    .O(__3059__)
  );
  LUT5 #(
    .INIT(32'h3ff38888)
  ) __6440__ (
    .I4(__803__),
    .I3(__436__),
    .I2(__1687__),
    .I1(g35),
    .I0(__2307__),
    .O(__3060__)
  );
  LUT6 #(
    .INIT(64'h0fff7f0070ff0000)
  ) __6441__ (
    .I5(__691__),
    .I4(__1180__),
    .I3(g35),
    .I2(__1438__),
    .I1(__1338__),
    .I0(__1437__),
    .O(__3061__)
  );
  LUT4 #(
    .INIT(16'h3caa)
  ) __6442__ (
    .I3(g35),
    .I2(__2779__),
    .I1(__271__),
    .I0(__424__),
    .O(__3062__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6443__ (
    .I5(g35),
    .I4(__157__),
    .I3(__2448__),
    .I2(__1079__),
    .I1(__335__),
    .I0(__1391__),
    .O(__3063__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6444__ (
    .I1(__507__),
    .I0(__1032__),
    .O(__3064__)
  );
  LUT6 #(
    .INIT(64'haaf0f0f0cccccccc)
  ) __6445__ (
    .I5(g35),
    .I4(__3064__),
    .I3(__364__),
    .I2(__1018__),
    .I1(__1263__),
    .I0(__396__),
    .O(__3065__)
  );
  LUT6 #(
    .INIT(64'h3fffc000aaaaaaaa)
  ) __6446__ (
    .I5(g35),
    .I4(__1175__),
    .I3(__157__),
    .I2(__561__),
    .I1(__863__),
    .I0(__300__),
    .O(__3066__)
  );
  LUT6 #(
    .INIT(64'hc0c0c0cd00000000)
  ) __6447__ (
    .I5(g35),
    .I4(__318__),
    .I3(__2461__),
    .I2(__1638__),
    .I1(__1269__),
    .I0(__617__),
    .O(__3067__)
  );
  LUT3 #(
    .INIT(8'h35)
  ) __6448__ (
    .I2(__1193__),
    .I1(__2868__),
    .I0(__2867__),
    .O(__3068__)
  );
  LUT6 #(
    .INIT(64'h8cffc80050ff0500)
  ) __6449__ (
    .I5(__11__),
    .I4(__246__),
    .I3(g35),
    .I2(__1193__),
    .I1(__2866__),
    .I0(__3068__),
    .O(__3069__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __6450__ (
    .I1(__209__),
    .I0(g35),
    .O(__3070__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6451__ (
    .I5(g35),
    .I4(__623__),
    .I3(__1946__),
    .I2(__202__),
    .I1(__477__),
    .I0(__1391__),
    .O(__3071__)
  );
  LUT2 #(
    .INIT(4'hb)
  ) __6452__ (
    .I1(__680__),
    .I0(__2109__),
    .O(__3072__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6453__ (
    .I5(g35),
    .I4(__1145__),
    .I3(__1394__),
    .I2(__921__),
    .I1(__86__),
    .I0(__1391__),
    .O(__3073__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6454__ (
    .I5(g35),
    .I4(__1969__),
    .I3(__2690__),
    .I2(__89__),
    .I1(__531__),
    .I0(__1391__),
    .O(__3074__)
  );
  LUT6 #(
    .INIT(64'hefffefffffff0000)
  ) __6455__ (
    .I5(g35),
    .I4(__429__),
    .I3(__2837__),
    .I2(__2835__),
    .I1(__2836__),
    .I0(__722__),
    .O(__3075__)
  );
  LUT6 #(
    .INIT(64'h06cc0000aaaaaaaa)
  ) __6456__ (
    .I5(g35),
    .I4(__758__),
    .I3(__1452__),
    .I2(__1450__),
    .I1(__698__),
    .I0(__397__),
    .O(__3076__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6457__ (
    .I1(__653__),
    .I0(__1237__),
    .O(__3077__)
  );
  LUT6 #(
    .INIT(64'hc3aaaaaaf0f0f0f0)
  ) __6458__ (
    .I5(g35),
    .I4(__3077__),
    .I3(__1708__),
    .I2(__877__),
    .I1(__969__),
    .I0(__1045__),
    .O(__3078__)
  );
  LUT5 #(
    .INIT(32'hd2dd0000)
  ) __6459__ (
    .I4(g35),
    .I3(__1248__),
    .I2(__1245__),
    .I1(__2057__),
    .I0(__539__),
    .O(__3079__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __6460__ (
    .I1(__631__),
    .I0(__736__),
    .O(__3080__)
  );
  LUT6 #(
    .INIT(64'hff004c80f0f0f0f0)
  ) __6461__ (
    .I5(g35),
    .I4(__3080__),
    .I3(__289__),
    .I2(__413__),
    .I1(__1832__),
    .I0(__555__),
    .O(__3081__)
  );
  LUT6 #(
    .INIT(64'h0000ff000000efef)
  ) __6462__ (
    .I5(__1596__),
    .I4(__1600__),
    .I3(__666__),
    .I2(__1248__),
    .I1(__1485__),
    .I0(__1599__),
    .O(__3082__)
  );
  LUT6 #(
    .INIT(64'h6666666affff0000)
  ) __6463__ (
    .I5(g35),
    .I4(__944__),
    .I3(__296__),
    .I2(__1600__),
    .I1(__55__),
    .I0(__3082__),
    .O(__3083__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6464__ (
    .I5(g35),
    .I4(__412__),
    .I3(__2839__),
    .I2(__1136__),
    .I1(__283__),
    .I0(__1391__),
    .O(__3084__)
  );
  LUT6 #(
    .INIT(64'hccccccacaaaaaaaa)
  ) __6465__ (
    .I5(g35),
    .I4(__881__),
    .I3(__660__),
    .I2(__580__),
    .I1(__152__),
    .I0(__985__),
    .O(__3085__)
  );
  LUT6 #(
    .INIT(64'h3fffc000aaaaaaaa)
  ) __6466__ (
    .I5(g35),
    .I4(__1232__),
    .I3(__313__),
    .I2(__569__),
    .I1(__989__),
    .I0(__1008__),
    .O(__3086__)
  );
  LUT6 #(
    .INIT(64'h373fbb330c0c0000)
  ) __6467__ (
    .I5(__33__),
    .I4(__744__),
    .I3(__981__),
    .I2(__1788__),
    .I1(g35),
    .I0(__1455__),
    .O(__3087__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6468__ (
    .I5(g35),
    .I4(__1853__),
    .I3(__1417__),
    .I2(__1047__),
    .I1(__1246__),
    .I0(__1391__),
    .O(__3088__)
  );
  LUT4 #(
    .INIT(16'heef0)
  ) __6469__ (
    .I3(g35),
    .I2(__806__),
    .I1(__968__),
    .I0(__904__),
    .O(__3089__)
  );
  LUT6 #(
    .INIT(64'h77ff0800ff00ff00)
  ) __6470__ (
    .I5(g35),
    .I4(__423__),
    .I3(__952__),
    .I2(__992__),
    .I1(__206__),
    .I0(__878__),
    .O(__3090__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __6471__ (
    .I1(__112__),
    .I0(__1521__),
    .O(__3091__)
  );
  LUT6 #(
    .INIT(64'hf055f0f0cccccccc)
  ) __6472__ (
    .I5(g35),
    .I4(__3091__),
    .I3(__540__),
    .I2(__837__),
    .I1(__1051__),
    .I0(__1827__),
    .O(__3092__)
  );
  LUT3 #(
    .INIT(8'he0)
  ) __6473__ (
    .I2(g35),
    .I1(__662__),
    .I0(__610__),
    .O(__3093__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __6474__ (
    .I1(__122__),
    .I0(__155__),
    .O(__3094__)
  );
  LUT6 #(
    .INIT(64'h0a03000000000000)
  ) __6475__ (
    .I5(g35),
    .I4(__3094__),
    .I3(__474__),
    .I2(__759__),
    .I1(__724__),
    .I0(__379__),
    .O(__3095__)
  );
  LUT3 #(
    .INIT(8'h78)
  ) __6476__ (
    .I2(__276__),
    .I1(g35),
    .I0(__328__),
    .O(__3096__)
  );
  LUT6 #(
    .INIT(64'h40004000ffff0000)
  ) __6477__ (
    .I5(g35),
    .I4(__701__),
    .I3(__10__),
    .I2(__2308__),
    .I1(__2891__),
    .I0(__702__),
    .O(__3097__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6478__ (
    .I5(g35),
    .I4(__898__),
    .I3(__2304__),
    .I2(__699__),
    .I1(__1176__),
    .I0(__1391__),
    .O(__3098__)
  );
  LUT2 #(
    .INIT(4'h2)
  ) __6479__ (
    .I1(__617__),
    .I0(__318__),
    .O(__3099__)
  );
  LUT5 #(
    .INIT(32'h00000008)
  ) __6480__ (
    .I4(g113),
    .I3(__1283__),
    .I2(__779__),
    .I1(__1636__),
    .I0(__1409__),
    .O(__3100__)
  );
  LUT6 #(
    .INIT(64'h0ff0aaaacccccccc)
  ) __6481__ (
    .I5(g35),
    .I4(__3100__),
    .I3(__1060__),
    .I2(__3099__),
    .I1(__1269__),
    .I0(__651__),
    .O(__3101__)
  );
  LUT5 #(
    .INIT(32'hff44f0f0)
  ) __6482__ (
    .I4(g35),
    .I3(__1915__),
    .I2(__1226__),
    .I1(__809__),
    .I0(__1896__),
    .O(__3102__)
  );
  LUT5 #(
    .INIT(32'hccaaf0f0)
  ) __6483__ (
    .I4(g35),
    .I3(__54__),
    .I2(__610__),
    .I1(g116),
    .I0(g114),
    .O(__3103__)
  );
  LUT5 #(
    .INIT(32'h7fff0000)
  ) __6484__ (
    .I4(__747__),
    .I3(g35),
    .I2(__1240__),
    .I1(__1567__),
    .I0(__1696__),
    .O(__3104__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __6485__ (
    .I1(__544__),
    .I0(__646__),
    .O(__3105__)
  );
  LUT6 #(
    .INIT(64'hff004c80f0f0f0f0)
  ) __6486__ (
    .I5(g35),
    .I4(__3105__),
    .I3(__1105__),
    .I2(__775__),
    .I1(__1813__),
    .I0(__1036__),
    .O(__3106__)
  );
  LUT6 #(
    .INIT(64'hff00df10ffff0000)
  ) __6487__ (
    .I5(g35),
    .I4(__569__),
    .I3(__598__),
    .I2(__1794__),
    .I1(__313__),
    .I0(__1391__),
    .O(__3107__)
  );
  LUT6 #(
    .INIT(64'h06666666aaaaaaaa)
  ) __6488__ (
    .I5(g35),
    .I4(__1303__),
    .I3(__810__),
    .I2(__1294__),
    .I1(__463__),
    .I0(__120__),
    .O(__3108__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6489__ (
    .I5(g35),
    .I4(__2952__),
    .I3(__1946__),
    .I2(__274__),
    .I1(__853__),
    .I0(__1391__),
    .O(__3109__)
  );
  LUT4 #(
    .INIT(16'h7f00)
  ) __6490__ (
    .I3(__1258__),
    .I2(g35),
    .I1(__847__),
    .I0(__1594__),
    .O(__3110__)
  );
  LUT6 #(
    .INIT(64'h3fffc000aaaaaaaa)
  ) __6491__ (
    .I5(g35),
    .I4(__395__),
    .I3(__56__),
    .I2(__635__),
    .I1(__1491__),
    .I0(__59__),
    .O(__3111__)
  );
  LUT6 #(
    .INIT(64'haaaaaaaccccccccc)
  ) __6492__ (
    .I5(g35),
    .I4(__860__),
    .I3(__1111__),
    .I2(__1782__),
    .I1(__743__),
    .I0(__562__),
    .O(__3112__)
  );
  LUT6 #(
    .INIT(64'h0fff7f0070ff0000)
  ) __6493__ (
    .I5(__527__),
    .I4(__254__),
    .I3(g35),
    .I2(__1630__),
    .I1(__1338__),
    .I0(__1569__),
    .O(__3113__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __6494__ (
    .I1(__198__),
    .I0(__410__),
    .O(__3114__)
  );
  LUT6 #(
    .INIT(64'h6996966996696996)
  ) __6495__ (
    .I5(__22__),
    .I4(__501__),
    .I3(__439__),
    .I2(__34__),
    .I1(__149__),
    .I0(__3114__),
    .O(__3115__)
  );
  LUT4 #(
    .INIT(16'hb400)
  ) __6496__ (
    .I3(g35),
    .I2(__3115__),
    .I1(__781__),
    .I0(__1532__),
    .O(__3116__)
  );
  LUT5 #(
    .INIT(32'hccaaf0f0)
  ) __6497__ (
    .I4(g35),
    .I3(__1864__),
    .I2(__149__),
    .I1(__80__),
    .I0(__439__),
    .O(__3117__)
  );
  LUT6 #(
    .INIT(64'h45aa45aaffff0000)
  ) __6498__ (
    .I5(g35),
    .I4(__525__),
    .I3(__1078__),
    .I2(__973__),
    .I1(__279__),
    .I0(__1819__),
    .O(__3118__)
  );
  LUT4 #(
    .INIT(16'h7580)
  ) __6499__ (
    .I3(__614__),
    .I2(__752__),
    .I1(__1190__),
    .I0(g35),
    .O(__3119__)
  );
  LUT5 #(
    .INIT(32'h73bbc000)
  ) __6500__ (
    .I4(__564__),
    .I3(__592__),
    .I2(__1147__),
    .I1(g35),
    .I0(__2587__),
    .O(__3120__)
  );
  LUT4 #(
    .INIT(16'h44f0)
  ) __6501__ (
    .I3(g35),
    .I2(__752__),
    .I1(__665__),
    .I0(__1082__),
    .O(__3121__)
  );
  LUT2 #(
    .INIT(4'hb)
  ) __6502__ (
    .I1(__680__),
    .I0(__2121__),
    .O(__3122__)
  );
  LUT6 #(
    .INIT(64'h3fffc000aaaaaaaa)
  ) __6503__ (
    .I5(g35),
    .I4(__816__),
    .I3(__723__),
    .I2(__518__),
    .I1(__1684__),
    .I0(__416__),
    .O(__3123__)
  );
  LUT6 #(
    .INIT(64'h0000000000000008)
  ) __6504__ (
    .I5(g113),
    .I4(__1283__),
    .I3(__779__),
    .I2(__639__),
    .I1(__1483__),
    .I0(__1598__),
    .O(__3124__)
  );
  LUT6 #(
    .INIT(64'h0ff0aaaacccccccc)
  ) __6505__ (
    .I5(g35),
    .I4(__3124__),
    .I3(__1060__),
    .I2(__1407__),
    .I1(__296__),
    .I0(__228__),
    .O(__3125__)
  );
  LUT6 #(
    .INIT(64'hf055f0f0cccccccc)
  ) __6506__ (
    .I5(g35),
    .I4(__2641__),
    .I3(__746__),
    .I2(__988__),
    .I1(__358__),
    .I0(__1552__),
    .O(__3126__)
  );
  LUT4 #(
    .INIT(16'hbbf0)
  ) __6507__ (
    .I3(g35),
    .I2(__1118__),
    .I1(__99__),
    .I0(__428__),
    .O(__3127__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6508__ (
    .I1(g35),
    .I0(__219__),
    .O(__3128__)
  );
  LUT5 #(
    .INIT(32'h7df05500)
  ) __6509__ (
    .I4(__1549__),
    .I3(__265__),
    .I2(__695__),
    .I1(__1451__),
    .I0(g35),
    .O(__3129__)
  );
  LUT6 #(
    .INIT(64'hc94ccccccccccccc)
  ) __6510__ (
    .I5(g35),
    .I4(__1399__),
    .I3(__631__),
    .I2(__299__),
    .I1(__736__),
    .I0(__90__),
    .O(__3130__)
  );
  LUT4 #(
    .INIT(16'h1f30)
  ) __6511__ (
    .I3(__62__),
    .I2(g35),
    .I1(__1261__),
    .I0(__1306__),
    .O(__3131__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6512__ (
    .I5(g35),
    .I4(__2264__),
    .I3(__2158__),
    .I2(__326__),
    .I1(__879__),
    .I0(__1391__),
    .O(__3132__)
  );
  LUT5 #(
    .INIT(32'hacaacccc)
  ) __6513__ (
    .I4(g35),
    .I3(__1531__),
    .I2(__1476__),
    .I1(__1013__),
    .I0(__584__),
    .O(__3133__)
  );
  LUT4 #(
    .INIT(16'h7f00)
  ) __6514__ (
    .I3(__741__),
    .I2(g35),
    .I1(__840__),
    .I0(__2012__),
    .O(__3134__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6515__ (
    .I5(g35),
    .I4(__2952__),
    .I3(__1728__),
    .I2(__1166__),
    .I1(__686__),
    .I0(__1391__),
    .O(__3135__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6516__ (
    .I2(g35),
    .I1(__1035__),
    .I0(__1153__),
    .O(__3136__)
  );
  LUT4 #(
    .INIT(16'h7da0)
  ) __6517__ (
    .I3(__206__),
    .I2(__952__),
    .I1(__878__),
    .I0(g35),
    .O(__3137__)
  );
  LUT5 #(
    .INIT(32'habff5400)
  ) __6518__ (
    .I4(__583__),
    .I3(__1041__),
    .I2(__1207__),
    .I1(__936__),
    .I0(__983__),
    .O(__3138__)
  );
  LUT6 #(
    .INIT(64'hfa00f0f0cccccccc)
  ) __6519__ (
    .I5(g35),
    .I4(__1883__),
    .I3(__3138__),
    .I2(__275__),
    .I1(__334__),
    .I0(__2367__),
    .O(__3139__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6520__ (
    .I2(g35),
    .I1(__232__),
    .I0(__415__),
    .O(__3140__)
  );
  LUT6 #(
    .INIT(64'heaaa2aaaffff0000)
  ) __6521__ (
    .I5(g35),
    .I4(__1134__),
    .I3(__1164__),
    .I2(__964__),
    .I1(__1383__),
    .I0(__131__),
    .O(__3141__)
  );
  LUT5 #(
    .INIT(32'h10ff0000)
  ) __6522__ (
    .I4(__357__),
    .I3(g35),
    .I2(__613__),
    .I1(__623__),
    .I0(__2877__),
    .O(__3142__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __6523__ (
    .I2(__795__),
    .I1(__718__),
    .I0(__465__),
    .O(__3143__)
  );
  LUT5 #(
    .INIT(32'h78ccffcc)
  ) __6524__ (
    .I4(__650__),
    .I3(g35),
    .I2(__1227__),
    .I1(__842__),
    .I0(__3143__),
    .O(__3144__)
  );
  LUT6 #(
    .INIT(64'h50ffaaff3000cc00)
  ) __6525__ (
    .I5(__1193__),
    .I4(__246__),
    .I3(g35),
    .I2(__2866__),
    .I1(__2867__),
    .I0(__2868__),
    .O(__3145__)
  );
  LUT6 #(
    .INIT(64'h0000000000000004)
  ) __6526__ (
    .I5(__640__),
    .I4(__1441__),
    .I3(__1876__),
    .I2(__678__),
    .I1(g35),
    .I0(__747__),
    .O(__3146__)
  );
  LUT5 #(
    .INIT(32'habff5400)
  ) __6527__ (
    .I4(__245__),
    .I3(__1041__),
    .I2(__1207__),
    .I1(__936__),
    .I0(__983__),
    .O(__3147__)
  );
  LUT6 #(
    .INIT(64'hfa00f0f0cccccccc)
  ) __6528__ (
    .I5(g35),
    .I4(__1694__),
    .I3(__3147__),
    .I2(__731__),
    .I1(__583__),
    .I0(__2367__),
    .O(__3148__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6529__ (
    .I5(g35),
    .I4(__2448__),
    .I3(__2163__),
    .I2(__647__),
    .I1(__176__),
    .I0(__1391__),
    .O(__3149__)
  );
  LUT6 #(
    .INIT(64'haaaaaaaccccccccc)
  ) __6530__ (
    .I5(g35),
    .I4(__950__),
    .I3(__645__),
    .I2(__1473__),
    .I1(__102__),
    .I0(__146__),
    .O(__3150__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6531__ (
    .I1(g35),
    .I0(g6745),
    .O(__3151__)
  );
  LUT6 #(
    .INIT(64'h000000000000bf00)
  ) __6532__ (
    .I5(__1145__),
    .I4(__798__),
    .I3(g35),
    .I2(__1303__),
    .I1(__1302__),
    .I0(__810__),
    .O(__3152__)
  );
  LUT6 #(
    .INIT(64'hefefff00ff00ff00)
  ) __6533__ (
    .I5(g35),
    .I4(__341__),
    .I3(__438__),
    .I2(g72),
    .I1(g73),
    .I0(__824__),
    .O(__3153__)
  );
  LUT4 #(
    .INIT(16'hca00)
  ) __6534__ (
    .I3(g35),
    .I2(__1477__),
    .I1(__1046__),
    .I0(__939__),
    .O(__3154__)
  );
  LUT6 #(
    .INIT(64'hc0c0c0cd00000000)
  ) __6535__ (
    .I5(g35),
    .I4(__746__),
    .I3(__2601__),
    .I2(__1555__),
    .I1(__793__),
    .I0(__352__),
    .O(__3155__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __6536__ (
    .I2(g35),
    .I1(__1247__),
    .I0(__166__),
    .O(__3156__)
  );
  LUT6 #(
    .INIT(64'h23af8c00ff00ff00)
  ) __6537__ (
    .I5(g35),
    .I4(__633__),
    .I3(__587__),
    .I2(__973__),
    .I1(__1816__),
    .I0(__279__),
    .O(__3157__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6538__ (
    .I5(g35),
    .I4(__2839__),
    .I3(__1712__),
    .I2(__841__),
    .I1(__1096__),
    .I0(__1391__),
    .O(__3158__)
  );
  LUT4 #(
    .INIT(16'heef0)
  ) __6539__ (
    .I3(g35),
    .I2(__662__),
    .I1(__888__),
    .I0(__200__),
    .O(__3159__)
  );
  LUT5 #(
    .INIT(32'hcaccffff)
  ) __6540__ (
    .I4(g35),
    .I3(__913__),
    .I2(__100__),
    .I1(__1257__),
    .I0(g113),
    .O(__3160__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6541__ (
    .I5(g35),
    .I4(__1028__),
    .I3(__2023__),
    .I2(__1050__),
    .I1(__922__),
    .I0(__1980__),
    .O(__3161__)
  );
  LUT5 #(
    .INIT(32'hbf80aaaa)
  ) __6542__ (
    .I4(g35),
    .I3(__339__),
    .I2(__1674__),
    .I1(__1673__),
    .I0(__1175__),
    .O(__3162__)
  );
  LUT5 #(
    .INIT(32'hccaaf0f0)
  ) __6543__ (
    .I4(g35),
    .I3(__1531__),
    .I2(__127__),
    .I1(__198__),
    .I0(__627__),
    .O(__3163__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6544__ (
    .I2(__696__),
    .I1(__18__),
    .I0(__261__),
    .O(__3164__)
  );
  LUT6 #(
    .INIT(64'hebaa00aa00000000)
  ) __6545__ (
    .I5(g35),
    .I4(__2967__),
    .I3(__1311__),
    .I2(__557__),
    .I1(__3164__),
    .I0(__572__),
    .O(__3165__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6546__ (
    .I2(g35),
    .I1(__785__),
    .I0(__1099__),
    .O(__3166__)
  );
  LUT6 #(
    .INIT(64'hc94ccccccccccccc)
  ) __6547__ (
    .I5(g35),
    .I4(__2187__),
    .I3(__544__),
    .I2(__396__),
    .I1(__646__),
    .I0(__262__),
    .O(__3167__)
  );
  LUT6 #(
    .INIT(64'hff3fffc0aaaaaaaa)
  ) __6548__ (
    .I5(g35),
    .I4(__702__),
    .I3(__1776__),
    .I2(__1268__),
    .I1(__2861__),
    .I0(__10__),
    .O(__3168__)
  );
  LUT4 #(
    .INIT(16'h8000)
  ) __6549__ (
    .I3(__972__),
    .I2(__1503__),
    .I1(__1718__),
    .I0(__1298__),
    .O(__3169__)
  );
  LUT6 #(
    .INIT(64'hf30caaaaf0f0f0f0)
  ) __6550__ (
    .I5(g35),
    .I4(__3169__),
    .I3(__749__),
    .I2(__91__),
    .I1(__13__),
    .I0(__792__),
    .O(__3170__)
  );
  LUT6 #(
    .INIT(64'hcf0f33ff0fafff55)
  ) __6551__ (
    .I5(__1205__),
    .I4(__1070__),
    .I3(__838__),
    .I2(__2866__),
    .I1(__959__),
    .I0(__492__),
    .O(__3171__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __6552__ (
    .I2(g35),
    .I1(__3171__),
    .I0(__838__),
    .O(__3172__)
  );
  LUT5 #(
    .INIT(32'h00000080)
  ) __6553__ (
    .I4(__1110__),
    .I3(__596__),
    .I2(__762__),
    .I1(__1251__),
    .I0(__639__),
    .O(__3173__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __6554__ (
    .I1(__599__),
    .I0(__461__),
    .O(__3174__)
  );
  LUT6 #(
    .INIT(64'hdddfececf0f0f0f0)
  ) __6555__ (
    .I5(g35),
    .I4(__1030__),
    .I3(__456__),
    .I2(__845__),
    .I1(__3174__),
    .I0(__3173__),
    .O(__3175__)
  );
  LUT6 #(
    .INIT(64'hff00df10ffff0000)
  ) __6556__ (
    .I5(g35),
    .I4(__468__),
    .I3(__826__),
    .I2(__2806__),
    .I1(__704__),
    .I0(__1391__),
    .O(__3176__)
  );
  LUT4 #(
    .INIT(16'h7f00)
  ) __6557__ (
    .I3(__865__),
    .I2(g35),
    .I1(__1187__),
    .I0(__1885__),
    .O(__3177__)
  );
  LUT4 #(
    .INIT(16'h11f0)
  ) __6558__ (
    .I3(g35),
    .I2(__1247__),
    .I1(__14__),
    .I0(__772__),
    .O(__3178__)
  );
  LUT4 #(
    .INIT(16'h3caa)
  ) __6559__ (
    .I3(g35),
    .I2(__1089__),
    .I1(__1897__),
    .I0(__368__),
    .O(__3179__)
  );
  LUT6 #(
    .INIT(64'haaaaaaaccccccccc)
  ) __6560__ (
    .I5(g35),
    .I4(__728__),
    .I3(__1348__),
    .I2(__801__),
    .I1(__1119__),
    .I0(__360__),
    .O(__3180__)
  );
  LUT5 #(
    .INIT(32'hccaaf0f0)
  ) __6561__ (
    .I4(g35),
    .I3(__1451__),
    .I2(__237__),
    .I1(__1648__),
    .I0(__1183__),
    .O(__3181__)
  );
  LUT6 #(
    .INIT(64'heaaa2aaaffff0000)
  ) __6562__ (
    .I5(g35),
    .I4(__76__),
    .I3(__468__),
    .I2(__704__),
    .I1(__898__),
    .I0(__195__),
    .O(__3182__)
  );
  LUT6 #(
    .INIT(64'h7f80f0f0fffff0f0)
  ) __6563__ (
    .I5(__752__),
    .I4(g35),
    .I3(__519__),
    .I2(__1224__),
    .I1(__1190__),
    .I0(__614__),
    .O(__3183__)
  );
  LUT6 #(
    .INIT(64'h5adaaa2affff0000)
  ) __6564__ (
    .I5(g35),
    .I4(__295__),
    .I3(__1197__),
    .I2(__1299__),
    .I1(__760__),
    .I0(__692__),
    .O(__3184__)
  );
  LUT6 #(
    .INIT(64'h0fff7f0070ff0000)
  ) __6565__ (
    .I5(__870__),
    .I4(__648__),
    .I3(g35),
    .I2(__1896__),
    .I1(__1338__),
    .I0(__1568__),
    .O(__3185__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6566__ (
    .I2(g35),
    .I1(__62__),
    .I0(__435__),
    .O(__3186__)
  );
  LUT5 #(
    .INIT(32'hff44f0f0)
  ) __6567__ (
    .I4(g35),
    .I3(__2299__),
    .I2(__740__),
    .I1(__250__),
    .I0(__1678__),
    .O(__3187__)
  );
  LUT6 #(
    .INIT(64'h55df557500aa0000)
  ) __6568__ (
    .I5(__776__),
    .I4(__269__),
    .I3(__544__),
    .I2(__1147__),
    .I1(__1700__),
    .I0(g35),
    .O(__3188__)
  );
  LUT5 #(
    .INIT(32'hbf80aaaa)
  ) __6569__ (
    .I4(g35),
    .I3(__523__),
    .I2(__2557__),
    .I1(__1438__),
    .I0(__872__),
    .O(__3189__)
  );
  LUT6 #(
    .INIT(64'h3fffc000aaaaaaaa)
  ) __6570__ (
    .I5(g35),
    .I4(__434__),
    .I3(__468__),
    .I2(__704__),
    .I1(__898__),
    .I0(__1081__),
    .O(__3190__)
  );
  LUT5 #(
    .INIT(32'hccaaf0f0)
  ) __6571__ (
    .I4(g35),
    .I3(__1864__),
    .I2(__22__),
    .I1(__48__),
    .I0(__501__),
    .O(__3191__)
  );
  LUT5 #(
    .INIT(32'hc3aaf0f0)
  ) __6572__ (
    .I4(g35),
    .I3(__1936__),
    .I2(__139__),
    .I1(__454__),
    .I0(__183__),
    .O(__3192__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6573__ (
    .I2(g35),
    .I1(__1170__),
    .I0(__884__),
    .O(__3193__)
  );
  LUT6 #(
    .INIT(64'hffff44f400f000f0)
  ) __6574__ (
    .I5(__1389__),
    .I4(__607__),
    .I3(g35),
    .I2(__1101__),
    .I1(__1388__),
    .I0(__1080__),
    .O(__3194__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6575__ (
    .I5(g35),
    .I4(__1880__),
    .I3(__2451__),
    .I2(__354__),
    .I1(__212__),
    .I0(__1391__),
    .O(__3195__)
  );
  LUT6 #(
    .INIT(64'heaaa2aaaffff0000)
  ) __6576__ (
    .I5(g35),
    .I4(__220__),
    .I3(__412__),
    .I2(__900__),
    .I1(__817__),
    .I0(__375__),
    .O(__3196__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6577__ (
    .I5(g35),
    .I4(__2451__),
    .I3(__1633__),
    .I2(__212__),
    .I1(__136__),
    .I0(__1391__),
    .O(__3197__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6578__ (
    .I5(g35),
    .I4(__1969__),
    .I3(__1558__),
    .I2(__531__),
    .I1(__286__),
    .I0(__1391__),
    .O(__3198__)
  );
  LUT6 #(
    .INIT(64'hccccf0aaf0f0f0f0)
  ) __6579__ (
    .I5(g35),
    .I4(__1609__),
    .I3(__2592__),
    .I2(__906__),
    .I1(__515__),
    .I0(__409__),
    .O(__3199__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6580__ (
    .I1(__760__),
    .I0(__431__),
    .O(__3200__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __6581__ (
    .I1(__922__),
    .I0(__760__),
    .O(__3201__)
  );
  LUT6 #(
    .INIT(64'hffccff00f0f0fafa)
  ) __6582__ (
    .I5(__1197__),
    .I4(__541__),
    .I3(__3201__),
    .I2(__3200__),
    .I1(__800__),
    .I0(__1050__),
    .O(__3202__)
  );
  LUT5 #(
    .INIT(32'h0f05030f)
  ) __6583__ (
    .I4(__541__),
    .I3(__760__),
    .I2(__3202__),
    .I1(__411__),
    .I0(__64__),
    .O(__3203__)
  );
  LUT5 #(
    .INIT(32'h33aaf0f0)
  ) __6584__ (
    .I4(g35),
    .I3(__1299__),
    .I2(__541__),
    .I1(__3203__),
    .I0(__295__),
    .O(__3204__)
  );
  LUT6 #(
    .INIT(64'h50ffaaff3000cc00)
  ) __6585__ (
    .I5(__1205__),
    .I4(__838__),
    .I3(g35),
    .I2(__2866__),
    .I1(__492__),
    .I0(__959__),
    .O(__3205__)
  );
  LUT4 #(
    .INIT(16'h44f0)
  ) __6586__ (
    .I3(g35),
    .I2(__650__),
    .I1(__85__),
    .I0(__551__),
    .O(__3206__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6587__ (
    .I5(g35),
    .I4(__2839__),
    .I3(__2061__),
    .I2(__283__),
    .I1(__841__),
    .I0(__1391__),
    .O(__3207__)
  );
  LUT5 #(
    .INIT(32'hecffea00)
  ) __6588__ (
    .I4(__448__),
    .I3(g35),
    .I2(__1142__),
    .I1(__384__),
    .I0(__550__),
    .O(__3208__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6589__ (
    .I5(g35),
    .I4(__2027__),
    .I3(__2266__),
    .I2(__95__),
    .I1(__29__),
    .I0(__1391__),
    .O(__3209__)
  );
  LUT5 #(
    .INIT(32'h5f3f0000)
  ) __6590__ (
    .I4(__588__),
    .I3(__734__),
    .I2(g35),
    .I1(__1003__),
    .I0(__1011__),
    .O(__3210__)
  );
  LUT4 #(
    .INIT(16'h1f30)
  ) __6591__ (
    .I3(__847__),
    .I2(g35),
    .I1(__1156__),
    .I0(__1594__),
    .O(__3211__)
  );
  LUT6 #(
    .INIT(64'hc0c0c0cd00000000)
  ) __6592__ (
    .I5(g35),
    .I4(__196__),
    .I3(__1484__),
    .I2(__1489__),
    .I1(__1028__),
    .I0(__190__),
    .O(__3212__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6593__ (
    .I2(g35),
    .I1(g6748),
    .I0(__1087__),
    .O(__3213__)
  );
  LUT3 #(
    .INIT(8'h08)
  ) __6594__ (
    .I2(__881__),
    .I1(__660__),
    .I0(__580__),
    .O(__3214__)
  );
  LUT6 #(
    .INIT(64'hdfff7555aaaa0000)
  ) __6595__ (
    .I5(__1243__),
    .I4(__500__),
    .I3(__3214__),
    .I2(__152__),
    .I1(__985__),
    .I0(g35),
    .O(__3215__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __6596__ (
    .I1(__728__),
    .I0(__1348__),
    .O(__3216__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6597__ (
    .I5(g35),
    .I4(__179__),
    .I3(__3216__),
    .I2(__763__),
    .I1(__506__),
    .I0(__1344__),
    .O(__3217__)
  );
  LUT3 #(
    .INIT(8'hd0)
  ) __6598__ (
    .I2(__1003__),
    .I1(__1011__),
    .I0(g35),
    .O(__3218__)
  );
  LUT5 #(
    .INIT(32'h7fd5aa00)
  ) __6599__ (
    .I4(__652__),
    .I3(__166__),
    .I2(__585__),
    .I1(__1068__),
    .I0(g35),
    .O(__3219__)
  );
  LUT5 #(
    .INIT(32'h3caaf0f0)
  ) __6600__ (
    .I4(g35),
    .I3(__2779__),
    .I2(__609__),
    .I1(__195__),
    .I0(__1081__),
    .O(__3220__)
  );
  LUT5 #(
    .INIT(32'habff5400)
  ) __6601__ (
    .I4(__943__),
    .I3(__1115__),
    .I2(__35__),
    .I1(__437__),
    .I0(__667__),
    .O(__3221__)
  );
  LUT6 #(
    .INIT(64'hfa00f0f0cccccccc)
  ) __6602__ (
    .I5(g35),
    .I4(__1759__),
    .I3(__3221__),
    .I2(__137__),
    .I1(__710__),
    .I0(__1497__),
    .O(__3222__)
  );
  LUT5 #(
    .INIT(32'h00cef0f0)
  ) __6603__ (
    .I4(g35),
    .I3(__401__),
    .I2(__1106__),
    .I1(__492__),
    .I0(__559__),
    .O(__3223__)
  );
  LUT6 #(
    .INIT(64'heeeef0f0ff00ff00)
  ) __6604__ (
    .I5(g35),
    .I4(__1383__),
    .I3(__984__),
    .I2(__1164__),
    .I1(__2268__),
    .I0(__1114__),
    .O(__3224__)
  );
  LUT6 #(
    .INIT(64'hf055f0f0cccccccc)
  ) __6605__ (
    .I5(g35),
    .I4(__2965__),
    .I3(__112__),
    .I2(__608__),
    .I1(__26__),
    .I0(__1827__),
    .O(__3225__)
  );
  LUT3 #(
    .INIT(8'h78)
  ) __6606__ (
    .I2(__734__),
    .I1(g35),
    .I0(__725__),
    .O(__3226__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6607__ (
    .I1(g35),
    .I0(__954__),
    .O(__3227__)
  );
  LUT5 #(
    .INIT(32'h0af0cccc)
  ) __6608__ (
    .I4(g35),
    .I3(__2616__),
    .I2(__331__),
    .I1(__1275__),
    .I0(__1207__),
    .O(__3228__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6609__ (
    .I5(g35),
    .I4(__2000__),
    .I3(__1621__),
    .I2(__475__),
    .I1(__1042__),
    .I0(__1391__),
    .O(__3229__)
  );
  LUT5 #(
    .INIT(32'h33aaf0f0)
  ) __6610__ (
    .I4(g35),
    .I3(__2935__),
    .I2(__273__),
    .I1(__2034__),
    .I0(__7__),
    .O(__3230__)
  );
  LUT5 #(
    .INIT(32'h575d0a00)
  ) __6611__ (
    .I4(__1067__),
    .I3(__498__),
    .I2(__2190__),
    .I1(__2191__),
    .I0(g35),
    .O(__3231__)
  );
  LUT6 #(
    .INIT(64'hee22eeeef0f0f0f0)
  ) __6612__ (
    .I5(g35),
    .I4(__1248__),
    .I3(__1245__),
    .I2(__404__),
    .I1(__2057__),
    .I0(__1278__),
    .O(__3232__)
  );
  LUT6 #(
    .INIT(64'h7fd55555aa000000)
  ) __6613__ (
    .I5(__445__),
    .I4(__752__),
    .I3(__810__),
    .I2(__519__),
    .I1(__2770__),
    .I0(g35),
    .O(__3233__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6614__ (
    .I5(g35),
    .I4(__1625__),
    .I3(__2690__),
    .I2(__852__),
    .I1(__67__),
    .I0(__1391__),
    .O(__3234__)
  );
  LUT6 #(
    .INIT(64'h2aaad55500000000)
  ) __6615__ (
    .I5(g35),
    .I4(__1391__),
    .I3(__457__),
    .I2(__874__),
    .I1(__1264__),
    .I0(__110__),
    .O(__3235__)
  );
  LUT4 #(
    .INIT(16'hbbf0)
  ) __6616__ (
    .I3(g35),
    .I2(__441__),
    .I1(__1018__),
    .I0(__224__),
    .O(__3236__)
  );
  LUT4 #(
    .INIT(16'hbbf0)
  ) __6617__ (
    .I3(g35),
    .I2(__1250__),
    .I1(__941__),
    .I0(__340__),
    .O(__3237__)
  );
  LUT5 #(
    .INIT(32'hc3aaf0f0)
  ) __6618__ (
    .I4(g35),
    .I3(__1528__),
    .I2(__1198__),
    .I1(__60__),
    .I0(__1076__),
    .O(__3238__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6619__ (
    .I5(g35),
    .I4(__2184__),
    .I3(__2543__),
    .I2(__172__),
    .I1(__37__),
    .I0(__1391__),
    .O(__3239__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6620__ (
    .I2(g35),
    .I1(__221__),
    .I0(__340__),
    .O(__3240__)
  );
  LUT4 #(
    .INIT(16'h0777)
  ) __6621__ (
    .I3(__1200__),
    .I2(__345__),
    .I1(__1153__),
    .I0(__44__),
    .O(__3241__)
  );
  LUT6 #(
    .INIT(64'h0000077707770777)
  ) __6622__ (
    .I5(__1159__),
    .I4(__388__),
    .I3(__291__),
    .I2(__694__),
    .I1(__1035__),
    .I0(__264__),
    .O(__3242__)
  );
  LUT6 #(
    .INIT(64'h153f000000000000)
  ) __6623__ (
    .I5(__3242__),
    .I4(__3241__),
    .I3(__40__),
    .I2(__209__),
    .I1(__1260__),
    .I0(__773__),
    .O(__3243__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6624__ (
    .I2(__2331__),
    .I1(__446__),
    .I0(__942__),
    .O(__3244__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6625__ (
    .I1(g35),
    .I0(__494__),
    .O(__3245__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6626__ (
    .I5(g35),
    .I4(__2184__),
    .I3(__1692__),
    .I2(__1132__),
    .I1(__715__),
    .I0(__1391__),
    .O(__3246__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6627__ (
    .I5(g35),
    .I4(__1866__),
    .I3(__2806__),
    .I2(__677__),
    .I1(__699__),
    .I0(__1391__),
    .O(__3247__)
  );
  LUT6 #(
    .INIT(64'h7f80f0f0fffff0f0)
  ) __6628__ (
    .I5(__752__),
    .I4(g35),
    .I3(__664__),
    .I2(__629__),
    .I1(__605__),
    .I0(__2006__),
    .O(__3248__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6629__ (
    .I5(g35),
    .I4(__1394__),
    .I3(__2690__),
    .I2(__86__),
    .I1(__1007__),
    .I0(__1391__),
    .O(__3249__)
  );
  LUT4 #(
    .INIT(16'h7da0)
  ) __6630__ (
    .I3(__1110__),
    .I2(__1251__),
    .I1(__762__),
    .I0(g35),
    .O(__3250__)
  );
  LUT5 #(
    .INIT(32'h7d55a000)
  ) __6631__ (
    .I4(__482__),
    .I3(__1432__),
    .I2(__1268__),
    .I1(__794__),
    .I0(g35),
    .O(__3251__)
  );
  LUT5 #(
    .INIT(32'hff44f0f0)
  ) __6632__ (
    .I4(g35),
    .I3(__2637__),
    .I2(__1212__),
    .I1(__733__),
    .I0(__1630__),
    .O(__3252__)
  );
  LUT6 #(
    .INIT(64'hbfff0000bfffbfff)
  ) __6633__ (
    .I5(__758__),
    .I4(__875__),
    .I3(__265__),
    .I2(__403__),
    .I1(__1125__),
    .I0(__671__),
    .O(__3253__)
  );
  LUT6 #(
    .INIT(64'h4cccffccf0f0f0f0)
  ) __6634__ (
    .I5(g35),
    .I4(__3253__),
    .I3(__1451__),
    .I2(__671__),
    .I1(__758__),
    .I0(__177__),
    .O(__3254__)
  );
  LUT5 #(
    .INIT(32'hc3aaf0f0)
  ) __6635__ (
    .I4(g35),
    .I3(__2056__),
    .I2(__375__),
    .I1(__220__),
    .I0(__455__),
    .O(__3255__)
  );
  LUT6 #(
    .INIT(64'hee22eeeef0f0f0f0)
  ) __6636__ (
    .I5(g35),
    .I4(__1248__),
    .I3(__1245__),
    .I2(__109__),
    .I1(__2051__),
    .I0(__1226__),
    .O(__3256__)
  );
  LUT6 #(
    .INIT(64'hf7f3ff0000000000)
  ) __6637__ (
    .I5(g35),
    .I4(__1586__),
    .I3(__53__),
    .I2(__3174__),
    .I1(__639__),
    .I0(__596__),
    .O(__3257__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6638__ (
    .I2(__511__),
    .I1(__31__),
    .I0(__865__),
    .O(__3258__)
  );
  LUT5 #(
    .INIT(32'h00000080)
  ) __6639__ (
    .I4(__282__),
    .I3(__452__),
    .I2(__132__),
    .I1(__32__),
    .I0(__347__),
    .O(__3259__)
  );
  LUT6 #(
    .INIT(64'hebaa00aa00000000)
  ) __6640__ (
    .I5(g35),
    .I4(__3259__),
    .I3(__1673__),
    .I2(__820__),
    .I1(__3258__),
    .I0(__504__),
    .O(__3260__)
  );
  LUT5 #(
    .INIT(32'hccaaf0f0)
  ) __6641__ (
    .I4(g35),
    .I3(__998__),
    .I2(__666__),
    .I1(__1147__),
    .I0(__966__),
    .O(__3261__)
  );
  LUT5 #(
    .INIT(32'h7d55a000)
  ) __6642__ (
    .I4(__203__),
    .I3(__2765__),
    .I2(__1235__),
    .I1(__706__),
    .I0(g35),
    .O(__3262__)
  );
  LUT6 #(
    .INIT(64'h3fffc000aaaaaaaa)
  ) __6643__ (
    .I5(g35),
    .I4(__102__),
    .I3(__1643__),
    .I2(__191__),
    .I1(__958__),
    .I0(__745__),
    .O(__3263__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __6644__ (
    .I1(__819__),
    .I0(__769__),
    .O(__3264__)
  );
  LUT6 #(
    .INIT(64'h3caaaaaaf0f0f0f0)
  ) __6645__ (
    .I5(g35),
    .I4(__3264__),
    .I3(__1286__),
    .I2(__1194__),
    .I1(__946__),
    .I0(__16__),
    .O(__3265__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6646__ (
    .I5(g35),
    .I4(__1880__),
    .I3(__1866__),
    .I2(__1010__),
    .I1(__377__),
    .I0(__1391__),
    .O(__3266__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6647__ (
    .I2(g35),
    .I1(__913__),
    .I0(__100__),
    .O(__3267__)
  );
  LUT6 #(
    .INIT(64'heeeef0f0ff00ff00)
  ) __6648__ (
    .I5(g35),
    .I4(__1643__),
    .I3(__141__),
    .I2(__191__),
    .I1(__2541__),
    .I0(__1208__),
    .O(__3268__)
  );
  LUT5 #(
    .INIT(32'h575d0a00)
  ) __6649__ (
    .I4(__1034__),
    .I3(__962__),
    .I2(__2940__),
    .I1(__1145__),
    .I0(g35),
    .O(__3269__)
  );
  LUT6 #(
    .INIT(64'h8000000000000000)
  ) __6650__ (
    .I5(__252__),
    .I4(__175__),
    .I3(__642__),
    .I2(__790__),
    .I1(__459__),
    .I0(__2324__),
    .O(__3270__)
  );
  LUT6 #(
    .INIT(64'h45aa45aaffff0000)
  ) __6651__ (
    .I5(g35),
    .I4(__459__),
    .I3(__525__),
    .I2(__973__),
    .I1(__279__),
    .I0(__3270__),
    .O(__3271__)
  );
  LUT5 #(
    .INIT(32'h00cef0f0)
  ) __6652__ (
    .I4(g35),
    .I3(__618__),
    .I2(__1254__),
    .I1(__435__),
    .I0(__106__),
    .O(__3272__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6653__ (
    .I5(g35),
    .I4(__2026__),
    .I3(__1791__),
    .I2(__408__),
    .I1(__953__),
    .I0(__1391__),
    .O(__3273__)
  );
  LUT6 #(
    .INIT(64'h000000000000bf00)
  ) __6654__ (
    .I5(__688__),
    .I4(__457__),
    .I3(g35),
    .I2(__1303__),
    .I1(__1294__),
    .I0(__810__),
    .O(__3274__)
  );
  LUT3 #(
    .INIT(8'h08)
  ) __6655__ (
    .I2(__546__),
    .I1(g35),
    .I0(__214__),
    .O(__3275__)
  );
  LUT5 #(
    .INIT(32'hefffffff)
  ) __6656__ (
    .I4(__680__),
    .I3(__2138__),
    .I2(__2137__),
    .I1(__2133__),
    .I0(__2128__),
    .O(__3276__)
  );
  LUT6 #(
    .INIT(64'hcfcccfcc4544cfcc)
  ) __6657__ (
    .I5(__972__),
    .I4(__1444__),
    .I3(__23__),
    .I2(__243__),
    .I1(__142__),
    .I0(__1465__),
    .O(__3277__)
  );
  LUT5 #(
    .INIT(32'h33aaf0f0)
  ) __6658__ (
    .I4(g35),
    .I3(__1430__),
    .I2(__1080__),
    .I1(__3277__),
    .I0(__243__),
    .O(__3278__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6659__ (
    .I2(g35),
    .I1(__376__),
    .I0(__362__),
    .O(__3279__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6660__ (
    .I5(g35),
    .I4(__2000__),
    .I3(__1743__),
    .I2(__1042__),
    .I1(__487__),
    .I0(__1391__),
    .O(__3280__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6661__ (
    .I5(g35),
    .I4(__1837__),
    .I3(__1625__),
    .I2(__150__),
    .I1(__1053__),
    .I0(__1391__),
    .O(__3281__)
  );
  LUT4 #(
    .INIT(16'hb000)
  ) __6662__ (
    .I3(g35),
    .I2(__786__),
    .I1(__973__),
    .I0(__279__),
    .O(__3282__)
  );
  LUT6 #(
    .INIT(64'hffff80ffffff0000)
  ) __6663__ (
    .I5(__693__),
    .I4(__3282__),
    .I3(g35),
    .I2(__1078__),
    .I1(__251__),
    .I0(__1819__),
    .O(__3283__)
  );
  LUT6 #(
    .INIT(64'haaaaaaaccccccccc)
  ) __6664__ (
    .I5(g35),
    .I4(__944__),
    .I3(__296__),
    .I2(__1600__),
    .I1(__55__),
    .I0(__946__),
    .O(__3284__)
  );
  LUT6 #(
    .INIT(64'h70f0f07000000000)
  ) __6665__ (
    .I5(g35),
    .I4(__584__),
    .I3(__77__),
    .I2(__758__),
    .I1(__1452__),
    .I0(__1449__),
    .O(__3285__)
  );
  LUT6 #(
    .INIT(64'h7fffd50055005500)
  ) __6666__ (
    .I5(__3285__),
    .I4(__916__),
    .I3(__698__),
    .I2(__1452__),
    .I1(__397__),
    .I0(g35),
    .O(__3286__)
  );
  LUT6 #(
    .INIT(64'hffff44f400f000f0)
  ) __6667__ (
    .I5(__1389__),
    .I4(__933__),
    .I3(g35),
    .I2(__851__),
    .I1(__1388__),
    .I0(__41__),
    .O(__3287__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6668__ (
    .I5(g35),
    .I4(__2952__),
    .I3(__2361__),
    .I2(__1218__),
    .I1(__156__),
    .I0(__1391__),
    .O(__3288__)
  );
  LUT6 #(
    .INIT(64'hf0f04444ff00ff00)
  ) __6669__ (
    .I5(g35),
    .I4(__1521__),
    .I3(__907__),
    .I2(__540__),
    .I1(__112__),
    .I0(__1523__),
    .O(__3289__)
  );
  LUT5 #(
    .INIT(32'h575d0a00)
  ) __6670__ (
    .I4(__313__),
    .I3(__569__),
    .I2(__1386__),
    .I1(__989__),
    .I0(g35),
    .O(__3290__)
  );
  LUT5 #(
    .INIT(32'h6ff6ff00)
  ) __6671__ (
    .I4(g35),
    .I3(__337__),
    .I2(__604__),
    .I1(__756__),
    .I0(__1031__),
    .O(__3291__)
  );
  LUT5 #(
    .INIT(32'h73bbc000)
  ) __6672__ (
    .I4(__575__),
    .I3(__510__),
    .I2(__2372__),
    .I1(g35),
    .I0(__2373__),
    .O(__3292__)
  );
  LUT6 #(
    .INIT(64'h3fc0bfc8f0f0f0f0)
  ) __6673__ (
    .I5(g35),
    .I4(__1041__),
    .I3(__507__),
    .I2(__1032__),
    .I1(__364__),
    .I0(__2189__),
    .O(__3293__)
  );
  LUT4 #(
    .INIT(16'h3caa)
  ) __6674__ (
    .I3(g35),
    .I2(__2281__),
    .I1(__220__),
    .I0(__1171__),
    .O(__3294__)
  );
  LUT6 #(
    .INIT(64'hc3aaaaaaf0f0f0f0)
  ) __6675__ (
    .I5(g35),
    .I4(__2465__),
    .I3(__2301__),
    .I2(__1093__),
    .I1(__658__),
    .I0(__971__),
    .O(__3295__)
  );
  LUT5 #(
    .INIT(32'hccaaf0f0)
  ) __6676__ (
    .I4(g35),
    .I3(__1864__),
    .I2(__198__),
    .I1(__538__),
    .I0(__1046__),
    .O(__3296__)
  );
  LUT6 #(
    .INIT(64'hccccf0aaf0f0f0f0)
  ) __6677__ (
    .I5(g35),
    .I4(__1609__),
    .I3(__3259__),
    .I2(__504__),
    .I1(__515__),
    .I0(__374__),
    .O(__3297__)
  );
  LUT6 #(
    .INIT(64'h3bcc3bcc00000000)
  ) __6678__ (
    .I5(g35),
    .I4(__507__),
    .I3(__1032__),
    .I2(__1041__),
    .I1(__364__),
    .I0(__2189__),
    .O(__3298__)
  );
  LUT3 #(
    .INIT(8'h8f)
  ) __6679__ (
    .I2(g35),
    .I1(__123__),
    .I0(__799__),
    .O(__3299__)
  );
  LUT6 #(
    .INIT(64'h505050f350f35050)
  ) __6680__ (
    .I5(__185__),
    .I4(__1351__),
    .I3(__3299__),
    .I2(__869__),
    .I1(__751__),
    .I0(g35),
    .O(__3300__)
  );
  LUT6 #(
    .INIT(64'hccccccacaaaaaaaa)
  ) __6681__ (
    .I5(g35),
    .I4(__881__),
    .I3(__660__),
    .I2(__580__),
    .I1(__985__),
    .I0(__365__),
    .O(__3301__)
  );
  LUT6 #(
    .INIT(64'h3caaaaaaf0f0f0f0)
  ) __6682__ (
    .I5(g35),
    .I4(__1674__),
    .I3(__1673__),
    .I2(__290__),
    .I1(__787__),
    .I0(__300__),
    .O(__3302__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __6683__ (
    .I1(g35),
    .I0(__684__),
    .O(__3303__)
  );
  LUT6 #(
    .INIT(64'h000c000500000000)
  ) __6684__ (
    .I5(__3303__),
    .I4(__351__),
    .I3(__1063__),
    .I2(__1123__),
    .I1(__1040__),
    .I0(__1074__),
    .O(__3304__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6685__ (
    .I1(__784__),
    .I0(__462__),
    .O(__3305__)
  );
  LUT6 #(
    .INIT(64'hc3aaaaaaf0f0f0f0)
  ) __6686__ (
    .I5(g35),
    .I4(__3305__),
    .I3(__1446__),
    .I2(__1148__),
    .I1(__931__),
    .I0(__836__),
    .O(__3306__)
  );
  LUT5 #(
    .INIT(32'h7f300000)
  ) __6687__ (
    .I4(g35),
    .I3(__365__),
    .I2(__1499__),
    .I1(__152__),
    .I0(__985__),
    .O(__3307__)
  );
  LUT3 #(
    .INIT(8'hf4)
  ) __6688__ (
    .I2(__2212__),
    .I1(__535__),
    .I0(g35),
    .O(__3308__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6689__ (
    .I1(g35),
    .I0(__242__),
    .O(__3309__)
  );
  LUT5 #(
    .INIT(32'hccaaf0f0)
  ) __6690__ (
    .I4(g35),
    .I3(__1531__),
    .I2(__700__),
    .I1(__1046__),
    .I0(__942__),
    .O(__3310__)
  );
  LUT5 #(
    .INIT(32'h7d55a000)
  ) __6691__ (
    .I4(__606__),
    .I3(__214__),
    .I2(__719__),
    .I1(__546__),
    .I0(g35),
    .O(__3311__)
  );
  LUT6 #(
    .INIT(64'h0001ffffffffffff)
  ) __6692__ (
    .I5(g35),
    .I4(__2906__),
    .I3(__844__),
    .I2(__947__),
    .I1(__1094__),
    .I0(__745__),
    .O(__3312__)
  );
  LUT4 #(
    .INIT(16'hf800)
  ) __6693__ (
    .I3(__3173__),
    .I2(__845__),
    .I1(__1030__),
    .I0(__456__),
    .O(__3313__)
  );
  LUT6 #(
    .INIT(64'h05050404ff00ff00)
  ) __6694__ (
    .I5(g35),
    .I4(__845__),
    .I3(__639__),
    .I2(__3174__),
    .I1(__3173__),
    .I0(__3313__),
    .O(__3314__)
  );
  LUT5 #(
    .INIT(32'hc3aaf0f0)
  ) __6695__ (
    .I4(g35),
    .I3(__2512__),
    .I2(__1141__),
    .I1(__1253__),
    .I0(__697__),
    .O(__3315__)
  );
  LUT6 #(
    .INIT(64'hefefff00ff00ff00)
  ) __6696__ (
    .I5(g35),
    .I4(__341__),
    .I3(__344__),
    .I2(g73),
    .I1(g72),
    .I0(__824__),
    .O(__3316__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6697__ (
    .I5(g35),
    .I4(__1969__),
    .I3(__1837__),
    .I2(__286__),
    .I1(__929__),
    .I0(__1391__),
    .O(__3317__)
  );
  LUT6 #(
    .INIT(64'h001c00ccf0f0f0f0)
  ) __6698__ (
    .I5(g35),
    .I4(__1698__),
    .I3(__1697__),
    .I2(__32__),
    .I1(__452__),
    .I0(__347__),
    .O(__3318__)
  );
  LUT6 #(
    .INIT(64'hffff44f400f000f0)
  ) __6699__ (
    .I5(__1389__),
    .I4(__993__),
    .I3(g35),
    .I2(__278__),
    .I1(__1388__),
    .I0(__737__),
    .O(__3319__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6700__ (
    .I5(g35),
    .I4(__2027__),
    .I3(__2448__),
    .I2(__79__),
    .I1(__647__),
    .I0(__1391__),
    .O(__3320__)
  );
  LUT6 #(
    .INIT(64'h000078f0aaaaaaaa)
  ) __6701__ (
    .I5(g35),
    .I4(__1776__),
    .I3(__976__),
    .I2(__871__),
    .I1(__1775__),
    .I0(__738__),
    .O(__3321__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6702__ (
    .I1(__881__),
    .I0(__660__),
    .O(__3322__)
  );
  LUT6 #(
    .INIT(64'haaf0f0f0cccccccc)
  ) __6703__ (
    .I5(g35),
    .I4(__3322__),
    .I3(__170__),
    .I2(__99__),
    .I1(__204__),
    .I0(__299__),
    .O(__3323__)
  );
  LUT5 #(
    .INIT(32'hff44f0f0)
  ) __6704__ (
    .I4(g35),
    .I3(__2568__),
    .I2(__1219__),
    .I1(__382__),
    .I0(__1438__),
    .O(__3324__)
  );
  LUT6 #(
    .INIT(64'h3fffc000aaaaaaaa)
  ) __6705__ (
    .I5(g35),
    .I4(__1043__),
    .I3(__1110__),
    .I2(__1251__),
    .I1(__547__),
    .I0(__762__),
    .O(__3325__)
  );
  LUT5 #(
    .INIT(32'h33aaf0f0)
  ) __6706__ (
    .I4(g35),
    .I3(__2487__),
    .I2(__225__),
    .I1(__1733__),
    .I0(__649__),
    .O(__3326__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6707__ (
    .I2(g35),
    .I1(__1159__),
    .I0(__1200__),
    .O(__3327__)
  );
  LUT6 #(
    .INIT(64'hefefff00ff00ff00)
  ) __6708__ (
    .I5(g35),
    .I4(__341__),
    .I3(__814__),
    .I2(g73),
    .I1(g72),
    .I0(__390__),
    .O(__3328__)
  );
  LUT6 #(
    .INIT(64'heaaa2aaaffff0000)
  ) __6709__ (
    .I5(g35),
    .I4(__1150__),
    .I3(__962__),
    .I2(__1145__),
    .I1(__1034__),
    .I0(__1037__),
    .O(__3329__)
  );
  LUT6 #(
    .INIT(64'h007f00ffffff0000)
  ) __6710__ (
    .I5(g35),
    .I4(__816__),
    .I3(__1066__),
    .I2(__723__),
    .I1(__518__),
    .I0(__1684__),
    .O(__3330__)
  );
  LUT6 #(
    .INIT(64'h2aaad55500000000)
  ) __6711__ (
    .I5(g35),
    .I4(__1391__),
    .I3(__962__),
    .I2(__1145__),
    .I1(__1034__),
    .I0(__314__),
    .O(__3331__)
  );
  LUT6 #(
    .INIT(64'h00ff33330f0f5555)
  ) __6712__ (
    .I5(g72),
    .I4(g73),
    .I3(__149__),
    .I2(__22__),
    .I1(__410__),
    .I0(__198__),
    .O(__3332__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __6713__ (
    .I2(g35),
    .I1(__3332__),
    .I0(__417__),
    .O(__3333__)
  );
  LUT5 #(
    .INIT(32'hbf80aaaa)
  ) __6714__ (
    .I4(g35),
    .I3(__1221__),
    .I2(__2288__),
    .I1(__1678__),
    .I0(__1206__),
    .O(__3334__)
  );
  LUT6 #(
    .INIT(64'h45aa45aaffff0000)
  ) __6715__ (
    .I5(g35),
    .I4(__175__),
    .I3(__252__),
    .I2(__973__),
    .I1(__279__),
    .I0(__1818__),
    .O(__3335__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __6716__ (
    .I1(__595__),
    .I0(__540__),
    .O(__3336__)
  );
  LUT6 #(
    .INIT(64'h0000000000008000)
  ) __6717__ (
    .I5(g113),
    .I4(__1283__),
    .I3(__779__),
    .I2(__1522__),
    .I1(__639__),
    .I0(__1520__),
    .O(__3337__)
  );
  LUT6 #(
    .INIT(64'h0ff0aaaacccccccc)
  ) __6718__ (
    .I5(g35),
    .I4(__3337__),
    .I3(__1060__),
    .I2(__3336__),
    .I1(__112__),
    .I0(__907__),
    .O(__3338__)
  );
  LUT6 #(
    .INIT(64'hddecffccffff0000)
  ) __6719__ (
    .I5(g35),
    .I4(__1030__),
    .I3(__456__),
    .I2(__845__),
    .I1(__3174__),
    .I0(__3173__),
    .O(__3339__)
  );
  LUT5 #(
    .INIT(32'h05f0cccc)
  ) __6720__ (
    .I4(g35),
    .I3(__1757__),
    .I2(__659__),
    .I1(__75__),
    .I0(__1144__),
    .O(__3340__)
  );
  LUT6 #(
    .INIT(64'hc3aaaaaaf0f0f0f0)
  ) __6721__ (
    .I5(g35),
    .I4(__1847__),
    .I3(__1630__),
    .I2(__258__),
    .I1(__235__),
    .I0(__903__),
    .O(__3341__)
  );
  LUT6 #(
    .INIT(64'h3fffc000aaaaaaaa)
  ) __6722__ (
    .I5(g35),
    .I4(__1223__),
    .I3(__509__),
    .I2(__306__),
    .I1(__705__),
    .I0(__20__),
    .O(__3342__)
  );
  LUT6 #(
    .INIT(64'h12121030ffff0000)
  ) __6723__ (
    .I5(g35),
    .I4(__1240__),
    .I3(__738__),
    .I2(__976__),
    .I1(__1776__),
    .I0(__1775__),
    .O(__3343__)
  );
  LUT6 #(
    .INIT(64'hff80808080808080)
  ) __6724__ (
    .I5(__1440__),
    .I4(__1876__),
    .I3(__2178__),
    .I2(__1698__),
    .I1(__1608__),
    .I0(__1396__),
    .O(__3344__)
  );
  LUT6 #(
    .INIT(64'hff07ffffffffffff)
  ) __6725__ (
    .I5(g113),
    .I4(__1567__),
    .I3(__3344__),
    .I2(g134),
    .I1(__884__),
    .I0(g99),
    .O(__3345__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __6726__ (
    .I1(__746__),
    .I0(__352__),
    .O(__3346__)
  );
  LUT5 #(
    .INIT(32'h00000008)
  ) __6727__ (
    .I4(g113),
    .I3(__1283__),
    .I2(__779__),
    .I1(__1411__),
    .I0(__1554__),
    .O(__3347__)
  );
  LUT6 #(
    .INIT(64'h0ff0aaaacccccccc)
  ) __6728__ (
    .I5(g35),
    .I4(__3347__),
    .I3(__1060__),
    .I2(__3346__),
    .I1(__793__),
    .I0(__422__),
    .O(__3348__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6729__ (
    .I2(g35),
    .I1(__65__),
    .I0(__493__),
    .O(__3349__)
  );
  LUT6 #(
    .INIT(64'hc3aaaaaaf0f0f0f0)
  ) __6730__ (
    .I5(g35),
    .I4(__2557__),
    .I3(__1438__),
    .I2(__523__),
    .I1(__872__),
    .I0(__201__),
    .O(__3350__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __6731__ (
    .I1(g35),
    .I0(__1006__),
    .O(__3351__)
  );
  LUT6 #(
    .INIT(64'h000c000500000000)
  ) __6732__ (
    .I5(__3351__),
    .I4(__901__),
    .I3(__723__),
    .I2(__644__),
    .I1(__68__),
    .I0(__518__),
    .O(__3352__)
  );
  LUT6 #(
    .INIT(64'haaaaaaaccccccccc)
  ) __6733__ (
    .I5(g35),
    .I4(__196__),
    .I3(__1028__),
    .I2(__1489__),
    .I1(__1253__),
    .I0(__1141__),
    .O(__3353__)
  );
  LUT6 #(
    .INIT(64'h80008000ffff0000)
  ) __6734__ (
    .I5(g35),
    .I4(__529__),
    .I3(__1539__),
    .I2(__210__),
    .I1(__381__),
    .I0(__333__),
    .O(__3354__)
  );
  LUT5 #(
    .INIT(32'habff5400)
  ) __6735__ (
    .I4(__500__),
    .I3(__1115__),
    .I2(__35__),
    .I1(__437__),
    .I0(__667__),
    .O(__3355__)
  );
  LUT6 #(
    .INIT(64'hcd00ccccf0f0f0f0)
  ) __6736__ (
    .I5(g35),
    .I4(__3214__),
    .I3(__3355__),
    .I2(__152__),
    .I1(__1243__),
    .I0(__365__),
    .O(__3356__)
  );
  LUT5 #(
    .INIT(32'hccaaf0f0)
  ) __6737__ (
    .I4(g35),
    .I3(__1451__),
    .I2(__996__),
    .I1(__198__),
    .I0(__657__),
    .O(__3357__)
  );
  LUT6 #(
    .INIT(64'hcaaaaaaacccccccc)
  ) __6738__ (
    .I5(g35),
    .I4(__13__),
    .I3(__711__),
    .I2(__1718__),
    .I1(__460__),
    .I0(__1140__),
    .O(__3358__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __6739__ (
    .I1(__196__),
    .I0(__190__),
    .O(__3359__)
  );
  LUT6 #(
    .INIT(64'h0000000000008000)
  ) __6740__ (
    .I5(g113),
    .I4(__1283__),
    .I3(__779__),
    .I2(__639__),
    .I1(__1488__),
    .I0(__1483__),
    .O(__3360__)
  );
  LUT6 #(
    .INIT(64'h0ff0aaaacccccccc)
  ) __6741__ (
    .I5(g35),
    .I4(__3360__),
    .I3(__1060__),
    .I2(__3359__),
    .I1(__1028__),
    .I0(__1128__),
    .O(__3361__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6742__ (
    .I2(g35),
    .I1(__508__),
    .I0(__1039__),
    .O(__3362__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6743__ (
    .I2(g35),
    .I1(__73__),
    .I0(__992__),
    .O(__3363__)
  );
  LUT5 #(
    .INIT(32'hff44f0f0)
  ) __6744__ (
    .I4(g35),
    .I3(__1477__),
    .I2(__560__),
    .I1(__1124__),
    .I0(__1451__),
    .O(__3364__)
  );
  LUT6 #(
    .INIT(64'hffff44f400f000f0)
  ) __6745__ (
    .I5(__1389__),
    .I4(__278__),
    .I3(g35),
    .I2(__611__),
    .I1(__1388__),
    .I0(__453__),
    .O(__3365__)
  );
  LUT6 #(
    .INIT(64'habffabffffff0000)
  ) __6746__ (
    .I5(g35),
    .I4(__620__),
    .I3(__1041__),
    .I2(__1207__),
    .I1(__936__),
    .I0(__216__),
    .O(__3366__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __6747__ (
    .I1(__1269__),
    .I0(__1638__),
    .O(__3367__)
  );
  LUT6 #(
    .INIT(64'hf055f0f0cccccccc)
  ) __6748__ (
    .I5(g35),
    .I4(__3367__),
    .I3(__617__),
    .I2(__1252__),
    .I1(__649__),
    .I0(__1733__),
    .O(__3368__)
  );
  LUT5 #(
    .INIT(32'h10ff0000)
  ) __6749__ (
    .I4(__267__),
    .I3(g35),
    .I2(__425__),
    .I1(__157__),
    .I0(__1894__),
    .O(__3369__)
  );
  LUT6 #(
    .INIT(64'hefffffff00000000)
  ) __6750__ (
    .I5(__640__),
    .I4(g35),
    .I3(__1440__),
    .I2(__15__),
    .I1(g113),
    .I0(__1283__),
    .O(__3370__)
  );
  LUT6 #(
    .INIT(64'h7fd55555aa000000)
  ) __6751__ (
    .I5(__1004__),
    .I4(__1147__),
    .I3(__637__),
    .I2(__914__),
    .I1(__342__),
    .I0(g35),
    .O(__3371__)
  );
  LUT6 #(
    .INIT(64'h55f0f0f0cccccccc)
  ) __6752__ (
    .I5(g35),
    .I4(__2046__),
    .I3(__1965__),
    .I2(__1262__),
    .I1(__565__),
    .I0(__1391__),
    .O(__3372__)
  );
  LUT5 #(
    .INIT(32'h7fd50000)
  ) __6753__ (
    .I4(__875__),
    .I3(__400__),
    .I2(__1451__),
    .I1(__671__),
    .I0(g35),
    .O(__3373__)
  );
  LUT6 #(
    .INIT(64'hc0c0c0cd00000000)
  ) __6754__ (
    .I5(g35),
    .I4(__1983__),
    .I3(__728__),
    .I2(__1348__),
    .I1(__801__),
    .I0(__179__),
    .O(__3374__)
  );
  LUT3 #(
    .INIT(8'h3a)
  ) __6755__ (
    .I2(g35),
    .I1(__1681__),
    .I0(__1011__),
    .O(__3375__)
  );
  LUT6 #(
    .INIT(64'heaaa2aaaffff0000)
  ) __6756__ (
    .I5(g35),
    .I4(__643__),
    .I3(__313__),
    .I2(__569__),
    .I1(__989__),
    .I0(__449__),
    .O(__3376__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6757__ (
    .I2(__1766__),
    .I1(__495__),
    .I0(__657__),
    .O(__3377__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6758__ (
    .I1(__1164__),
    .I0(__964__),
    .O(__3378__)
  );
  LUT6 #(
    .INIT(64'hc3aaaaaaf0f0f0f0)
  ) __6759__ (
    .I5(g35),
    .I4(__3378__),
    .I3(__1383__),
    .I2(__131__),
    .I1(__1134__),
    .I0(__1091__),
    .O(__3379__)
  );
  assign g20652 = __1170__;
  assign g29214 = __1170__;
  assign g16624 = __1217__;
  assign g17845 = __398__;
  assign g13881 = __520__;
  assign g33636 = __1988__;
  assign g17320 = __674__;
  assign g14673 = __991__;
  assign g16874 = __774__;
  assign g28030 = __2838__;
  assign g9680 = __74__;
  assign g12833 = __5__;
  assign g9251 = __117__;
  assign g28041 = __2820__;
  assign g21245 = __809__;
  assign g29220 = __809__;
  assign g21270 = __87__;
  assign g29217 = __87__;
  assign g11349 = __451__;
  assign g13272 = __709__;
  assign g13906 = __215__;
  assign g17604 = __833__;
  assign g12184 = __28__;
  assign g18095 = g6749;
  assign g14779 = __901__;
  assign g8291 = __712__;
  assign g17787 = __133__;
  assign g13085 = __1006__;
  assign g14694 = __1199__;
  assign g23002 = __6__;
  assign g30327 = __6__;
  assign g20763 = __218__;
  assign g29211 = __218__;
  assign g14451 = __573__;
  assign g17674 = __724__;
  assign g12350 = __612__;
  assign g10527 = __966__;
  assign g25114 = __1566__;
  assign g31860 = __1566__;
  assign g34917 = __3039__;
  assign g14147 = __330__;
  assign g34921 = __3011__;
  assign g8235 = __230__;
  assign g18099 = g6745;
  assign g8344 = __867__;
  assign g18092 = g6753;
  assign g14201 = __80__;
  assign g34927 = __2387__;
  assign g16659 = __442__;
  assign g9615 = __618__;
  assign g24162 = g54;
  assign g16722 = __1169__;
  assign g24183 = g134;
  assign g14518 = __259__;
  assign g17404 = __380__;
  assign g24185 = g44;
  assign g17400 = __1009__;
  assign g34425 = __1746__;
  assign g34839 = __1397__;
  assign g34956 = __1397__;
  assign g34923 = __3276__;
  assign g17739 = __873__;
  assign g24168 = g84;
  assign g7243 = __967__;
  assign g16656 = __217__;
  assign g16775 = __160__;
  assign g34925 = __2930__;
  assign g24181 = g126;
  assign g8784 = __305__;
  assign g24151 = 1'b1;
  assign g25582 = 1'b1;
  assign g25583 = 1'b1;
  assign g25584 = 1'b1;
  assign g25585 = 1'b1;
  assign g25586 = 1'b1;
  assign g25587 = 1'b1;
  assign g25588 = 1'b1;
  assign g25589 = 1'b1;
  assign g25590 = 1'b1;
  assign g32429 = 1'b1;
  assign g32454 = 1'b1;
  assign g33945 = 1'b1;
  assign g33946 = 1'b1;
  assign g33947 = 1'b1;
  assign g33948 = 1'b1;
  assign g33949 = 1'b1;
  assign g33950 = 1'b1;
  assign g34232 = 1'b1;
  assign g34233 = 1'b1;
  assign g34234 = 1'b1;
  assign g34235 = 1'b1;
  assign g34236 = 1'b1;
  assign g34237 = 1'b1;
  assign g34238 = 1'b1;
  assign g34239 = 1'b1;
  assign g34240 = 1'b1;
  assign g16603 = __1162__;
  assign g17813 = __811__;
  assign g13926 = __30__;
  assign g17577 = __155__;
  assign g8920 = __1202__;
  assign g21727 = __2728__;
  assign g17711 = __103__;
  assign g17649 = __723__;
  assign g19357 = __321__;
  assign g7260 = __481__;
  assign g25259 = __1948__;
  assign g31862 = __1948__;
  assign g8132 = __19__;
  assign g27831 = __1471__;
  assign g33533 = __1471__;
  assign g8786 = __1102__;
  assign g20049 = __1280__;
  assign g29210 = __1280__;
  assign g24163 = g56;
  assign g24176 = g115;
  assign g8398 = __43__;
  assign g24182 = g127;
  assign g7245 = __1103__;
  assign g24171 = g92;
  assign g24178 = g120;
  assign g12919 = __214__;
  assign g17639 = __181__;
  assign g11418 = __502__;
  assign g21176 = __954__;
  assign g29216 = __954__;
  assign g9019 = __924__;
  assign g8839 = __328__;
  assign g9741 = __189__;
  assign g16748 = __1097__;
  assign g14738 = __394__;
  assign g26876 = __1725__;
  assign g8788 = __945__;
  assign g16924 = __450__;
  assign g9555 = __106__;
  assign g33435 = __2817__;
  assign g9817 = __542__;
  assign g17715 = __105__;
  assign g20901 = __73__;
  assign g29215 = __73__;
  assign g25167 = __1801__;
  assign g31863 = __1801__;
  assign g17871 = __263__;
  assign g23683 = __739__;
  assign g30332 = __739__;
  assign g24165 = g64;
  assign g17778 = __1074__;
  assign g24177 = g116;
  assign g31521 = __2421__;
  assign g34435 = __2421__;
  assign g14662 = __474__;
  assign g32185 = __3243__;
  assign g16627 = __56__;
  assign g9048 = __751__;
  assign g18101 = g6746;
  assign g14635 = __1135__;
  assign g16955 = __433__;
  assign g16686 = __1222__;
  assign g33894 = __2469__;
  assign g34788 = __2469__;
  assign g28042 = __1468__;
  assign g8917 = __49__;
  assign g8787 = __1272__;
  assign g14217 = __994__;
  assign g10306 = __1138__;
  assign g10500 = __42__;
  assign g24179 = g124;
  assign g17291 = __484__;
  assign g17722 = __1063__;
  assign g9617 = __193__;
  assign g34201 = __2504__;
  assign g13039 = __122__;
  assign g24170 = g91;
  assign g20899 = __941__;
  assign g29212 = __941__;
  assign g13895 = __302__;
  assign g20557 = __970__;
  assign g29213 = __970__;
  assign g17423 = __998__;
  assign g9743 = __128__;
  assign g17607 = __115__;
  assign g13068 = __979__;
  assign g8719 = __547__;
  assign g17760 = __518__;
  assign g18881 = __701__;
  assign g29218 = __701__;
  assign g24175 = g114;
  assign g8916 = __521__;
  assign g14125 = __371__;
  assign g26875 = __3312__;
  assign g31656 = __2434__;
  assign g34436 = __2434__;
  assign g17819 = __349__;
  assign g13865 = __366__;
  assign g7540 = __66__;
  assign g21698 = g36;
  assign g8783 = __526__;
  assign g12923 = __1147__;
  assign g7946 = __364__;
  assign g18094 = g6748;
  assign g14189 = __419__;
  assign g21292 = __221__;
  assign g29221 = __221__;
  assign g18098 = g6744;
  assign g34972 = __2252__;
  assign g11388 = __1276__;
  assign g13049 = __1216__;
  assign g18100 = g6751;
  assign g24167 = g73;
  assign g8358 = __294__;
  assign g14749 = __887__;
  assign g11770 = __554__;
  assign g8178 = __186__;
  assign g14167 = __528__;
  assign g8342 = __1270__;
  assign g8475 = __802__;
  assign g14421 = __1038__;
  assign g8277 = __1130__;
  assign g19334 = __1085__;
  assign g34383 = __1415__;
  assign g34919 = __3072__;
  assign g17580 = __187__;
  assign g12368 = __350__;
  assign g28753 = __1896__;
  assign g33959 = __1896__;
  assign g33874 = __1619__;
  assign g17316 = __168__;
  assign g8353 = __1005__;
  assign g17685 = __644__;
  assign g16718 = __935__;
  assign g34913 = __3122__;
  assign g10122 = __14__;
  assign g8283 = __287__;
  assign g33935 = __2017__;
  assign g12832 = __1267__;
  assign g12470 = __1040__;
  assign g24174 = g113;
  assign g33079 = __1623__;
  assign g17678 = __654__;
  assign g20654 = __930__;
  assign g29219 = __930__;
  assign g14597 = __208__;
  assign g9553 = __559__;
  assign g24164 = g57;
  assign g8279 = __624__;
  assign g8416 = __1177__;
  assign g24161 = g53;
  assign g24169 = g90;
  assign g17646 = __359__;
  assign g18097 = g6747;
  assign g25219 = __847__;
  assign g31861 = __847__;
  assign g17743 = __312__;
  assign g33659 = __2060__;
  assign g24172 = g99;
  assign g31793 = __1428__;
  assign g8870 = __815__;
  assign g12238 = __379__;
  assign g12422 = __68__;
  assign g8789 = __71__;
  assign g7257 = __239__;
  assign g17764 = __72__;
  assign g13099 = __684__;
  assign g34221 = __3345__;
  assign g8785 = __813__;
  assign g16744 = __635__;
  assign g14828 = __351__;
  assign g24173 = g100;
  assign g12300 = __823__;
  assign g14705 = __98__;
  assign g8215 = __859__;
  assign g11447 = __1112__;
  assign g17519 = __759__;
  assign g8918 = __257__;
  assign g17688 = __1123__;
  assign g31665 = __2411__;
  assign g34437 = __2411__;
  assign g24180 = g125;
  assign g23759 = __2__;
  assign g30331 = __2__;
  assign g13966 = __45__;
  assign g26801 = __2051__;
  assign g32975 = __2051__;
  assign g24184 = g135;
  assign g8403 = __990__;
  assign g23652 = __3__;
  assign g30330 = __3__;
  assign g11678 = __973__;
  assign g24166 = g72;
  assign g26877 = __1844__;
  assign g9682 = __1184__;
  assign g7916 = __170__;
  assign g9497 = __401__;
  assign g13259 = __580__;
  assign g23612 = __4__;
  assign g30329 = __4__;
  assign g14096 = __48__;
  assign g34915 = __1382__;
  assign g16693 = __661__;
  assign g8915 = __1157__;
  assign g8919 = __169__;
  assign g23190 = 1'b0;
  assign g34597 = 1'b0;
  assign g18096 = g6750;
endmodule
