module s1423 (
  CK,
  G0,
  G1,
  G10,
  G11,
  G12,
  G13,
  G14,
  G15,
  G16,
  G2,
  G3,
  G4,
  G5,
  G6,
  G7,
  G8,
  G9,
  G729,
  G727,
  G702,
  G726,
  G701BF
);
  input CK;
  wire CK;
  input G0;
  wire G0;
  input G1;
  wire G1;
  input G10;
  wire G10;
  input G11;
  wire G11;
  input G12;
  wire G12;
  input G13;
  wire G13;
  input G14;
  wire G14;
  input G15;
  wire G15;
  input G16;
  wire G16;
  input G2;
  wire G2;
  input G3;
  wire G3;
  input G4;
  wire G4;
  input G5;
  wire G5;
  input G6;
  wire G6;
  input G7;
  wire G7;
  input G8;
  wire G8;
  input G9;
  wire G9;
  output G729;
  wire G729;
  output G727;
  wire G727;
  output G702;
  wire G702;
  output G726;
  wire G726;
  output G701BF;
  wire G701BF;
  wire __0__;
  wire __1__;
  wire __2__;
  wire __3__;
  wire __4__;
  wire __5__;
  wire __6__;
  wire __7__;
  wire __8__;
  wire __9__;
  wire __10__;
  wire __11__;
  wire __12__;
  wire __13__;
  wire __14__;
  wire __15__;
  wire __16__;
  wire __17__;
  wire __18__;
  wire __19__;
  wire __20__;
  wire __21__;
  wire __22__;
  wire __23__;
  wire __24__;
  wire __25__;
  wire __26__;
  wire __27__;
  wire __28__;
  wire __29__;
  wire __30__;
  wire __31__;
  wire __32__;
  wire __33__;
  wire __34__;
  wire __35__;
  wire __36__;
  wire __37__;
  wire __38__;
  wire __39__;
  wire __40__;
  wire __41__;
  wire __42__;
  wire __43__;
  wire __44__;
  wire __45__;
  wire __46__;
  wire __47__;
  wire __48__;
  wire __49__;
  wire __50__;
  wire __51__;
  wire __52__;
  wire __53__;
  wire __54__;
  wire __55__;
  wire __56__;
  wire __57__;
  wire __58__;
  wire __59__;
  wire __60__;
  wire __61__;
  wire __62__;
  wire __63__;
  wire __64__;
  wire __65__;
  wire __66__;
  wire __67__;
  wire __68__;
  wire __69__;
  wire __70__;
  wire __71__;
  wire __72__;
  wire __73__;
  wire __74__;
  wire __75__;
  wire __76__;
  wire __77__;
  wire __80__;
  wire __81__;
  wire __82__;
  wire __83__;
  wire __84__;
  wire __85__;
  wire __86__;
  wire __87__;
  wire __88__;
  wire __89__;
  wire __90__;
  wire __91__;
  wire __92__;
  wire __93__;
  wire __94__;
  wire __95__;
  wire __96__;
  wire __97__;
  wire __98__;
  wire __99__;
  wire __100__;
  wire __101__;
  wire __102__;
  wire __103__;
  wire __104__;
  wire __105__;
  wire __106__;
  wire __107__;
  wire __108__;
  wire __109__;
  wire __110__;
  wire __111__;
  wire __112__;
  wire __113__;
  wire __114__;
  wire __115__;
  wire __116__;
  wire __117__;
  wire __118__;
  wire __119__;
  wire __120__;
  wire __121__;
  wire __122__;
  wire __123__;
  wire __124__;
  wire __125__;
  wire __126__;
  wire __127__;
  wire __128__;
  wire __129__;
  wire __130__;
  wire __131__;
  wire __132__;
  wire __133__;
  wire __134__;
  wire __135__;
  wire __136__;
  wire __137__;
  wire __138__;
  wire __139__;
  wire __140__;
  wire __141__;
  wire __142__;
  wire __143__;
  wire __144__;
  wire __145__;
  wire __146__;
  wire __147__;
  wire __148__;
  wire __149__;
  wire __150__;
  wire __151__;
  wire __152__;
  wire __153__;
  wire __154__;
  wire __155__;
  wire __156__;
  wire __157__;
  wire __158__;
  wire __159__;
  wire __160__;
  wire __161__;
  wire __162__;
  wire __163__;
  wire __164__;
  wire __165__;
  wire __166__;
  wire __167__;
  wire __168__;
  wire __169__;
  wire __170__;
  wire __171__;
  wire __172__;
  wire __173__;
  wire __174__;
  wire __175__;
  wire __176__;
  wire __177__;
  wire __178__;
  wire __179__;
  wire __180__;
  wire __181__;
  wire __182__;
  wire __183__;
  wire __184__;
  wire __185__;
  wire __186__;
  wire __187__;
  wire __188__;
  wire __189__;
  wire __190__;
  wire __191__;
  wire __192__;
  wire __193__;
  wire __194__;
  wire __195__;
  wire __196__;
  wire __197__;
  wire __198__;
  wire __199__;
  wire __200__;
  wire __201__;
  wire __202__;
  wire __203__;
  wire __204__;
  wire __205__;
  INV __206__ (
    .I(G15),
    .O(__0__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __207__ (
    .D(__198__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __208__ (
    .D(__114__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__2__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __209__ (
    .D(__183__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__3__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __210__ (
    .D(__144__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__4__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __211__ (
    .D(__181__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__5__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __212__ (
    .D(__116__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__6__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __213__ (
    .D(__204__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__7__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __214__ (
    .D(__182__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__8__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __215__ (
    .D(__147__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__9__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __216__ (
    .D(__112__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__10__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __217__ (
    .D(__155__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__11__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __218__ (
    .D(__131__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__12__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __219__ (
    .D(__111__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__13__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __220__ (
    .D(__125__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__14__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __221__ (
    .D(__191__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__15__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __222__ (
    .D(__193__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__16__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __223__ (
    .D(__145__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__17__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __224__ (
    .D(__200__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__18__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __225__ (
    .D(__174__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__19__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __226__ (
    .D(__202__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__20__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __227__ (
    .D(__177__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__21__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __228__ (
    .D(__127__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__22__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __229__ (
    .D(__161__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__23__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __230__ (
    .D(__171__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__24__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __231__ (
    .D(__168__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__25__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __232__ (
    .D(__173__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__26__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __233__ (
    .D(__124__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__27__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __234__ (
    .D(__185__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__28__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __235__ (
    .D(__159__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__29__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __236__ (
    .D(__120__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__30__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __237__ (
    .D(__199__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__31__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __238__ (
    .D(__195__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__32__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __239__ (
    .D(__165__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__33__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __240__ (
    .D(__188__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__34__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __241__ (
    .D(__192__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__35__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __242__ (
    .D(__167__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__36__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __243__ (
    .D(__164__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__37__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __244__ (
    .D(__179__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__38__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __245__ (
    .D(__156__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__39__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __246__ (
    .D(__190__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__40__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __247__ (
    .D(__121__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__41__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __248__ (
    .D(__203__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__42__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __249__ (
    .D(__201__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__43__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __250__ (
    .D(__133__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__44__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __251__ (
    .D(__146__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__45__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __252__ (
    .D(__178__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__46__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __253__ (
    .D(__162__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__47__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __254__ (
    .D(__158__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__48__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __255__ (
    .D(__109__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__49__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __256__ (
    .D(__184__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__50__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __257__ (
    .D(__172__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__51__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __258__ (
    .D(__129__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__52__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __259__ (
    .D(__113__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__53__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __260__ (
    .D(__132__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__54__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __261__ (
    .D(__175__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__55__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __262__ (
    .D(__104__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__56__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __263__ (
    .D(__180__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__57__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __264__ (
    .D(__176__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__58__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __265__ (
    .D(__118__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__59__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __266__ (
    .D(__77__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__60__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __267__ (
    .D(__130__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__61__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __268__ (
    .D(__166__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__62__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __269__ (
    .D(__187__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__63__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __270__ (
    .D(__194__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__64__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __271__ (
    .D(__196__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__65__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __272__ (
    .D(__157__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__66__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __273__ (
    .D(__186__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__67__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __274__ (
    .D(__122__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__68__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __275__ (
    .D(__189__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__69__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __276__ (
    .D(__205__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__70__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __277__ (
    .D(__119__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__71__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __278__ (
    .D(__143__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__72__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __279__ (
    .D(__169__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__73__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __280__ (
    .D(__154__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__74__)
  );
  LUT4 #(
    .INIT(16'h9009)
  ) __281__ (
    .I3(__52__),
    .I2(__48__),
    .I1(__51__),
    .I0(__47__),
    .O(__75__)
  );
  LUT6 #(
    .INIT(64'h0001f00e00000000)
  ) __282__ (
    .I5(__75__),
    .I4(__49__),
    .I3(__46__),
    .I2(__50__),
    .I1(__52__),
    .I0(__51__),
    .O(__76__)
  );
  LUT5 #(
    .INIT(32'hb8f0aaaa)
  ) __283__ (
    .I4(G14),
    .I3(__70__),
    .I2(__60__),
    .I1(__76__),
    .I0(G8),
    .O(__77__)
  );
  LUT5 #(
    .INIT(32'hee44cfc0)
  ) __286__ (
    .I4(__69__),
    .I3(__64__),
    .I2(G8),
    .I1(__63__),
    .I0(__43__),
    .O(__80__)
  );
  LUT5 #(
    .INIT(32'h0088000f)
  ) __287__ (
    .I4(__69__),
    .I3(__25__),
    .I2(G4),
    .I1(__57__),
    .I0(__80__),
    .O(__81__)
  );
  LUT5 #(
    .INIT(32'hca000000)
  ) __288__ (
    .I4(__69__),
    .I3(__54__),
    .I2(__43__),
    .I1(__64__),
    .I0(__63__),
    .O(__82__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __289__ (
    .I1(__69__),
    .I0(G1),
    .O(__83__)
  );
  LUT5 #(
    .INIT(32'hca000000)
  ) __290__ (
    .I4(__69__),
    .I3(__53__),
    .I2(__43__),
    .I1(__64__),
    .I0(__63__),
    .O(__84__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __291__ (
    .I1(__69__),
    .I0(G0),
    .O(__85__)
  );
  LUT6 #(
    .INIT(64'h020202ab02020202)
  ) __292__ (
    .I5(__21__),
    .I4(__85__),
    .I3(__84__),
    .I2(__83__),
    .I1(__82__),
    .I0(__22__),
    .O(__86__)
  );
  LUT5 #(
    .INIT(32'hc0553faa)
  ) __293__ (
    .I4(__23__),
    .I3(__69__),
    .I2(__80__),
    .I1(__55__),
    .I0(G2),
    .O(__87__)
  );
  LUT4 #(
    .INIT(16'h77f0)
  ) __294__ (
    .I3(__69__),
    .I2(G3),
    .I1(__80__),
    .I0(__56__),
    .O(__88__)
  );
  LUT5 #(
    .INIT(32'hc0553faa)
  ) __295__ (
    .I4(__25__),
    .I3(__69__),
    .I2(__57__),
    .I1(__80__),
    .I0(G4),
    .O(__89__)
  );
  LUT6 #(
    .INIT(64'h044f0000077f0000)
  ) __296__ (
    .I5(__23__),
    .I4(__89__),
    .I3(__24__),
    .I2(__88__),
    .I1(__87__),
    .I0(__86__),
    .O(__90__)
  );
  LUT6 #(
    .INIT(64'h000e000000000000)
  ) __297__ (
    .I5(__19__),
    .I4(__16__),
    .I3(__10__),
    .I2(__13__),
    .I1(__90__),
    .I0(__81__),
    .O(__91__)
  );
  LUT6 #(
    .INIT(64'h008f000000000000)
  ) __298__ (
    .I5(__7__),
    .I4(__6__),
    .I3(__8__),
    .I2(__71__),
    .I1(__9__),
    .I0(__91__),
    .O(__92__)
  );
  LUT6 #(
    .INIT(64'h000000004000ffff)
  ) __299__ (
    .I5(__17__),
    .I4(__71__),
    .I3(__5__),
    .I2(__11__),
    .I1(__92__),
    .I0(__4__),
    .O(__93__)
  );
  LUT6 #(
    .INIT(64'h000040ff00000000)
  ) __300__ (
    .I5(__1__),
    .I4(__2__),
    .I3(__70__),
    .I2(__20__),
    .I1(__93__),
    .I0(__12__),
    .O(__94__)
  );
  LUT3 #(
    .INIT(8'h80)
  ) __301__ (
    .I2(__5__),
    .I1(__11__),
    .I0(__92__),
    .O(__95__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __302__ (
    .I1(__55__),
    .I0(__60__),
    .O(__96__)
  );
  LUT2 #(
    .INIT(4'h6)
  ) __303__ (
    .I1(__56__),
    .I0(__61__),
    .O(__97__)
  );
  LUT6 #(
    .INIT(64'h1001000000001001)
  ) __304__ (
    .I5(__53__),
    .I4(__58__),
    .I3(__54__),
    .I2(__59__),
    .I1(__97__),
    .I0(__96__),
    .O(__98__)
  );
  LUT6 #(
    .INIT(64'h0001fffe00000000)
  ) __305__ (
    .I5(__98__),
    .I4(__57__),
    .I3(__59__),
    .I2(__58__),
    .I1(__61__),
    .I0(__60__),
    .O(__99__)
  );
  LUT5 #(
    .INIT(32'hefff0000)
  ) __306__ (
    .I4(__69__),
    .I3(G16),
    .I2(__99__),
    .I1(__62__),
    .I0(__45__),
    .O(__100__)
  );
  LUT6 #(
    .INIT(64'hbbbbbbbb0fff0000)
  ) __307__ (
    .I5(__100__),
    .I4(__71__),
    .I3(__4__),
    .I2(__95__),
    .I1(__94__),
    .I0(__18__),
    .O(__101__)
  );
  LUT3 #(
    .INIT(8'h04)
  ) __308__ (
    .I2(__99__),
    .I1(__53__),
    .I0(__101__),
    .O(__102__)
  );
  LUT4 #(
    .INIT(16'hcafa)
  ) __309__ (
    .I3(G14),
    .I2(__69__),
    .I1(__76__),
    .I0(G9),
    .O(__103__)
  );
  LUT5 #(
    .INIT(32'h007f0080)
  ) __310__ (
    .I4(__56__),
    .I3(__103__),
    .I2(__55__),
    .I1(__54__),
    .I0(__102__),
    .O(__104__)
  );
  LUT5 #(
    .INIT(32'hbfff0000)
  ) __311__ (
    .I4(__71__),
    .I3(__5__),
    .I2(__11__),
    .I1(__92__),
    .I0(__4__),
    .O(__105__)
  );
  LUT6 #(
    .INIT(64'h880f000000000000)
  ) __312__ (
    .I5(__38__),
    .I4(__37__),
    .I3(__100__),
    .I2(__105__),
    .I1(__18__),
    .I0(__94__),
    .O(__106__)
  );
  LUT6 #(
    .INIT(64'h7f000000ffff0000)
  ) __313__ (
    .I5(__106__),
    .I4(__69__),
    .I3(__70__),
    .I2(__32__),
    .I1(__40__),
    .I0(__41__),
    .O(__107__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __314__ (
    .I1(G14),
    .I0(__76__),
    .O(__108__)
  );
  LUT6 #(
    .INIT(64'hbfff400000000000)
  ) __315__ (
    .I5(__108__),
    .I4(__49__),
    .I3(__48__),
    .I2(__47__),
    .I1(__46__),
    .I0(__107__),
    .O(__109__)
  );
  LUT6 #(
    .INIT(64'h5555055555554444)
  ) __316__ (
    .I5(__69__),
    .I4(__25__),
    .I3(__57__),
    .I2(__80__),
    .I1(G4),
    .I0(__90__),
    .O(__110__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __317__ (
    .I2(G14),
    .I1(__13__),
    .I0(__110__),
    .O(__111__)
  );
  LUT6 #(
    .INIT(64'he1f0f0f000000000)
  ) __318__ (
    .I5(G14),
    .I4(__19__),
    .I3(__16__),
    .I2(__10__),
    .I1(__13__),
    .I0(__110__),
    .O(__112__)
  );
  LUT4 #(
    .INIT(16'h0e01)
  ) __319__ (
    .I3(__53__),
    .I2(__103__),
    .I1(__99__),
    .I0(__101__),
    .O(__113__)
  );
  LUT6 #(
    .INIT(64'h9aaa555500000000)
  ) __320__ (
    .I5(G14),
    .I4(__70__),
    .I3(__20__),
    .I2(__93__),
    .I1(__12__),
    .I0(__2__),
    .O(__114__)
  );
  LUT4 #(
    .INIT(16'h008f)
  ) __321__ (
    .I3(__8__),
    .I2(__71__),
    .I1(__9__),
    .I0(__91__),
    .O(__115__)
  );
  LUT4 #(
    .INIT(16'h7800)
  ) __322__ (
    .I3(G14),
    .I2(__6__),
    .I1(__7__),
    .I0(__115__),
    .O(__116__)
  );
  LUT3 #(
    .INIT(8'h0b)
  ) __323__ (
    .I2(__69__),
    .I1(G14),
    .I0(__76__),
    .O(__117__)
  );
  LUT5 #(
    .INIT(32'hb8f0aaaa)
  ) __324__ (
    .I4(G14),
    .I3(__70__),
    .I2(__59__),
    .I1(__76__),
    .I0(G7),
    .O(__118__)
  );
  LUT6 #(
    .INIT(64'ha0c0ffffffffffff)
  ) __325__ (
    .I5(G13),
    .I4(G14),
    .I3(G10),
    .I2(__65__),
    .I1(__71__),
    .I0(__70__),
    .O(__119__)
  );
  LUT5 #(
    .INIT(32'h50230000)
  ) __326__ (
    .I4(G14),
    .I3(__30__),
    .I2(__70__),
    .I1(__32__),
    .I0(__106__),
    .O(__120__)
  );
  LUT6 #(
    .INIT(64'h4fffb00000000000)
  ) __327__ (
    .I5(G14),
    .I4(__41__),
    .I3(__32__),
    .I2(__40__),
    .I1(__70__),
    .I0(__106__),
    .O(__121__)
  );
  LUT4 #(
    .INIT(16'hca00)
  ) __328__ (
    .I3(G14),
    .I2(G11),
    .I1(__67__),
    .I0(__68__),
    .O(__122__)
  );
  LUT6 #(
    .INIT(64'h00008000aaaaaaaa)
  ) __329__ (
    .I5(__71__),
    .I4(__4__),
    .I3(__5__),
    .I2(__11__),
    .I1(__92__),
    .I0(__33__),
    .O(__123__)
  );
  LUT6 #(
    .INIT(64'hcaaacccc00000000)
  ) __330__ (
    .I5(G14),
    .I4(__70__),
    .I3(__123__),
    .I2(__35__),
    .I1(__26__),
    .I0(__27__),
    .O(__124__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __331__ (
    .I2(G15),
    .I1(__15__),
    .I0(__14__),
    .O(__125__)
  );
  LUT6 #(
    .INIT(64'h4000000000000000)
  ) __332__ (
    .I5(__21__),
    .I4(__26__),
    .I3(__27__),
    .I2(__28__),
    .I1(__29__),
    .I0(__125__),
    .O(__126__)
  );
  LUT6 #(
    .INIT(64'h050a112200001122)
  ) __333__ (
    .I5(G14),
    .I4(__69__),
    .I3(__22__),
    .I2(__76__),
    .I1(G7),
    .I0(__126__),
    .O(__127__)
  );
  LUT3 #(
    .INIT(8'h70)
  ) __334__ (
    .I2(G14),
    .I1(__69__),
    .I0(__76__),
    .O(__128__)
  );
  LUT5 #(
    .INIT(32'hf0f0ccaa)
  ) __335__ (
    .I4(__128__),
    .I3(__42__),
    .I2(__52__),
    .I1(G5),
    .I0(G2),
    .O(__129__)
  );
  LUT5 #(
    .INIT(32'hb8f0aaaa)
  ) __336__ (
    .I4(G14),
    .I3(__70__),
    .I2(__61__),
    .I1(__76__),
    .I0(G9),
    .O(__130__)
  );
  LUT3 #(
    .INIT(8'h60)
  ) __337__ (
    .I2(G14),
    .I1(__93__),
    .I0(__12__),
    .O(__131__)
  );
  LUT5 #(
    .INIT(32'h32013300)
  ) __338__ (
    .I4(__53__),
    .I3(__54__),
    .I2(__99__),
    .I1(__103__),
    .I0(__101__),
    .O(__132__)
  );
  LUT3 #(
    .INIT(8'he0)
  ) __339__ (
    .I2(G14),
    .I1(__76__),
    .I0(__44__),
    .O(__133__)
  );
  LUT6 #(
    .INIT(64'h555ff5ffcccccccc)
  ) __340__ (
    .I5(__69__),
    .I4(__64__),
    .I3(__63__),
    .I2(__43__),
    .I1(G0),
    .I0(__53__),
    .O(__134__)
  );
  LUT3 #(
    .INIT(8'he0)
  ) __341__ (
    .I2(__89__),
    .I1(__21__),
    .I0(__134__),
    .O(__135__)
  );
  LUT6 #(
    .INIT(64'h882200aa0aa00aa0)
  ) __342__ (
    .I5(__69__),
    .I4(__80__),
    .I3(__24__),
    .I2(G3),
    .I1(__56__),
    .I0(__87__),
    .O(__136__)
  );
  LUT6 #(
    .INIT(64'h4141c3c34144c3cc)
  ) __343__ (
    .I5(__69__),
    .I4(__21__),
    .I3(G1),
    .I2(__82__),
    .I1(__22__),
    .I0(__134__),
    .O(__137__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __344__ (
    .I1(__99__),
    .I0(__62__),
    .O(__138__)
  );
  LUT6 #(
    .INIT(64'h7f7f0000007f007f)
  ) __345__ (
    .I5(__69__),
    .I4(__138__),
    .I3(G5),
    .I2(__137__),
    .I1(__136__),
    .I0(__135__),
    .O(__139__)
  );
  LUT5 #(
    .INIT(32'hf0f055cc)
  ) __346__ (
    .I4(__100__),
    .I3(__71__),
    .I2(__18__),
    .I1(__3__),
    .I0(__4__),
    .O(__140__)
  );
  LUT5 #(
    .INIT(32'h33550f0f)
  ) __347__ (
    .I4(__69__),
    .I3(__70__),
    .I2(__3__),
    .I1(__41__),
    .I0(__38__),
    .O(__141__)
  );
  LUT6 #(
    .INIT(64'h03000000aaaaaaaa)
  ) __348__ (
    .I5(__69__),
    .I4(G16),
    .I3(__99__),
    .I2(__62__),
    .I1(__45__),
    .I0(G6),
    .O(__142__)
  );
  LUT6 #(
    .INIT(64'h0f0f00bb00000000)
  ) __349__ (
    .I5(G14),
    .I4(__142__),
    .I3(__110__),
    .I2(__141__),
    .I1(__140__),
    .I0(__139__),
    .O(__143__)
  );
  LUT5 #(
    .INIT(32'h7f800000)
  ) __350__ (
    .I4(G14),
    .I3(__4__),
    .I2(__5__),
    .I1(__11__),
    .I0(__92__),
    .O(__144__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __351__ (
    .I2(G14),
    .I1(__17__),
    .I0(__105__),
    .O(__145__)
  );
  LUT4 #(
    .INIT(16'hca00)
  ) __352__ (
    .I3(G14),
    .I2(__76__),
    .I1(__44__),
    .I0(__45__),
    .O(__146__)
  );
  LUT3 #(
    .INIT(8'h60)
  ) __353__ (
    .I2(G14),
    .I1(__9__),
    .I0(__91__),
    .O(__147__)
  );
  LUT6 #(
    .INIT(64'hd000000000000000)
  ) __354__ (
    .I5(__32__),
    .I4(__40__),
    .I3(__41__),
    .I2(__68__),
    .I1(__106__),
    .I0(__70__),
    .O(__148__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __355__ (
    .I1(__9__),
    .I0(__91__),
    .O(__149__)
  );
  LUT3 #(
    .INIT(8'h08)
  ) __356__ (
    .I2(__12__),
    .I1(__20__),
    .I0(__93__),
    .O(__150__)
  );
  LUT5 #(
    .INIT(32'h40000000)
  ) __357__ (
    .I4(__5__),
    .I3(__11__),
    .I2(__92__),
    .I1(__66__),
    .I0(__4__),
    .O(__151__)
  );
  LUT6 #(
    .INIT(64'h0000000000005f13)
  ) __358__ (
    .I5(__69__),
    .I4(__151__),
    .I3(__73__),
    .I2(__150__),
    .I1(__149__),
    .I0(__67__),
    .O(__152__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __359__ (
    .I1(__152__),
    .I0(__148__),
    .O(__153__)
  );
  LUT4 #(
    .INIT(16'h8000)
  ) __360__ (
    .I3(G14),
    .I2(__80__),
    .I1(__62__),
    .I0(__140__),
    .O(__154__)
  );
  LUT3 #(
    .INIT(8'h60)
  ) __361__ (
    .I2(G14),
    .I1(__11__),
    .I0(__92__),
    .O(__155__)
  );
  LUT6 #(
    .INIT(64'h44ff0b0000000000)
  ) __362__ (
    .I5(G14),
    .I4(__39__),
    .I3(__32__),
    .I2(__40__),
    .I1(__70__),
    .I0(__106__),
    .O(__156__)
  );
  LUT4 #(
    .INIT(16'h5c00)
  ) __363__ (
    .I3(G14),
    .I2(G11),
    .I1(__66__),
    .I0(__73__),
    .O(__157__)
  );
  LUT6 #(
    .INIT(64'h00000000bf400000)
  ) __364__ (
    .I5(__76__),
    .I4(G14),
    .I3(__48__),
    .I2(__47__),
    .I1(__46__),
    .I0(__107__),
    .O(__158__)
  );
  LUT6 #(
    .INIT(64'hcaaacccc00000000)
  ) __365__ (
    .I5(G14),
    .I4(__70__),
    .I3(__123__),
    .I2(__35__),
    .I1(__28__),
    .I0(__29__),
    .O(__159__)
  );
  LUT4 #(
    .INIT(16'hcafa)
  ) __366__ (
    .I3(G14),
    .I2(__69__),
    .I1(__76__),
    .I0(G7),
    .O(__160__)
  );
  LUT4 #(
    .INIT(16'h0708)
  ) __367__ (
    .I3(__23__),
    .I2(__160__),
    .I1(__22__),
    .I0(__126__),
    .O(__161__)
  );
  LUT5 #(
    .INIT(32'h0000b400)
  ) __368__ (
    .I4(__76__),
    .I3(G14),
    .I2(__47__),
    .I1(__46__),
    .I0(__107__),
    .O(__162__)
  );
  LUT4 #(
    .INIT(16'h880f)
  ) __369__ (
    .I3(__100__),
    .I2(__105__),
    .I1(__18__),
    .I0(__94__),
    .O(__163__)
  );
  LUT4 #(
    .INIT(16'h2c00)
  ) __370__ (
    .I3(G14),
    .I2(__163__),
    .I1(__37__),
    .I0(__36__),
    .O(__164__)
  );
  LUT4 #(
    .INIT(16'hc300)
  ) __371__ (
    .I3(G14),
    .I2(__105__),
    .I1(__33__),
    .I0(__35__),
    .O(__165__)
  );
  LUT5 #(
    .INIT(32'h0000af03)
  ) __372__ (
    .I4(__103__),
    .I3(__62__),
    .I2(__99__),
    .I1(__101__),
    .I0(__140__),
    .O(__166__)
  );
  LUT4 #(
    .INIT(16'h1c00)
  ) __373__ (
    .I3(G14),
    .I2(__163__),
    .I1(__36__),
    .I0(__37__),
    .O(__167__)
  );
  LUT6 #(
    .INIT(64'h00007fff00008000)
  ) __374__ (
    .I5(__25__),
    .I4(__160__),
    .I3(__23__),
    .I2(__24__),
    .I1(__22__),
    .I0(__126__),
    .O(__168__)
  );
  LUT4 #(
    .INIT(16'h5c00)
  ) __375__ (
    .I3(G14),
    .I2(G11),
    .I1(__73__),
    .I0(__68__),
    .O(__169__)
  );
  LUT5 #(
    .INIT(32'h40000000)
  ) __376__ (
    .I4(__26__),
    .I3(__27__),
    .I2(__28__),
    .I1(__29__),
    .I0(__125__),
    .O(__170__)
  );
  LUT6 #(
    .INIT(64'h00007fff00008000)
  ) __377__ (
    .I5(__24__),
    .I4(__160__),
    .I3(__23__),
    .I2(__21__),
    .I1(__22__),
    .I0(__170__),
    .O(__171__)
  );
  LUT5 #(
    .INIT(32'hf0f0ccaa)
  ) __378__ (
    .I4(__128__),
    .I3(__42__),
    .I2(__51__),
    .I1(G4),
    .I0(G1),
    .O(__172__)
  );
  LUT6 #(
    .INIT(64'hcaaacccc00000000)
  ) __379__ (
    .I5(G14),
    .I4(__70__),
    .I3(__123__),
    .I2(__35__),
    .I1(G12),
    .I0(__26__),
    .O(__173__)
  );
  LUT5 #(
    .INIT(32'hef100000)
  ) __380__ (
    .I4(G14),
    .I3(__19__),
    .I2(__16__),
    .I1(__13__),
    .I0(__110__),
    .O(__174__)
  );
  LUT6 #(
    .INIT(64'h3233333301000000)
  ) __381__ (
    .I5(__55__),
    .I4(__53__),
    .I3(__54__),
    .I2(__99__),
    .I1(__103__),
    .I0(__101__),
    .O(__175__)
  );
  LUT5 #(
    .INIT(32'hb8f0aaaa)
  ) __382__ (
    .I4(G14),
    .I3(__70__),
    .I2(__58__),
    .I1(__76__),
    .I0(G6),
    .O(__176__)
  );
  LUT6 #(
    .INIT(64'h050a112200001122)
  ) __383__ (
    .I5(G14),
    .I4(__69__),
    .I3(__21__),
    .I2(__76__),
    .I1(G7),
    .I0(__170__),
    .O(__177__)
  );
  LUT4 #(
    .INIT(16'h0090)
  ) __384__ (
    .I3(__76__),
    .I2(G14),
    .I1(__46__),
    .I0(__107__),
    .O(__178__)
  );
  LUT4 #(
    .INIT(16'h7800)
  ) __385__ (
    .I3(G14),
    .I2(__38__),
    .I1(__37__),
    .I0(__163__),
    .O(__179__)
  );
  LUT6 #(
    .INIT(64'h00007fff00008000)
  ) __386__ (
    .I5(__57__),
    .I4(__103__),
    .I3(__56__),
    .I2(__55__),
    .I1(__54__),
    .I0(__102__),
    .O(__180__)
  );
  LUT4 #(
    .INIT(16'h7800)
  ) __387__ (
    .I3(G14),
    .I2(__5__),
    .I1(__11__),
    .I0(__92__),
    .O(__181__)
  );
  LUT5 #(
    .INIT(32'h6a550000)
  ) __388__ (
    .I4(G14),
    .I3(__71__),
    .I2(__9__),
    .I1(__91__),
    .I0(__8__),
    .O(__182__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __389__ (
    .I1(G14),
    .I0(__3__),
    .O(__183__)
  );
  LUT5 #(
    .INIT(32'hf0f0ccaa)
  ) __390__ (
    .I4(__128__),
    .I3(__42__),
    .I2(__50__),
    .I1(G3),
    .I0(G0),
    .O(__184__)
  );
  LUT6 #(
    .INIT(64'hcaaacccc00000000)
  ) __391__ (
    .I5(G14),
    .I4(__70__),
    .I3(__123__),
    .I2(__35__),
    .I1(__27__),
    .I0(__28__),
    .O(__185__)
  );
  LUT4 #(
    .INIT(16'hca00)
  ) __392__ (
    .I3(G14),
    .I2(G11),
    .I1(__66__),
    .I0(__67__),
    .O(__186__)
  );
  LUT5 #(
    .INIT(32'hb8f0aaaa)
  ) __393__ (
    .I4(G14),
    .I3(__70__),
    .I2(__63__),
    .I1(__76__),
    .I0(G10),
    .O(__187__)
  );
  LUT4 #(
    .INIT(16'h1c00)
  ) __394__ (
    .I3(G14),
    .I2(__123__),
    .I1(__34__),
    .I0(__35__),
    .O(__188__)
  );
  LUT5 #(
    .INIT(32'he0ffffff)
  ) __395__ (
    .I4(G13),
    .I3(G14),
    .I2(__65__),
    .I1(G10),
    .I0(__69__),
    .O(__189__)
  );
  LUT6 #(
    .INIT(64'h44ffb00000000000)
  ) __396__ (
    .I5(G14),
    .I4(__40__),
    .I3(__32__),
    .I2(__39__),
    .I1(__70__),
    .I0(__106__),
    .O(__190__)
  );
  LUT6 #(
    .INIT(64'hfffffffe40000000)
  ) __397__ (
    .I5(__15__),
    .I4(__26__),
    .I3(__27__),
    .I2(__28__),
    .I1(__29__),
    .I0(G15),
    .O(__191__)
  );
  LUT4 #(
    .INIT(16'h2c00)
  ) __398__ (
    .I3(G14),
    .I2(__123__),
    .I1(__35__),
    .I0(__34__),
    .O(__192__)
  );
  LUT4 #(
    .INIT(16'he100)
  ) __399__ (
    .I3(G14),
    .I2(__16__),
    .I1(__13__),
    .I0(__110__),
    .O(__193__)
  );
  LUT5 #(
    .INIT(32'hb8f0aaaa)
  ) __400__ (
    .I4(G14),
    .I3(__70__),
    .I2(__64__),
    .I1(__76__),
    .I0(G11),
    .O(__194__)
  );
  LUT6 #(
    .INIT(64'h4444b00000000000)
  ) __401__ (
    .I5(G14),
    .I4(__32__),
    .I3(__31__),
    .I2(__30__),
    .I1(__70__),
    .I0(__106__),
    .O(__195__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __402__ (
    .I1(G13),
    .I0(G14),
    .O(__196__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __403__ (
    .I1(__93__),
    .I0(__12__),
    .O(__197__)
  );
  LUT6 #(
    .INIT(64'hff70008f00000000)
  ) __404__ (
    .I5(G14),
    .I4(__1__),
    .I3(__2__),
    .I2(__70__),
    .I1(__20__),
    .I0(__197__),
    .O(__198__)
  );
  LUT6 #(
    .INIT(64'h444f0b0000000000)
  ) __405__ (
    .I5(G14),
    .I4(__31__),
    .I3(__30__),
    .I2(__32__),
    .I1(__70__),
    .I0(__106__),
    .O(__199__)
  );
  LUT3 #(
    .INIT(8'h60)
  ) __406__ (
    .I2(G14),
    .I1(__18__),
    .I0(__94__),
    .O(__200__)
  );
  LUT4 #(
    .INIT(16'hca00)
  ) __407__ (
    .I3(G14),
    .I2(__76__),
    .I1(__42__),
    .I0(__43__),
    .O(__201__)
  );
  LUT4 #(
    .INIT(16'hb400)
  ) __408__ (
    .I3(G14),
    .I2(__20__),
    .I1(__93__),
    .I0(__12__),
    .O(__202__)
  );
  LUT3 #(
    .INIT(8'he0)
  ) __409__ (
    .I2(G14),
    .I1(__140__),
    .I0(__42__),
    .O(__203__)
  );
  LUT6 #(
    .INIT(64'hff70008f00000000)
  ) __410__ (
    .I5(G14),
    .I4(__7__),
    .I3(__8__),
    .I2(__71__),
    .I1(__9__),
    .I0(__91__),
    .O(__204__)
  );
  LUT6 #(
    .INIT(64'ha0c0ffffffffffff)
  ) __411__ (
    .I5(G13),
    .I4(G14),
    .I3(G10),
    .I2(__65__),
    .I1(__70__),
    .I0(__69__),
    .O(__205__)
  );
  assign G729 = __74__;
  assign G727 = __117__;
  assign G702 = __153__;
  assign G726 = __72__;
  assign G701BF = __0__;
endmodule
