module max512 (
    x0,
    x1,
    x2,
    x3,
    x4,
    x5,
    x6,
    x7,
    x8,
    y0,
    y1,
    y2,
    y3,
    y4,
    y5
);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8;
  output y0, y1, y2, y3, y4, y5;
  wire n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 ;
  assign n10  = x5 & x7;
  assign n11  = (~x4 & x6) | (~x4 & n10) | (x6 & n10);
  assign n12  = x4 & n11;
  assign n13  = x2 & x3;
  assign n14  = (x0 & n12) | (x0 & n13) | (n12 & n13);
  assign n15  = x1 & ~n14;
  assign n16  = (x0 & x1) | (x0 & ~n15) | (x1 & ~n15);
  assign n17  = (x2 & ~x6) | (x2 & x7) | (~x6 & x7);
  assign n18  = (x3 & x7) | (x3 & ~n17) | (x7 & ~n17);
  assign n19  = (~x2 & x3) | (~x2 & n17) | (x3 & n17);
  assign n20  = n18 & ~n19;
  assign n21  = x1 & x5;
  assign n22  = (x4 & ~n20) | (x4 & n21) | (~n20 & n21);
  assign n23  = n20 & n22;
  assign n47  = x0 & n23;
  assign n24  = ~x0 & x2;
  assign n25  = x1 & n24;
  assign n26  = x5 & ~x6;
  assign n27  = x4 & n26;
  assign n28  = (x3 & ~n25) | (x3 & n27) | (~n25 & n27);
  assign n29  = n25 & n28;
  assign n37  = ~x0 & x1;
  assign n38  = x1 & ~x3;
  assign n39  = (x0 & x2) | (x0 & n38) | (x2 & n38);
  assign n40  = (~x2 & x3) | (~x2 & n39) | (x3 & n39);
  assign n41  = (x1 & n39) | (x1 & n40) | (n39 & n40);
  assign n35  = x2 & ~x4;
  assign n36  = x3 & n35;
  assign n42  = n36 | n41;
  assign n43  = (n37 & n41) | (n37 & n42) | (n41 & n42);
  assign n30  = (x0 & x1) | (x0 & x5) | (x1 & x5);
  assign n31  = (x1 & ~x3) | (x1 & n30) | (~x3 & n30);
  assign n32  = x1 & ~n31;
  assign n33  = n31 | n32;
  assign n34  = (~x1 & n32) | (~x1 & n33) | (n32 & n33);
  assign n44  = (x2 & n34) | (x2 & n43) | (n34 & n43);
  assign n45  = x4 & ~n44;
  assign n46  = (x4 & n43) | (x4 & ~n45) | (n43 & ~n45);
  assign n48  = n29 | n46;
  assign n49  = (n23 & ~n47) | (n23 & n48) | (~n47 & n48);
  assign n54  = x6 | x7;
  assign n55  = x5 | n54;
  assign n56  = x4 & ~n55;
  assign n57  = (x0 & x2) | (x0 & n56) | (x2 & n56);
  assign n58  = ~x0 & n57;
  assign n50  = x6 & n10;
  assign n51  = x0 & ~x4;
  assign n52  = (x2 & n50) | (x2 & n51) | (n50 & n51);
  assign n53  = ~x2 & n52;
  assign n59  = n53 & ~n58;
  assign n60  = ~x3 & x8;
  assign n61  = (n58 & n59) | (n58 & n60) | (n59 & n60);
  assign n126 = ~x1 & n61;
  assign n65  = (x2 & ~x3) | (x2 & x6) | (~x3 & x6);
  assign n66  = (x1 & ~x6) | (x1 & n65) | (~x6 & n65);
  assign n67  = (x2 & ~x3) | (x2 & n66) | (~x3 & n66);
  assign n68  = ~n65 & n67;
  assign n69  = (~n66 & n67) | (~n66 & n68) | (n67 & n68);
  assign n70  = x4 & n69;
  assign n71  = x0 | n70;
  assign n62  = x1 | x2;
  assign n63  = ~x4 & x6;
  assign n64  = x3 & n63;
  assign n72  = ~n62 & n64;
  assign n73  = x0 & ~n72;
  assign n74  = n71 & ~n73;
  assign n102 = ~x5 & n74;
  assign n75  = ~x3 & x4;
  assign n76  = ~x5 & x6;
  assign n77  = n25 & n76;
  assign n78  = n75 & n77;
  assign n79  = (x2 & x3) | (x2 & ~x4) | (x3 & ~x4);
  assign n80  = (x0 & ~x3) | (x0 & n79) | (~x3 & n79);
  assign n81  = (~x2 & x3) | (~x2 & n80) | (x3 & n80);
  assign n82  = n79 & ~n81;
  assign n83  = (x0 & ~n80) | (x0 & n82) | (~n80 & n82);
  assign n89  = (~x2 & x3) | (~x2 & x5) | (x3 & x5);
  assign n90  = x2 & ~x5;
  assign n91  = (x1 & x3) | (x1 & ~n90) | (x3 & ~n90);
  assign n92  = ~n89 & n91;
  assign n96  = (x0 & x4) | (x0 & n92) | (x4 & n92);
  assign n93  = x0 & ~x1;
  assign n94  = (x3 & n90) | (x3 & n93) | (n90 & n93);
  assign n95  = ~x3 & n94;
  assign n97  = x4 & n95;
  assign n98  = (~x0 & n96) | (~x0 & n97) | (n96 & n97);
  assign n99  = (~x1 & n83) | (~x1 & n98) | (n83 & n98);
  assign n84  = ~x0 & x4;
  assign n85  = (x0 & x2) | (x0 & x3) | (x2 & x3);
  assign n86  = (x0 & x2) | (x0 & ~x4) | (x2 & ~x4);
  assign n87  = x3 | n86;
  assign n88  = (n84 & ~n85) | (n84 & n87) | (~n85 & n87);
  assign n100 = (x1 & ~n88) | (x1 & n98) | (~n88 & n98);
  assign n101 = n99 | n100;
  assign n103 = n78 | n101;
  assign n104 = (n74 & ~n102) | (n74 & n103) | (~n102 & n103);
  assign n117 = ~x6 & x7;
  assign n118 = (x4 & x5) | (x4 & n117) | (x5 & n117);
  assign n119 = ~x4 & n118;
  assign n120 = x3 & n119;
  assign n121 = (x2 & n93) | (x2 & n120) | (n93 & n120);
  assign n122 = ~x2 & n121;
  assign n105 = (x3 & ~x5) | (x3 & x7) | (~x5 & x7);
  assign n106 = (x3 & ~x6) | (x3 & n105) | (~x6 & n105);
  assign n107 = x3 & ~n106;
  assign n108 = n106 | n107;
  assign n109 = (~x3 & n107) | (~x3 & n108) | (n107 & n108);
  assign n114 = (x2 & x4) | (x2 & ~n109) | (x4 & ~n109);
  assign n110 = x2 | x3;
  assign n111 = x5 & ~n110;
  assign n112 = (x6 & x7) | (x6 & n111) | (x7 & n111);
  assign n113 = ~x7 & n112;
  assign n115 = x4 & n113;
  assign n116 = (n109 & n114) | (n109 & n115) | (n114 & n115);
  assign n123 = (~x0 & n116) | (~x0 & n122) | (n116 & n122);
  assign n124 = x1 & ~n123;
  assign n125 = (x1 & n122) | (x1 & ~n124) | (n122 & ~n124);
  assign n127 = n104 | n125;
  assign n128 = (n61 & ~n126) | (n61 & n127) | (~n126 & n127);
  assign n145 = (~x2 & x3) | (~x2 & x4) | (x3 & x4);
  assign n146 = (~x2 & x5) | (~x2 & n145) | (x5 & n145);
  assign n147 = (x4 & x5) | (x4 & ~n146) | (x5 & ~n146);
  assign n148 = x3 & n147;
  assign n149 = (x2 & n146) | (x2 & ~n148) | (n146 & ~n148);
  assign n150 = x0 & ~n149;
  assign n143 = x3 & x5;
  assign n144 = (~x3 & n35) | (~x3 & n143) | (n35 & n143);
  assign n151 = x0 | n144;
  assign n152 = (~x0 & n150) | (~x0 & n151) | (n150 & n151);
  assign n153 = x1 & ~n152;
  assign n139 = (x3 & x4) | (x3 & x5) | (x4 & x5);
  assign n140 = (x0 & x3) | (x0 & ~x4) | (x3 & ~x4);
  assign n141 = n139 | n140;
  assign n142 = (~x5 & n139) | (~x5 & n141) | (n139 & n141);
  assign n154 = x2 & ~n142;
  assign n155 = x1 | n154;
  assign n156 = ~n153 & n155;
  assign n134 = x4 & x5;
  assign n135 = x3 & ~n134;
  assign n136 = (x1 & x3) | (x1 & ~n134) | (x3 & ~n134);
  assign n137 = ~n135 & n136;
  assign n138 = (x3 & ~n135) | (x3 & n137) | (~n135 & n137);
  assign n157 = (~x0 & x2) | (~x0 & n138) | (x2 & n138);
  assign n158 = (~n24 & n156) | (~n24 & n157) | (n156 & n157);
  assign n159 = ~x1 & x2;
  assign n129 = (x0 & x4) | (x0 & x5) | (x4 & x5);
  assign n130 = (x3 & ~x5) | (x3 & n129) | (~x5 & n129);
  assign n131 = (x0 & x4) | (x0 & n130) | (x4 & n130);
  assign n132 = ~n129 & n131;
  assign n133 = (~n130 & n131) | (~n130 & n132) | (n131 & n132);
  assign n160 = (~x1 & x2) | (~x1 & n133) | (x2 & n133);
  assign n161 = (n158 & ~n159) | (n158 & n160) | (~n159 & n160);
  assign n188 = x7 & x8;
  assign n189 = ~x6 & n188;
  assign n190 = (x4 & x5) | (x4 & n189) | (x5 & n189);
  assign n191 = ~x4 & n190;
  assign n206 = x6 | x8;
  assign n207 = (~x5 & x7) | (~x5 & n206) | (x7 & n206);
  assign n208 = x5 | n207;
  assign n209 = x4 & ~n208;
  assign n210 = (x2 & ~n37) | (x2 & n209) | (~n37 & n209);
  assign n211 = n37 & n210;
  assign n198 = ~x6 & x8;
  assign n199 = ~x7 & n198;
  assign n200 = ~x5 & n199;
  assign n201 = (x1 & x2) | (x1 & n200) | (x2 & n200);
  assign n202 = ~x1 & n201;
  assign n195 = ~x2 & x5;
  assign n196 = x1 & n195;
  assign n197 = x7 & ~x8;
  assign n203 = (n196 & n197) | (n196 & n202) | (n197 & n202);
  assign n204 = x6 & ~n203;
  assign n205 = (x6 & n202) | (x6 & ~n204) | (n202 & ~n204);
  assign n212 = (~x4 & n205) | (~x4 & n211) | (n205 & n211);
  assign n213 = x0 & ~n212;
  assign n214 = (x0 & n211) | (x0 & ~n213) | (n211 & ~n213);
  assign n215 = ~x3 & n214;
  assign n192 = x0 | x1;
  assign n193 = ~x2 & x3;
  assign n194 = ~n192 & n193;
  assign n216 = n194 | n215;
  assign n217 = (n191 & n215) | (n191 & n216) | (n215 & n216);
  assign n171 = (x3 & ~x4) | (x3 & x5) | (~x4 & x5);
  assign n172 = (x3 & ~x6) | (x3 & n171) | (~x6 & n171);
  assign n173 = x3 & ~n172;
  assign n174 = n172 | n173;
  assign n175 = (~x3 & n173) | (~x3 & n174) | (n173 & n174);
  assign n176 = x1 & ~n175;
  assign n170 = x4 & n76;
  assign n177 = ~x3 & n170;
  assign n178 = x1 | n177;
  assign n179 = ~n176 & n178;
  assign n180 = x2 | n179;
  assign n167 = (~x3 & x4) | (~x3 & x6) | (x4 & x6);
  assign n168 = (~x3 & x4) | (~x3 & x5) | (x4 & x5);
  assign n169 = n167 & ~n168;
  assign n181 = ~x1 & n169;
  assign n182 = x2 & ~n181;
  assign n183 = n180 & ~n182;
  assign n184 = x0 & ~n183;
  assign n162 = (x1 & x2) | (x1 & ~x3) | (x2 & ~x3);
  assign n163 = (x2 & x6) | (x2 & n38) | (x6 & n38);
  assign n164 = n162 & ~n163;
  assign n165 = x4 | n72;
  assign n166 = (n72 & n164) | (n72 & n165) | (n164 & n165);
  assign n185 = x5 & n166;
  assign n186 = x0 | n185;
  assign n187 = ~n184 & n186;
  assign n225 = (x3 & ~x4) | (x3 & x6) | (~x4 & x6);
  assign n226 = (x1 & ~x6) | (x1 & n225) | (~x6 & n225);
  assign n227 = (x1 & x3) | (x1 & ~n225) | (x3 & ~n225);
  assign n228 = n226 & ~n227;
  assign n229 = x0 & ~n228;
  assign n223 = ~x3 & x6;
  assign n224 = x4 & n223;
  assign n230 = x1 & n224;
  assign n231 = x0 | n230;
  assign n232 = ~n229 & n231;
  assign n236 = (x2 & x7) | (x2 & n232) | (x7 & n232);
  assign n233 = x3 & x6;
  assign n234 = (x4 & ~n25) | (x4 & n233) | (~n25 & n233);
  assign n235 = n25 & n234;
  assign n237 = ~x7 & n235;
  assign n238 = (n232 & ~n236) | (n232 & n237) | (~n236 & n237);
  assign n239 = x5 & n238;
  assign n218 = (~x3 & x4) | (~x3 & x7) | (x4 & x7);
  assign n219 = ~n167 & n218;
  assign n220 = ~x5 & n219;
  assign n221 = (x1 & x2) | (x1 & n220) | (x2 & n220);
  assign n222 = ~x1 & n221;
  assign n240 = n222 | n239;
  assign n241 = (x0 & n239) | (x0 & n240) | (n239 & n240);
  assign n242 = n187 | n241;
  assign n243 = (~n161 & n217) | (~n161 & n242) | (n217 & n242);
  assign n244 = n161 | n243;
  assign n271 = x3 & ~x5;
  assign n272 = ~x7 & n271;
  assign n273 = x0 & x2;
  assign n274 = (x1 & n272) | (x1 & n273) | (n272 & n273);
  assign n275 = ~x1 & n274;
  assign n276 = (x2 & ~x3) | (x2 & x7) | (~x3 & x7);
  assign n277 = (x5 & ~x7) | (x5 & n276) | (~x7 & n276);
  assign n278 = (x2 & x5) | (x2 & ~n276) | (x5 & ~n276);
  assign n279 = n277 & ~n278;
  assign n283 = (x0 & ~x1) | (x0 & n279) | (~x1 & n279);
  assign n280 = x3 & x7;
  assign n281 = x5 & n280;
  assign n282 = n159 & n281;
  assign n284 = ~x0 & n282;
  assign n285 = (n279 & ~n283) | (n279 & n284) | (~n283 & n284);
  assign n259 = x5 & ~x7;
  assign n286 = x3 & ~x7;
  assign n287 = ~x3 & x5;
  assign n288 = (~n259 & n286) | (~n259 & n287) | (n286 & n287);
  assign n289 = x4 & n288;
  assign n290 = x0 & ~x2;
  assign n291 = (x1 & n289) | (x1 & n290) | (n289 & n290);
  assign n292 = ~x1 & n291;
  assign n293 = (~n275 & n285) | (~n275 & n292) | (n285 & n292);
  assign n294 = x4 & ~n292;
  assign n295 = (n275 & n293) | (n275 & ~n294) | (n293 & ~n294);
  assign n296 = x6 & n295;
  assign n260 = ~x3 & n259;
  assign n261 = ~x4 & n260;
  assign n262 = x0 & n261;
  assign n263 = ~n62 & n262;
  assign n264 = (x2 & x5) | (x2 & ~x7) | (x5 & ~x7);
  assign n265 = (x4 & x5) | (x4 & ~n264) | (x5 & ~n264);
  assign n266 = (~x2 & x4) | (~x2 & n264) | (x4 & n264);
  assign n267 = n265 & ~n266;
  assign n268 = x3 & n267;
  assign n269 = (x0 & x1) | (x0 & n268) | (x1 & n268);
  assign n270 = ~x0 & n269;
  assign n297 = n263 | n270;
  assign n298 = ~x6 & n297;
  assign n299 = n296 | n298;
  assign n301 = ~x2 & x7;
  assign n302 = (x0 & ~x5) | (x0 & n301) | (~x5 & n301);
  assign n303 = (x2 & x5) | (x2 & n301) | (x5 & n301);
  assign n304 = (x0 & x7) | (x0 & ~n303) | (x7 & ~n303);
  assign n305 = ~n302 & n304;
  assign n306 = x4 | n305;
  assign n300 = x0 | x2;
  assign n307 = n259 & ~n300;
  assign n308 = x4 & ~n307;
  assign n309 = n306 & ~n308;
  assign n313 = (x3 & ~x6) | (x3 & n309) | (~x6 & n309);
  assign n310 = x4 & n259;
  assign n311 = (x0 & n13) | (x0 & n310) | (n13 & n310);
  assign n312 = ~x0 & n311;
  assign n314 = x6 & n312;
  assign n315 = (n309 & ~n313) | (n309 & n314) | (~n313 & n314);
  assign n365 = x2 | x5;
  assign n366 = (~x1 & x4) | (~x1 & n365) | (x4 & n365);
  assign n367 = x1 | n366;
  assign n359 = ~x1 & x5;
  assign n360 = ~x0 & x5;
  assign n361 = (n37 & n359) | (n37 & ~n360) | (n359 & ~n360);
  assign n362 = (x2 & x4) | (x2 & ~n361) | (x4 & ~n361);
  assign n363 = x2 & ~n362;
  assign n364 = (x4 & ~n362) | (x4 & n363) | (~n362 & n363);
  assign n368 = x0 & x1;
  assign n369 = ~x2 & x4;
  assign n370 = (n84 & n368) | (n84 & ~n369) | (n368 & ~n369);
  assign n371 = (~x1 & n368) | (~x1 & n370) | (n368 & n370);
  assign n372 = n364 | n371;
  assign n373 = n367 & ~n372;
  assign n383 = (x2 & n37) | (x2 & n287) | (n37 & n287);
  assign n384 = ~x2 & n383;
  assign n385 = x0 & ~x5;
  assign n386 = (n24 & ~n90) | (n24 & n385) | (~n90 & n385);
  assign n387 = (x1 & ~x3) | (x1 & n386) | (~x3 & n386);
  assign n388 = ~x1 & n387;
  assign n389 = (x3 & n387) | (x3 & n388) | (n387 & n388);
  assign n390 = (x3 & x5) | (x3 & x6) | (x5 & x6);
  assign n391 = ~x5 & n390;
  assign n392 = (~x3 & n390) | (~x3 & n391) | (n390 & n391);
  assign n393 = x2 & n392;
  assign n394 = (x0 & x1) | (x0 & n393) | (x1 & n393);
  assign n395 = ~x0 & n394;
  assign n396 = (~n384 & n389) | (~n384 & n395) | (n389 & n395);
  assign n397 = x6 & ~n395;
  assign n398 = (n384 & n396) | (n384 & ~n397) | (n396 & ~n397);
  assign n399 = x4 & ~n398;
  assign n374 = (~x0 & x1) | (~x0 & x6) | (x1 & x6);
  assign n375 = (x0 & ~x3) | (x0 & n374) | (~x3 & n374);
  assign n376 = (x1 & x6) | (x1 & n375) | (x6 & n375);
  assign n377 = ~n374 & n376;
  assign n378 = (~n375 & n376) | (~n375 & n377) | (n376 & n377);
  assign n379 = x2 | n378;
  assign n380 = n93 & n223;
  assign n381 = x2 & ~n380;
  assign n382 = n379 & ~n381;
  assign n400 = x5 & n382;
  assign n401 = x4 | n400;
  assign n402 = ~n399 & n401;
  assign n403 = (x3 & ~n373) | (x3 & n402) | (~n373 & n402);
  assign n352 = (~x1 & x5) | (~x1 & n37) | (x5 & n37);
  assign n353 = (x2 & n37) | (x2 & n352) | (n37 & n352);
  assign n354 = (x0 & ~x2) | (x0 & n353) | (~x2 & n353);
  assign n355 = n353 | n354;
  assign n356 = x4 & ~n355;
  assign n347 = x1 & ~x2;
  assign n348 = (x0 & x5) | (x0 & n347) | (x5 & n347);
  assign n349 = x5 | n348;
  assign n350 = x5 & n348;
  assign n351 = n349 & ~n350;
  assign n357 = x4 | n351;
  assign n358 = (~x4 & n356) | (~x4 & n357) | (n356 & n357);
  assign n404 = (~x3 & n358) | (~x3 & n402) | (n358 & n402);
  assign n405 = n403 | n404;
  assign n406 = (x1 & n315) | (x1 & n405) | (n315 & n405);
  assign n331 = (x3 & x5) | (x3 & x7) | (x5 & x7);
  assign n332 = (~x6 & x7) | (~x6 & n331) | (x7 & n331);
  assign n333 = x7 & ~n332;
  assign n334 = n332 | n333;
  assign n335 = (~x7 & n333) | (~x7 & n334) | (n333 & n334);
  assign n340 = (x2 & x4) | (x2 & n335) | (x4 & n335);
  assign n336 = ~x5 & x7;
  assign n337 = x6 & n336;
  assign n338 = ~x3 & n337;
  assign n339 = x2 & n338;
  assign n341 = ~x4 & n339;
  assign n342 = (n335 & ~n340) | (n335 & n341) | (~n340 & n341);
  assign n343 = ~x0 & n342;
  assign n316 = (x2 & x4) | (x2 & ~x6) | (x4 & ~x6);
  assign n317 = (x6 & x7) | (x6 & n316) | (x7 & n316);
  assign n318 = (x2 & x4) | (x2 & n317) | (x4 & n317);
  assign n319 = ~n316 & n318;
  assign n320 = (~n317 & n318) | (~n317 & n319) | (n318 & n319);
  assign n324 = (~x3 & x5) | (~x3 & n320) | (x5 & n320);
  assign n321 = ~x4 & x5;
  assign n322 = (x2 & ~n54) | (x2 & n321) | (~n54 & n321);
  assign n323 = ~x2 & n322;
  assign n325 = x3 & n323;
  assign n326 = (n320 & ~n324) | (n320 & n325) | (~n324 & n325);
  assign n327 = x5 & n117;
  assign n328 = ~x3 & n327;
  assign n329 = (x2 & ~x4) | (x2 & n328) | (~x4 & n328);
  assign n330 = ~x2 & n329;
  assign n344 = n326 | n330;
  assign n345 = x0 & n344;
  assign n346 = n343 | n345;
  assign n407 = (~x1 & n346) | (~x1 & n405) | (n346 & n405);
  assign n408 = n406 | n407;
  assign n409 = (x8 & n299) | (x8 & n408) | (n299 & n408);
  assign n250 = n25 & ~n54;
  assign n251 = (x4 & x5) | (x4 & n250) | (x5 & n250);
  assign n252 = ~x5 & n251;
  assign n245 = x1 & x2;
  assign n246 = x1 & ~n245;
  assign n247 = n50 & n246;
  assign n248 = (n55 & n245) | (n55 & ~n246) | (n245 & ~n246);
  assign n249 = (x2 & n247) | (x2 & ~n248) | (n247 & ~n248);
  assign n253 = (~x4 & n249) | (~x4 & n252) | (n249 & n252);
  assign n254 = x0 & ~n253;
  assign n255 = (x0 & n252) | (x0 & ~n254) | (n252 & ~n254);
  assign n256 = ~x3 & n255;
  assign n257 = n194 | n256;
  assign n258 = (n119 & n256) | (n119 & n257) | (n256 & n257);
  assign n410 = (~x8 & n258) | (~x8 & n408) | (n258 & n408);
  assign n411 = n409 | n410;
  assign n413 = ~x1 & x3;
  assign n414 = (n159 & n193) | (n159 & ~n413) | (n193 & ~n413);
  assign n415 = x0 & ~n414;
  assign n412 = ~x8 & n193;
  assign n416 = x1 & n412;
  assign n417 = x0 | n416;
  assign n418 = ~n415 & n417;
  assign n423 = (x6 & ~x7) | (x6 & n418) | (~x7 & n418);
  assign n419 = (x2 & x6) | (x2 & ~x8) | (x6 & ~x8);
  assign n420 = (x2 & x3) | (x2 & ~x8) | (x3 & ~x8);
  assign n421 = n419 & ~n420;
  assign n422 = n37 & n421;
  assign n424 = x7 & n422;
  assign n425 = (n418 & ~n423) | (n418 & n424) | (~n423 & n424);
  assign n426 = (x1 & x7) | (x1 & ~x8) | (x7 & ~x8);
  assign n427 = (~x3 & x7) | (~x3 & x8) | (x7 & x8);
  assign n428 = n426 | n427;
  assign n429 = x0 & ~x6;
  assign n430 = (x2 & ~n428) | (x2 & n429) | (~n428 & n429);
  assign n431 = ~x2 & n430;
  assign n432 = n425 | n431;
  assign n433 = (~x4 & x5) | (~x4 & n432) | (x5 & n432);
  assign n434 = (n321 & n432) | (n321 & ~n433) | (n432 & ~n433);
  assign n461 = n63 & n197;
  assign n465 = (~x0 & x7) | (~x0 & x8) | (x7 & x8);
  assign n466 = (x0 & ~x6) | (x0 & n465) | (~x6 & n465);
  assign n467 = (x7 & x8) | (x7 & n466) | (x8 & n466);
  assign n468 = ~n465 & n467;
  assign n469 = (~n466 & n467) | (~n466 & n468) | (n467 & n468);
  assign n470 = x1 | n469;
  assign n462 = (x6 & x7) | (x6 & x8) | (x7 & x8);
  assign n463 = x6 & ~n462;
  assign n464 = (x8 & ~n462) | (x8 & n463) | (~n462 & n463);
  assign n471 = ~x0 & n464;
  assign n472 = x1 & ~n471;
  assign n473 = n470 & ~n472;
  assign n476 = (x3 & x4) | (x3 & ~n473) | (x4 & ~n473);
  assign n460 = ~x3 & n37;
  assign n474 = ~x6 & n197;
  assign n475 = n460 & n474;
  assign n477 = x4 & n475;
  assign n478 = (n473 & n476) | (n473 & n477) | (n476 & n477);
  assign n479 = n460 | n478;
  assign n480 = (n461 & n478) | (n461 & n479) | (n478 & n479);
  assign n523 = (x2 & ~x5) | (x2 & n480) | (~x5 & n480);
  assign n507 = (x3 & ~x4) | (x3 & x8) | (~x4 & x8);
  assign n508 = (x3 & ~x7) | (x3 & n507) | (~x7 & n507);
  assign n509 = x3 & ~n508;
  assign n510 = n508 | n509;
  assign n511 = (~x3 & n509) | (~x3 & n510) | (n509 & n510);
  assign n512 = x1 & ~n511;
  assign n505 = x4 | x8;
  assign n506 = x7 | n505;
  assign n513 = x3 | n506;
  assign n514 = ~x1 & n513;
  assign n515 = n512 | n514;
  assign n516 = ~x6 & n515;
  assign n501 = (x3 & ~x7) | (x3 & x8) | (~x7 & x8);
  assign n502 = (x4 & ~x8) | (x4 & n501) | (~x8 & n501);
  assign n503 = (x3 & x4) | (x3 & ~n501) | (x4 & ~n501);
  assign n504 = n502 & ~n503;
  assign n517 = ~x1 & n504;
  assign n518 = x6 & ~n517;
  assign n519 = n516 | n518;
  assign n520 = x0 & ~n519;
  assign n455 = x7 | x8;
  assign n456 = (~x7 & n197) | (~x7 & n455) | (n197 & n455);
  assign n481 = (x1 & x6) | (x1 & n456) | (x6 & n456);
  assign n482 = (x3 & ~x6) | (x3 & n481) | (~x6 & n481);
  assign n483 = (x1 & x3) | (x1 & ~n481) | (x3 & ~n481);
  assign n484 = n482 & ~n483;
  assign n486 = (x3 & x6) | (x3 & ~x7) | (x6 & ~x7);
  assign n487 = (x3 & ~x8) | (x3 & n486) | (~x8 & n486);
  assign n488 = x3 & ~n487;
  assign n489 = n487 | n488;
  assign n490 = (~x3 & n488) | (~x3 & n489) | (n488 & n489);
  assign n491 = x1 & ~n490;
  assign n485 = x7 | n206;
  assign n492 = x3 | n485;
  assign n493 = ~x1 & n492;
  assign n494 = n491 | n493;
  assign n495 = x6 & n197;
  assign n496 = (x1 & n75) | (x1 & n495) | (n75 & n495);
  assign n497 = ~x1 & n496;
  assign n498 = (n484 & n494) | (n484 & ~n497) | (n494 & ~n497);
  assign n499 = x4 & ~n497;
  assign n500 = (~n484 & n498) | (~n484 & n499) | (n498 & n499);
  assign n521 = ~x0 & n500;
  assign n522 = (x0 & ~n520) | (x0 & n521) | (~n520 & n521);
  assign n524 = (x2 & x5) | (x2 & ~n522) | (x5 & ~n522);
  assign n525 = n523 & n524;
  assign n562 = (x2 & x3) | (x2 & ~x6) | (x3 & ~x6);
  assign n563 = (~x3 & x4) | (~x3 & n562) | (x4 & n562);
  assign n564 = (x2 & x4) | (x2 & ~n562) | (x4 & ~n562);
  assign n565 = n563 & ~n564;
  assign n566 = x1 & ~n565;
  assign n567 = x2 & n224;
  assign n568 = x1 | n567;
  assign n569 = ~n566 & n568;
  assign n570 = ~x5 & n569;
  assign n559 = x4 & x6;
  assign n560 = (x2 & x5) | (x2 & n559) | (x5 & n559);
  assign n561 = ~x2 & n560;
  assign n571 = n561 | n570;
  assign n572 = (~x1 & n570) | (~x1 & n571) | (n570 & n571);
  assign n573 = (x0 & x8) | (x0 & n572) | (x8 & n572);
  assign n574 = (x7 & ~x8) | (x7 & n573) | (~x8 & n573);
  assign n575 = (x0 & x7) | (x0 & ~n573) | (x7 & ~n573);
  assign n576 = n574 & ~n575;
  assign n537 = ~x7 & x8;
  assign n538 = x5 & n537;
  assign n539 = x4 & n538;
  assign n540 = x4 & x8;
  assign n541 = (x4 & x8) | (x4 & n288) | (x8 & n288);
  assign n542 = (n539 & ~n540) | (n539 & n541) | (~n540 & n541);
  assign n543 = x6 & ~n542;
  assign n534 = (~x3 & x5) | (~x3 & n501) | (x5 & n501);
  assign n535 = (~x5 & x7) | (~x5 & n501) | (x7 & n501);
  assign n536 = n534 & n535;
  assign n544 = x4 & n536;
  assign n545 = x6 | n544;
  assign n546 = ~n543 & n545;
  assign n547 = x0 & ~n546;
  assign n526 = (x6 & ~x7) | (x6 & x8) | (~x7 & x8);
  assign n527 = x6 & ~n526;
  assign n528 = (x3 & x8) | (x3 & n527) | (x8 & n527);
  assign n529 = (~n526 & n527) | (~n526 & n528) | (n527 & n528);
  assign n530 = x4 & ~n529;
  assign n531 = x3 & ~n485;
  assign n532 = x4 | n531;
  assign n533 = ~n530 & n532;
  assign n548 = x5 & n533;
  assign n549 = x0 | n548;
  assign n550 = ~n547 & n549;
  assign n556 = (x1 & x2) | (x1 & n550) | (x2 & n550);
  assign n551 = x1 & n75;
  assign n552 = x0 & n551;
  assign n553 = x6 & n188;
  assign n554 = (x5 & ~n552) | (x5 & n553) | (~n552 & n553);
  assign n555 = n552 & n554;
  assign n557 = ~x2 & n555;
  assign n558 = (n550 & ~n556) | (n550 & n557) | (~n556 & n557);
  assign n621 = (~x3 & x7) | (~x3 & n559) | (x7 & n559);
  assign n622 = (x3 & ~x6) | (x3 & n559) | (~x6 & n559);
  assign n623 = (x4 & x7) | (x4 & ~n622) | (x7 & ~n622);
  assign n624 = ~n621 & n623;
  assign n625 = ~x4 & n76;
  assign n626 = x3 & n625;
  assign n627 = x5 | n626;
  assign n628 = (n624 & n626) | (n624 & n627) | (n626 & n627);
  assign n629 = x0 | n628;
  assign n617 = (x4 & x5) | (x4 & x6) | (x5 & x6);
  assign n618 = (~x4 & x5) | (~x4 & x7) | (x5 & x7);
  assign n619 = ~n617 & n618;
  assign n620 = (x6 & ~n617) | (x6 & n619) | (~n617 & n619);
  assign n630 = ~x3 & n620;
  assign n631 = x0 & ~n630;
  assign n632 = n629 & ~n631;
  assign n633 = x2 & n632;
  assign n610 = (x4 & ~x6) | (x4 & x7) | (~x6 & x7);
  assign n611 = (x0 & x6) | (x0 & n610) | (x6 & n610);
  assign n612 = (x4 & x6) | (x4 & ~n611) | (x6 & ~n611);
  assign n613 = n610 | n612;
  assign n614 = (x0 & ~n611) | (x0 & n613) | (~n611 & n613);
  assign n615 = x5 & ~n614;
  assign n616 = x3 & n615;
  assign n634 = x2 | n616;
  assign n635 = (~x2 & n633) | (~x2 & n634) | (n633 & n634);
  assign n641 = (x1 & ~n110) | (x1 & n625) | (~n110 & n625);
  assign n642 = ~x1 & n641;
  assign n636 = (x3 & x4) | (x3 & x6) | (x4 & x6);
  assign n637 = (~x5 & x6) | (~x5 & n636) | (x6 & n636);
  assign n638 = x6 & ~n637;
  assign n639 = n637 | n638;
  assign n640 = (~x6 & n638) | (~x6 & n639) | (n638 & n639);
  assign n643 = (x1 & n640) | (x1 & n642) | (n640 & n642);
  assign n644 = x2 & ~n643;
  assign n645 = (x2 & n642) | (x2 & ~n644) | (n642 & ~n644);
  assign n646 = (x4 & ~x5) | (x4 & n636) | (~x5 & n636);
  assign n647 = x4 & ~n646;
  assign n648 = n646 | n647;
  assign n649 = (~x4 & n647) | (~x4 & n648) | (n647 & n648);
  assign n650 = ~x1 & x7;
  assign n651 = (x2 & n649) | (x2 & ~n650) | (n649 & ~n650);
  assign n652 = n649 & ~n651;
  assign n653 = x7 & ~n652;
  assign n654 = (n645 & n652) | (n645 & ~n653) | (n652 & ~n653);
  assign n655 = (x1 & n635) | (x1 & n654) | (n635 & n654);
  assign n596 = ~x3 & x7;
  assign n597 = (n287 & n336) | (n287 & ~n596) | (n336 & ~n596);
  assign n598 = x2 & x4;
  assign n599 = x2 & ~n598;
  assign n600 = n597 & n599;
  assign n601 = (n336 & ~n598) | (n336 & n599) | (~n598 & n599);
  assign n602 = (x4 & n600) | (x4 & n601) | (n600 & n601);
  assign n603 = x0 & n602;
  assign n592 = x2 | x4;
  assign n593 = x2 & ~x3;
  assign n594 = x5 & ~n593;
  assign n595 = (~n134 & n592) | (~n134 & n594) | (n592 & n594);
  assign n604 = ~x0 & n595;
  assign n605 = (x0 & ~n603) | (x0 & n604) | (~n603 & n604);
  assign n606 = x6 | n605;
  assign n577 = (x4 & ~x5) | (x4 & x7) | (~x5 & x7);
  assign n578 = x4 & ~n577;
  assign n579 = (x3 & ~x5) | (x3 & n578) | (~x5 & n578);
  assign n580 = (~n577 & n578) | (~n577 & n579) | (n578 & n579);
  assign n584 = (x0 & ~x2) | (x0 & n580) | (~x2 & n580);
  assign n581 = (~x3 & x4) | (~x3 & n105) | (x4 & n105);
  assign n582 = (~x4 & x5) | (~x4 & n105) | (x5 & n105);
  assign n583 = n581 & n582;
  assign n585 = (x0 & x2) | (x0 & ~n583) | (x2 & ~n583);
  assign n586 = n584 & ~n585;
  assign n587 = x4 & x7;
  assign n588 = x5 & n587;
  assign n589 = x0 & n588;
  assign n590 = (x2 & x3) | (x2 & n589) | (x3 & n589);
  assign n591 = ~x3 & n590;
  assign n607 = n586 | n591;
  assign n608 = x6 & n607;
  assign n609 = n606 & ~n608;
  assign n656 = (x1 & n609) | (x1 & ~n654) | (n609 & ~n654);
  assign n657 = ~n655 & n656;
  assign n658 = ~n558 & n657;
  assign n659 = (n525 & ~n576) | (n525 & n658) | (~n576 & n658);
  assign n660 = ~n525 & n659;
  assign n446 = (x1 & x3) | (x1 & x6) | (x3 & x6);
  assign n447 = (x5 & ~x6) | (x5 & n446) | (~x6 & n446);
  assign n448 = (x1 & x3) | (x1 & n447) | (x3 & n447);
  assign n449 = ~n446 & n448;
  assign n450 = (~n447 & n448) | (~n447 & n449) | (n448 & n449);
  assign n451 = x2 | n450;
  assign n443 = x5 | x6;
  assign n444 = x3 | n443;
  assign n445 = (~x3 & n271) | (~x3 & n444) | (n271 & n444);
  assign n452 = x1 | n445;
  assign n453 = x2 & n452;
  assign n454 = n451 & ~n453;
  assign n457 = (x0 & n454) | (x0 & n456) | (n454 & n456);
  assign n436 = (x3 & x6) | (x3 & n89) | (x6 & n89);
  assign n437 = n89 | n436;
  assign n438 = ~n193 & n437;
  assign n439 = x1 & ~n438;
  assign n435 = x5 & n233;
  assign n440 = x2 & n435;
  assign n441 = x1 | n440;
  assign n442 = ~n439 & n441;
  assign n458 = (~x0 & n442) | (~x0 & n456) | (n442 & n456);
  assign n459 = n457 & n458;
  assign n661 = x1 & ~x7;
  assign n662 = (x0 & ~x8) | (x0 & n661) | (~x8 & n661);
  assign n663 = (x7 & x8) | (x7 & n661) | (x8 & n661);
  assign n664 = (x0 & x1) | (x0 & ~n663) | (x1 & ~n663);
  assign n665 = ~n662 & n664;
  assign n666 = x3 & ~n665;
  assign n667 = n188 & ~n192;
  assign n668 = x3 | n667;
  assign n669 = ~n666 & n668;
  assign n676 = (x5 & x6) | (x5 & n669) | (x6 & n669);
  assign n670 = x5 | x8;
  assign n671 = (~n10 & n197) | (~n10 & n670) | (n197 & n670);
  assign n672 = (x1 & x3) | (x1 & ~n671) | (x3 & ~n671);
  assign n673 = (x0 & ~x3) | (x0 & n672) | (~x3 & n672);
  assign n674 = (x0 & x1) | (x0 & ~n672) | (x1 & ~n672);
  assign n675 = n673 & ~n674;
  assign n677 = ~x6 & n675;
  assign n678 = (n669 & ~n676) | (n669 & n677) | (~n676 & n677);
  assign n717 = ~x2 & n678;
  assign n690 = (x0 & x3) | (x0 & ~x7) | (x3 & ~x7);
  assign n691 = (~x0 & x5) | (~x0 & x7) | (x5 & x7);
  assign n692 = n690 | n691;
  assign n696 = (x1 & x2) | (x1 & ~n692) | (x2 & ~n692);
  assign n693 = x3 & n538;
  assign n694 = (x0 & x1) | (x0 & n693) | (x1 & n693);
  assign n695 = ~x0 & n694;
  assign n697 = x2 & n695;
  assign n698 = (~x1 & n696) | (~x1 & n697) | (n696 & n697);
  assign n679 = x3 & n192;
  assign n680 = (n13 & n347) | (n13 & ~n679) | (n347 & ~n679);
  assign n681 = (x5 & x8) | (x5 & n680) | (x8 & n680);
  assign n682 = (x7 & ~x8) | (x7 & n681) | (~x8 & n681);
  assign n683 = (x5 & x7) | (x5 & ~n681) | (x7 & ~n681);
  assign n684 = n682 & ~n683;
  assign n685 = (x3 & x5) | (x3 & n537) | (x5 & n537);
  assign n686 = ~x3 & n685;
  assign n687 = ~x2 & n686;
  assign n688 = (x0 & x1) | (x0 & n687) | (x1 & n687);
  assign n689 = ~x0 & n688;
  assign n699 = (x6 & n684) | (x6 & n689) | (n684 & n689);
  assign n700 = ~n698 & n699;
  assign n701 = (x6 & n698) | (x6 & n700) | (n698 & n700);
  assign n702 = (x1 & x5) | (x1 & x6) | (x5 & x6);
  assign n703 = x2 & n702;
  assign n709 = (~x0 & x3) | (~x0 & n703) | (x3 & n703);
  assign n704 = (x1 & x2) | (x1 & x6) | (x2 & x6);
  assign n705 = (x2 & ~x5) | (x2 & n704) | (~x5 & n704);
  assign n706 = x2 & ~n705;
  assign n707 = n705 | n706;
  assign n708 = (~x2 & n706) | (~x2 & n707) | (n706 & n707);
  assign n710 = (x0 & x3) | (x0 & n708) | (x3 & n708);
  assign n711 = n709 & n710;
  assign n712 = (x2 & n26) | (x2 & n38) | (n26 & n38);
  assign n713 = ~x2 & n712;
  assign n714 = n711 | n713;
  assign n715 = (x7 & x8) | (x7 & n714) | (x8 & n714);
  assign n716 = (n188 & n714) | (n188 & ~n715) | (n714 & ~n715);
  assign n718 = n701 | n716;
  assign n719 = (n678 & ~n717) | (n678 & n718) | (~n717 & n718);
  assign n720 = n459 | n719;
  assign n721 = (n434 & n660) | (n434 & ~n720) | (n660 & ~n720);
  assign n722 = ~n434 & n721;
  assign y0   = n16;
  assign y1   = n49;
  assign y2   = n128;
  assign y3   = n244;
  assign y4   = n411;
  assign y5   = ~n722;
endmodule
