// IWLS benchmark module "MinMax9b" printed on Wed May 29 22:12:27 2002
module mm9b(\1 , \2 , \3 , \4 , \5 , \6 , \7 , \8 , \9 , \10 , \11 , \12 , \39 , \40 , \41 , \42 , \43 , \44 , \45 , \46 , \47 );
input
  \1 ,
  \2 ,
  \3 ,
  \4 ,
  \5 ,
  \6 ,
  \7 ,
  \8 ,
  \9 ,
  \10 ,
  \11 ,
  \12 ;
output
  \39 ,
  \40 ,
  \41 ,
  \42 ,
  \43 ,
  \44 ,
  \45 ,
  \46 ,
  \47 ;
reg
  \13 ,
  \14 ,
  \15 ,
  \16 ,
  \17 ,
  \18 ,
  \19 ,
  \20 ,
  \21 ,
  \22 ,
  \23 ,
  \24 ,
  \25 ,
  \26 ,
  \27 ,
  \28 ,
  \29 ,
  \30 ,
  \31 ,
  \32 ,
  \33 ,
  \34 ,
  \35 ,
  \36 ,
  \37 ,
  \38 ;
wire
  \48 ,
  \49 ,
  \50 ,
  \51 ,
  \52 ,
  \53 ,
  \54 ,
  \55 ,
  \56 ,
  \57 ,
  \58 ,
  \59 ,
  \60 ,
  \61 ,
  \62 ,
  \63 ,
  \64 ,
  \65 ,
  \66 ,
  \67 ,
  \68 ,
  \69 ,
  \70 ,
  \71 ,
  \72 ,
  \73 ,
  \74 ,
  \75 ,
  \76 ,
  \77 ,
  \78 ,
  \79 ,
  \80 ,
  \81 ,
  \82 ,
  \83 ,
  \84 ,
  \85 ,
  \86 ,
  \87 ,
  \88 ,
  \89 ,
  \90 ,
  \91 ,
  \92 ,
  \93 ,
  \94 ,
  \95 ,
  \96 ,
  \97 ,
  \98 ,
  \99 ,
  \100 ,
  \101 ,
  \102 ,
  \103 ,
  \104 ,
  \105 ,
  \106 ,
  \107 ,
  \108 ,
  \109 ,
  \110 ,
  \111 ,
  \112 ,
  \113 ,
  \114 ,
  \115 ,
  \116 ,
  \117 ,
  \118 ,
  \119 ,
  \120 ,
  \121 ,
  \122 ,
  \123 ,
  \124 ,
  \125 ,
  \126 ,
  \127 ,
  \128 ,
  \129 ,
  \130 ,
  \131 ,
  \132 ,
  \133 ,
  \134 ,
  \135 ,
  \136 ,
  \137 ,
  \138 ,
  \139 ,
  \140 ,
  \141 ,
  \142 ,
  \143 ,
  \144 ,
  \145 ,
  \146 ,
  \147 ,
  \148 ,
  \149 ,
  \150 ,
  \151 ,
  \152 ,
  \153 ,
  \154 ,
  \155 ,
  \156 ,
  \157 ,
  \158 ,
  \159 ,
  \160 ,
  \161 ,
  \162 ,
  \163 ,
  \164 ,
  \165 ,
  \166 ,
  \167 ,
  \168 ,
  \169 ,
  \170 ,
  \171 ,
  \172 ,
  \173 ,
  \174 ,
  \175 ,
  \176 ,
  \177 ,
  \178 ,
  \179 ,
  \180 ,
  \181 ,
  \182 ,
  \183 ,
  \184 ,
  \185 ,
  \186 ,
  \187 ,
  \188 ,
  \189 ,
  \190 ,
  \191 ,
  \192 ,
  \193 ,
  \194 ,
  \195 ,
  \196 ,
  \197 ,
  \198 ,
  \199 ,
  \200 ,
  \201 ,
  \202 ,
  \203 ,
  \204 ,
  \205 ,
  \206 ,
  \207 ,
  \208 ,
  \209 ,
  \210 ,
  \211 ,
  \212 ,
  \213 ,
  \214 ,
  \215 ,
  \216 ,
  \217 ,
  \218 ,
  \219 ,
  \[26] ,
  \220 ,
  \221 ,
  \222 ,
  \223 ,
  \224 ,
  \225 ,
  \226 ,
  \227 ,
  \228 ,
  \229 ,
  \[27] ,
  \230 ,
  \231 ,
  \232 ,
  \233 ,
  \234 ,
  \235 ,
  \236 ,
  \237 ,
  \238 ,
  \239 ,
  \[28] ,
  \240 ,
  \241 ,
  \242 ,
  \243 ,
  \244 ,
  \245 ,
  \246 ,
  \247 ,
  \248 ,
  \249 ,
  \[29] ,
  \250 ,
  \251 ,
  \252 ,
  \253 ,
  \254 ,
  \255 ,
  \256 ,
  \257 ,
  \258 ,
  \259 ,
  \260 ,
  \261 ,
  \262 ,
  \263 ,
  \264 ,
  \265 ,
  \266 ,
  \267 ,
  \268 ,
  \269 ,
  \270 ,
  \271 ,
  \272 ,
  \273 ,
  \274 ,
  \275 ,
  \276 ,
  \277 ,
  \278 ,
  \279 ,
  \280 ,
  \281 ,
  \282 ,
  \283 ,
  \284 ,
  \285 ,
  \286 ,
  \287 ,
  \288 ,
  \289 ,
  \290 ,
  \291 ,
  \292 ,
  \293 ,
  \294 ,
  \295 ,
  \296 ,
  \297 ,
  \298 ,
  \299 ,
  \[30] ,
  \[31] ,
  \[32] ,
  \[33] ,
  \[34] ,
  \300 ,
  \301 ,
  \302 ,
  \303 ,
  \304 ,
  \305 ,
  \306 ,
  \307 ,
  \308 ,
  \309 ,
  \[35] ,
  \310 ,
  \311 ,
  \312 ,
  \313 ,
  \314 ,
  \315 ,
  \316 ,
  \317 ,
  \318 ,
  \319 ,
  \[36] ,
  \320 ,
  \321 ,
  \322 ,
  \323 ,
  \324 ,
  \325 ,
  \326 ,
  \327 ,
  \328 ,
  \329 ,
  \[37] ,
  \330 ,
  \331 ,
  \332 ,
  \333 ,
  \334 ,
  \335 ,
  \336 ,
  \337 ,
  \338 ,
  \339 ,
  \[38] ,
  \340 ,
  \341 ,
  \342 ,
  \343 ,
  \344 ,
  \345 ,
  \346 ,
  \347 ,
  \348 ,
  \349 ,
  \[39] ,
  \350 ,
  \351 ,
  \352 ,
  \353 ,
  \354 ,
  \355 ,
  \356 ,
  \357 ,
  \358 ,
  \359 ,
  \360 ,
  \361 ,
  \362 ,
  \363 ,
  \364 ,
  \365 ,
  \366 ,
  \367 ,
  \368 ,
  \369 ,
  \370 ,
  \371 ,
  \372 ,
  \373 ,
  \374 ,
  \375 ,
  \376 ,
  \377 ,
  \378 ,
  \379 ,
  \380 ,
  \381 ,
  \382 ,
  \383 ,
  \384 ,
  \385 ,
  \386 ,
  \387 ,
  \388 ,
  \389 ,
  \390 ,
  \391 ,
  \392 ,
  \393 ,
  \394 ,
  \395 ,
  \396 ,
  \397 ,
  \398 ,
  \399 ,
  \[40] ,
  \[41] ,
  \[42] ,
  \[43] ,
  \[44] ,
  \400 ,
  \401 ,
  \402 ,
  \403 ,
  \404 ,
  \405 ,
  \406 ,
  \407 ,
  \408 ,
  \409 ,
  \[45] ,
  \410 ,
  \411 ,
  \412 ,
  \413 ,
  \414 ,
  \415 ,
  \416 ,
  \417 ,
  \418 ,
  \419 ,
  \[46] ,
  \420 ,
  \421 ,
  \422 ,
  \423 ,
  \424 ,
  \425 ,
  \426 ,
  \427 ,
  \428 ,
  \429 ,
  \[47] ,
  \430 ,
  \431 ,
  \432 ,
  \433 ,
  \434 ,
  \435 ,
  \436 ,
  \437 ,
  \438 ,
  \439 ,
  \[48] ,
  \440 ,
  \441 ,
  \442 ,
  \443 ,
  \444 ,
  \445 ,
  \446 ,
  \447 ,
  \448 ,
  \449 ,
  \[49] ,
  \450 ,
  \451 ,
  \452 ,
  \453 ,
  \454 ,
  \455 ,
  \456 ,
  \457 ,
  \458 ,
  \459 ,
  \460 ,
  \461 ,
  \462 ,
  \463 ,
  \464 ,
  \465 ,
  \466 ,
  \467 ,
  \468 ,
  \469 ,
  \470 ,
  \471 ,
  \472 ,
  \473 ,
  \474 ,
  \475 ,
  \476 ,
  \477 ,
  \478 ,
  \479 ,
  \480 ,
  \481 ,
  \482 ,
  \483 ,
  \484 ,
  \485 ,
  \486 ,
  \487 ,
  \488 ,
  \489 ,
  \490 ,
  \491 ,
  \492 ,
  \493 ,
  \494 ,
  \495 ,
  \496 ,
  \497 ,
  \498 ,
  \499 ,
  \[50] ,
  \[51] ,
  \[52] ,
  \[53] ,
  \[54] ,
  \500 ,
  \501 ,
  \502 ,
  \503 ,
  \504 ,
  \505 ,
  \506 ,
  \507 ,
  \508 ,
  \509 ,
  \[55] ,
  \510 ,
  \511 ,
  \512 ,
  \513 ,
  \514 ,
  \515 ,
  \516 ,
  \517 ,
  \518 ,
  \519 ,
  \[56] ,
  \520 ,
  \521 ,
  \522 ,
  \523 ,
  \524 ,
  \525 ,
  \526 ,
  \527 ,
  \528 ,
  \529 ,
  \[57] ,
  \530 ,
  \531 ,
  \532 ,
  \533 ,
  \534 ,
  \535 ,
  \536 ,
  \537 ,
  \538 ,
  \539 ,
  \[58] ,
  \540 ,
  \541 ,
  \542 ,
  \543 ,
  \544 ,
  \545 ,
  \546 ,
  \547 ,
  \548 ,
  \549 ,
  \[59] ,
  \550 ,
  \551 ,
  \552 ,
  \553 ,
  \554 ,
  \555 ,
  \556 ,
  \557 ,
  \558 ,
  \559 ,
  \560 ,
  \561 ,
  \562 ,
  \563 ,
  \564 ,
  \565 ,
  \566 ,
  \567 ,
  \568 ,
  \569 ,
  \570 ,
  \571 ,
  \572 ,
  \573 ,
  \574 ,
  \575 ,
  \576 ,
  \577 ,
  \578 ,
  \579 ,
  \580 ,
  \581 ,
  \582 ,
  \583 ,
  \584 ,
  \585 ,
  \586 ,
  \587 ,
  \588 ,
  \589 ,
  \590 ,
  \591 ,
  \592 ,
  \593 ,
  \594 ,
  \595 ,
  \596 ,
  \597 ,
  \598 ,
  \599 ,
  \[60] ,
  \600 ,
  \601 ,
  \602 ,
  \603 ,
  \604 ,
  \605 ,
  \606 ,
  \607 ,
  \608 ,
  \609 ,
  \610 ,
  \611 ,
  \612 ,
  \613 ,
  \614 ,
  \615 ,
  \616 ,
  \617 ,
  \618 ,
  \619 ,
  \620 ,
  \621 ,
  \622 ,
  \623 ,
  \624 ,
  \625 ,
  \626 ,
  \627 ,
  \628 ,
  \629 ,
  \630 ,
  \631 ,
  \632 ,
  \633 ,
  \634 ,
  \635 ,
  \636 ,
  \637 ,
  \638 ,
  \639 ,
  \640 ,
  \641 ,
  \642 ,
  \643 ,
  \644 ,
  \645 ,
  \646 ,
  \647 ,
  \648 ,
  \649 ,
  \650 ,
  \651 ,
  \652 ,
  \653 ,
  \654 ,
  \655 ,
  \656 ,
  \657 ,
  \658 ,
  \659 ,
  \660 ,
  \661 ,
  \662 ,
  \663 ,
  \664 ,
  \665 ,
  \666 ,
  \667 ,
  \668 ,
  \669 ,
  \670 ,
  \671 ,
  \672 ,
  \673 ,
  \674 ,
  \675 ,
  \676 ,
  \677 ,
  \678 ,
  \679 ,
  \680 ,
  \681 ,
  \682 ,
  \683 ,
  \684 ,
  \685 ,
  \686 ,
  \687 ,
  \688 ,
  \689 ,
  \690 ,
  \691 ,
  \692 ,
  \693 ,
  \694 ,
  \695 ,
  \696 ,
  \697 ,
  \698 ,
  \699 ,
  \700 ,
  \701 ,
  \702 ,
  \703 ,
  \704 ,
  \705 ,
  \706 ,
  \707 ,
  \708 ,
  \709 ,
  \710 ,
  \711 ,
  \712 ,
  \713 ,
  \714 ,
  \715 ,
  \716 ,
  \717 ,
  \718 ,
  \719 ,
  \720 ,
  \721 ,
  \722 ,
  \723 ,
  \724 ,
  \725 ,
  \726 ,
  \727 ,
  \728 ,
  \729 ,
  \730 ,
  \731 ,
  \732 ,
  \733 ,
  \734 ,
  \735 ,
  \736 ,
  \737 ,
  \738 ,
  \739 ,
  \740 ,
  \741 ,
  \742 ,
  \743 ,
  \744 ,
  \745 ,
  \746 ,
  \747 ,
  \748 ,
  \749 ,
  \750 ,
  \751 ,
  \752 ,
  \753 ,
  \754 ,
  \755 ,
  \756 ,
  \757 ,
  \758 ,
  \759 ,
  \760 ,
  \761 ,
  \762 ,
  \763 ,
  \764 ,
  \765 ,
  \766 ,
  \767 ,
  \768 ,
  \769 ,
  \770 ,
  \771 ,
  \772 ,
  \773 ,
  \774 ,
  \775 ,
  \776 ,
  \777 ,
  \778 ,
  \779 ,
  \780 ,
  \781 ,
  \782 ,
  \783 ,
  \784 ,
  \785 ,
  \786 ,
  \787 ,
  \788 ,
  \789 ,
  \790 ,
  \791 ,
  \792 ,
  \793 ,
  \794 ,
  \795 ,
  \796 ,
  \797 ,
  \798 ,
  \799 ,
  \800 ,
  \801 ,
  \802 ,
  \803 ,
  \804 ,
  \805 ,
  \806 ,
  \807 ,
  \808 ,
  \809 ,
  \810 ,
  \811 ,
  \812 ,
  \813 ,
  \814 ,
  \815 ,
  \816 ,
  \817 ,
  \818 ,
  \819 ,
  \820 ,
  \821 ,
  \822 ,
  \823 ,
  \824 ,
  \825 ,
  \826 ,
  \827 ,
  \828 ,
  \829 ,
  \830 ,
  \831 ,
  \832 ,
  \833 ,
  \834 ,
  \835 ,
  \836 ,
  \837 ,
  \838 ,
  \839 ,
  \840 ,
  \841 ,
  \842 ,
  \843 ,
  \844 ,
  \845 ,
  \846 ,
  \847 ,
  \848 ,
  \849 ,
  \850 ,
  \851 ,
  \852 ,
  \853 ,
  \854 ,
  \855 ,
  \856 ,
  \857 ,
  \858 ,
  \859 ,
  \860 ,
  \861 ,
  \862 ,
  \863 ,
  \864 ,
  \865 ,
  \866 ,
  \867 ,
  \868 ,
  \869 ,
  \870 ,
  \871 ,
  \872 ,
  \873 ,
  \874 ,
  \875 ,
  \876 ,
  \877 ,
  \878 ,
  \879 ,
  \880 ,
  \881 ,
  \882 ,
  \883 ,
  \884 ,
  \885 ,
  \886 ,
  \887 ,
  \888 ,
  \889 ,
  \890 ,
  \891 ,
  \892 ,
  \893 ,
  \894 ,
  \895 ,
  \896 ,
  \897 ,
  \898 ,
  \899 ,
  \900 ,
  \901 ,
  \902 ,
  \903 ,
  \904 ,
  \905 ,
  \906 ,
  \907 ,
  \908 ,
  \909 ,
  \910 ,
  \911 ,
  \912 ,
  \913 ,
  \914 ,
  \915 ,
  \916 ,
  \917 ,
  \918 ,
  \919 ,
  \920 ,
  \921 ,
  \922 ,
  \923 ,
  \924 ,
  \925 ,
  \926 ,
  \927 ,
  \928 ,
  \929 ,
  \930 ,
  \931 ,
  \932 ,
  \933 ,
  \934 ,
  \935 ,
  \936 ,
  \937 ,
  \938 ,
  \939 ,
  \940 ,
  \941 ,
  \942 ,
  \943 ,
  \944 ,
  \945 ,
  \946 ,
  \947 ,
  \948 ,
  \949 ,
  \950 ,
  \951 ,
  \952 ,
  \953 ,
  \954 ;
assign
  \39  = \[26] ,
  \40  = \[27] ,
  \41  = \[28] ,
  \42  = \[29] ,
  \43  = \[30] ,
  \44  = \[31] ,
  \45  = \[32] ,
  \46  = \[33] ,
  \47  = \[34] ,
  \48  = \532  | \531 ,
  \49  = \537  | \536 ,
  \50  = \542  | \541 ,
  \51  = \547  | \546 ,
  \52  = \552  | \551 ,
  \53  = \557  | \556 ,
  \54  = \562  | \561 ,
  \55  = \567  | \566 ,
  \56  = \572  | \571 ,
  \57  = \580  | \579 ,
  \58  = \588  | \587 ,
  \59  = \596  | \595 ,
  \60  = \604  | \603 ,
  \61  = \612  | \611 ,
  \62  = \620  | \619 ,
  \63  = \628  | \627 ,
  \64  = \636  | \635 ,
  \65  = \644  | \643 ,
  \66  = \652  | \651 ,
  \67  = \660  | \659 ,
  \68  = \668  | \667 ,
  \69  = \676  | \675 ,
  \70  = \684  | \683 ,
  \71  = \692  | \691 ,
  \72  = \700  | \699 ,
  \73  = \711  | \710 ,
  \74  = ~\75 ,
  \75  = \1 ,
  \76  = ~\77 ,
  \77  = ~\2 ,
  \78  = ~\79 ,
  \79  = \3 ,
  \80  = ~\81 ,
  \81  = \406  & \404 ,
  \82  = ~\83 ,
  \83  = \408  & \407 ,
  \84  = ~\85 ,
  \85  = (~\409  & \12 ) | (\409  & ~\12 ),
  \86  = ~\87 ,
  \87  = (~\410  & \11 ) | (\410  & ~\11 ),
  \88  = ~\89 ,
  \89  = (~\411  & \10 ) | (\411  & ~\10 ),
  \90  = ~\91 ,
  \91  = (~\412  & \9 ) | (\412  & ~\9 ),
  \92  = ~\93 ,
  \93  = (~\413  & \8 ) | (\413  & ~\8 ),
  \94  = ~\95 ,
  \95  = (~\414  & \7 ) | (\414  & ~\7 ),
  \96  = ~\97 ,
  \97  = (~\415  & \6 ) | (\415  & ~\6 ),
  \98  = ~\99 ,
  \99  = (~\416  & \5 ) | (\416  & ~\5 ),
  \100  = ~\101 ,
  \101  = (~\417  & \4 ) | (\417  & ~\4 ),
  \102  = ~\103 ,
  \103  = \418 ,
  \104  = ~\105 ,
  \105  = (~\419  & \12 ) | (\419  & ~\12 ),
  \106  = ~\107 ,
  \107  = (~\420  & \11 ) | (\420  & ~\11 ),
  \108  = ~\109 ,
  \109  = (~\421  & \10 ) | (\421  & ~\10 ),
  \110  = ~\111 ,
  \111  = (~\422  & \9 ) | (\422  & ~\9 ),
  \112  = ~\113 ,
  \113  = (~\423  & \8 ) | (\423  & ~\8 ),
  \114  = ~\115 ,
  \115  = (~\424  & \7 ) | (\424  & ~\7 ),
  \116  = ~\117 ,
  \117  = (~\425  & \6 ) | (\425  & ~\6 ),
  \118  = ~\119 ,
  \119  = (~\426  & \5 ) | (\426  & ~\5 ),
  \120  = ~\121 ,
  \121  = (~\427  & \4 ) | (\427  & ~\4 ),
  \122  = ~\123 ,
  \123  = \428 ,
  \124  = ~\125 ,
  \125  = ~\12 ,
  \126  = 0,
  \127  = 0,
  \128  = 0,
  \129  = 0,
  \130  = 0,
  \131  = 0,
  \132  = 0,
  \133  = 0,
  \134  = 0,
  \135  = 0,
  \136  = 0,
  \137  = 0,
  \138  = 0,
  \139  = 0,
  \140  = 0,
  \141  = 0,
  \142  = 0,
  \143  = 0,
  \144  = 0,
  \145  = \4 ,
  \146  = \5 ,
  \147  = \6 ,
  \148  = \7 ,
  \149  = \8 ,
  \150  = \9 ,
  \151  = \10 ,
  \152  = \11 ,
  \153  = \12 ,
  \154  = \13 ,
  \155  = \14 ,
  \156  = \15 ,
  \157  = \16 ,
  \158  = \17 ,
  \159  = \18 ,
  \160  = \19 ,
  \161  = \20 ,
  \162  = \21 ,
  \163  = 1,
  \164  = 1,
  \165  = 1,
  \166  = 1,
  \167  = 1,
  \168  = 1,
  \169  = 1,
  \170  = 1,
  \171  = 0,
  \172  = 0,
  \173  = 0,
  \174  = 0,
  \175  = 0,
  \176  = 0,
  \177  = 0,
  \178  = 0,
  \179  = 0,
  \180  = \21 ,
  \181  = \4 ,
  \182  = \5 ,
  \183  = \6 ,
  \184  = \7 ,
  \185  = \8 ,
  \186  = \9 ,
  \187  = \10 ,
  \188  = \11 ,
  \189  = \12 ,
  \190  = 0,
  \191  = 0,
  \192  = 0,
  \193  = 0,
  \194  = 0,
  \195  = 0,
  \196  = 0,
  \197  = 0,
  \198  = \12 ,
  \199  = 1,
  \200  = 1,
  \201  = 1,
  \202  = 1,
  \203  = 1,
  \204  = 1,
  \205  = 1,
  \206  = 1,
  \207  = 1,
  \208  = 0,
  \209  = 0,
  \210  = 0,
  \211  = 0,
  \212  = 0,
  \213  = 0,
  \214  = 0,
  \215  = 0,
  \216  = \13 ,
  \217  = \14 ,
  \218  = \15 ,
  \219  = \16 ,
  \[26]  = \463  | \462 ,
  \220  = \17 ,
  \221  = \18 ,
  \222  = \19 ,
  \223  = \20 ,
  \224  = \21 ,
  \225  = 1,
  \226  = 1,
  \227  = 1,
  \228  = 1,
  \229  = 1,
  \[27]  = \471  | \470 ,
  \230  = 1,
  \231  = 1,
  \232  = 1,
  \233  = \21  & \38 ,
  \234  = 1,
  \235  = 1,
  \236  = 1,
  \237  = 1,
  \238  = 1,
  \239  = 1,
  \[28]  = \479  | \478 ,
  \240  = 1,
  \241  = 1,
  \242  = 1,
  \243  = \22 ,
  \244  = \23 ,
  \245  = \24 ,
  \246  = \25 ,
  \247  = \26 ,
  \248  = \27 ,
  \249  = \28 ,
  \[29]  = \487  | \486 ,
  \250  = \29 ,
  \251  = 0,
  \252  = 0,
  \253  = 0,
  \254  = 0,
  \255  = 0,
  \256  = 0,
  \257  = 0,
  \258  = 0,
  \259  = 0,
  \260  = \21  | \38 ,
  \261  = \30 ,
  \262  = \31 ,
  \263  = \32 ,
  \264  = \33 ,
  \265  = \34 ,
  \266  = \35 ,
  \267  = \36 ,
  \268  = \37 ,
  \269  = \12 ,
  \270  = \11 ,
  \271  = \10 ,
  \272  = \9 ,
  \273  = \8 ,
  \274  = \7 ,
  \275  = \6 ,
  \276  = \5 ,
  \277  = 0,
  \278  = \4 ,
  \279  = \417 ,
  \280  = \416 ,
  \281  = \415 ,
  \282  = \414 ,
  \283  = \413 ,
  \284  = \412 ,
  \285  = \411 ,
  \286  = \410 ,
  \287  = \409 ,
  \288  = \4 ,
  \289  = \5 ,
  \290  = \6 ,
  \291  = \7 ,
  \292  = \8 ,
  \293  = \9 ,
  \294  = \10 ,
  \295  = \11 ,
  \296  = \12 ,
  \297  = \12 ,
  \298  = \11 ,
  \299  = \10 ,
  \[30]  = \495  | \494 ,
  \[31]  = \503  | \502 ,
  \[32]  = \511  | \510 ,
  \[33]  = \519  | \518 ,
  \[34]  = \527  | \526 ,
  \300  = \9 ,
  \301  = \8 ,
  \302  = \7 ,
  \303  = \6 ,
  \304  = \5 ,
  \305  = 0,
  \306  = \4 ,
  \307  = \4 ,
  \308  = \5 ,
  \309  = \6 ,
  \[35]  = \48 ,
  \310  = \7 ,
  \311  = \8 ,
  \312  = \9 ,
  \313  = \10 ,
  \314  = \11 ,
  \315  = \12 ,
  \316  = \427 ,
  \317  = \426 ,
  \318  = \425 ,
  \319  = \424 ,
  \[36]  = \49 ,
  \320  = \423 ,
  \321  = \422 ,
  \322  = \421 ,
  \323  = \420 ,
  \324  = \419 ,
  \325  = (\455  & \454 ) | ((\455  & \453 ) | (\454  & \453 )),
  \326  = (~\434  & (~\433  & \432 )) | ((~\434  & (\433  & ~\432 )) | ((\434  & (~\433  & ~\432 )) | (\434  & (\433  & \432 )))),
  \327  = (~\437  & (~\436  & \435 )) | ((~\437  & (\436  & ~\435 )) | ((\437  & (~\436  & ~\435 )) | (\437  & (\436  & \435 )))),
  \328  = (~\440  & (~\439  & \438 )) | ((~\440  & (\439  & ~\438 )) | ((\440  & (~\439  & ~\438 )) | (\440  & (\439  & \438 )))),
  \329  = (~\443  & (~\442  & \441 )) | ((~\443  & (\442  & ~\441 )) | ((\443  & (~\442  & ~\441 )) | (\443  & (\442  & \441 )))),
  \[37]  = \50 ,
  \330  = (~\446  & (~\445  & \444 )) | ((~\446  & (\445  & ~\444 )) | ((\446  & (~\445  & ~\444 )) | (\446  & (\445  & \444 )))),
  \331  = (~\449  & (~\448  & \447 )) | ((~\449  & (\448  & ~\447 )) | ((\449  & (~\448  & ~\447 )) | (\449  & (\448  & \447 )))),
  \332  = (~\452  & (~\451  & \450 )) | ((~\452  & (\451  & ~\450 )) | ((\452  & (~\451  & ~\450 )) | (\452  & (\451  & \450 )))),
  \333  = (~\455  & (~\454  & \453 )) | ((~\455  & (\454  & ~\453 )) | ((\455  & (~\454  & ~\453 )) | (\455  & (\454  & \453 )))),
  \334  = \325 ,
  \335  = \326 ,
  \336  = \327 ,
  \337  = \328 ,
  \338  = \329 ,
  \339  = \330 ,
  \[38]  = \51 ,
  \340  = \331 ,
  \341  = \332 ,
  \342  = \333 ,
  \343  = \430 ,
  \344  = \433 ,
  \345  = \436 ,
  \346  = \439 ,
  \347  = \442 ,
  \348  = \445 ,
  \349  = \448 ,
  \[39]  = \52 ,
  \350  = \451 ,
  \351  = \431 ,
  \352  = \434 ,
  \353  = \437 ,
  \354  = \440 ,
  \355  = \443 ,
  \356  = \446 ,
  \357  = \449 ,
  \358  = \452 ,
  \359  = \455 ,
  \360  = \454 ,
  \361  = 0,
  \362  = (~\361  & ~\37 ) | (\361  & \37 ),
  \363  = 0,
  \364  = (~\363  & ~\36 ) | (\363  & \36 ),
  \365  = \364  & \362 ,
  \366  = 0,
  \367  = (~\366  & ~\35 ) | (\366  & \35 ),
  \368  = \367  & \365 ,
  \369  = 0,
  \370  = (~\369  & ~\34 ) | (\369  & \34 ),
  \371  = \370  & \368 ,
  \372  = 0,
  \373  = (~\372  & ~\33 ) | (\372  & \33 ),
  \374  = \373  & \371 ,
  \375  = 0,
  \376  = (~\375  & ~\32 ) | (\375  & \32 ),
  \377  = \376  & \374 ,
  \378  = 0,
  \379  = (~\378  & ~\31 ) | (\378  & \31 ),
  \380  = \379  & \377 ,
  \381  = 0,
  \382  = (~\381  & ~\30 ) | (\381  & \30 ),
  \383  = \382  & \380 ,
  \384  = 1,
  \385  = (~\384  & ~\29 ) | (\384  & \29 ),
  \386  = \385  & \383 ,
  \387  = 1,
  \388  = (~\387  & ~\28 ) | (\387  & \28 ),
  \389  = \388  & \386 ,
  \390  = 1,
  \391  = (~\390  & ~\27 ) | (\390  & \27 ),
  \392  = \391  & \389 ,
  \393  = 1,
  \394  = (~\393  & ~\26 ) | (\393  & \26 ),
  \395  = \394  & \392 ,
  \396  = 1,
  \397  = (~\396  & ~\25 ) | (\396  & \25 ),
  \398  = \397  & \395 ,
  \399  = 1,
  \[40]  = \53 ,
  \[41]  = \54 ,
  \[42]  = \55 ,
  \[43]  = \56 ,
  \[44]  = \57 ,
  \400  = (~\399  & ~\24 ) | (\399  & \24 ),
  \401  = \400  & \398 ,
  \402  = 1,
  \403  = (~\402  & ~\23 ) | (\402  & \23 ),
  \404  = \403  & \401 ,
  \405  = 1,
  \406  = (~\405  & ~\22 ) | (\405  & \22 ),
  \407  = (~\21  & ~\38 ) | (\21  & \38 ),
  \408  = \954  & \952 ,
  \409  = \949  & \947 ,
  \[45]  = \58 ,
  \410  = \944  & \942 ,
  \411  = \939  & \937 ,
  \412  = \934  & \932 ,
  \413  = \929  & \927 ,
  \414  = \924  & \922 ,
  \415  = \919  & \917 ,
  \416  = \914  & \912 ,
  \417  = \909  & \907 ,
  \418  = \904  & \902 ,
  \419  = \875  & \873 ,
  \[46]  = \59 ,
  \420  = \870  & \868 ,
  \421  = \865  & \863 ,
  \422  = \860  & \858 ,
  \423  = \855  & \853 ,
  \424  = \850  & \848 ,
  \425  = \845  & \843 ,
  \426  = \840  & \838 ,
  \427  = \835  & \833 ,
  \428  = \830  & \828 ,
  \429  = 0,
  \[47]  = \60 ,
  \430  = \801  & \799 ,
  \431  = \796  & \794 ,
  \432  = (\431  & \430 ) | ((\431  & \429 ) | (\430  & \429 )),
  \433  = \791  & \789 ,
  \434  = \786  & \784 ,
  \435  = (\434  & \433 ) | ((\434  & \432 ) | (\433  & \432 )),
  \436  = \781  & \779 ,
  \437  = \776  & \774 ,
  \438  = (\437  & \436 ) | ((\437  & \435 ) | (\436  & \435 )),
  \439  = \771  & \769 ,
  \[48]  = \61 ,
  \440  = \766  & \764 ,
  \441  = (\440  & \439 ) | ((\440  & \438 ) | (\439  & \438 )),
  \442  = \761  & \759 ,
  \443  = \756  & \754 ,
  \444  = (\443  & \442 ) | ((\443  & \441 ) | (\442  & \441 )),
  \445  = \751  & \749 ,
  \446  = \746  & \744 ,
  \447  = (\446  & \445 ) | ((\446  & \444 ) | (\445  & \444 )),
  \448  = \741  & \739 ,
  \449  = \736  & \734 ,
  \[49]  = \62 ,
  \450  = (\449  & \448 ) | ((\449  & \447 ) | (\448  & \447 )),
  \451  = \731  & \729 ,
  \452  = \726  & \724 ,
  \453  = (\452  & \451 ) | ((\452  & \450 ) | (\451  & \450 )),
  \454  = \721  & \719 ,
  \455  = \716  & \714 ,
  \456  = \335  & \78 ,
  \457  = \181  & \79 ,
  \458  = \457  | \456 ,
  \459  = \458  & \76 ,
  \460  = \154  & \77 ,
  \461  = \460  | \459 ,
  \462  = \461  & \74 ,
  \463  = \127  & \75 ,
  \464  = \336  & \78 ,
  \465  = \182  & \79 ,
  \466  = \465  | \464 ,
  \467  = \466  & \76 ,
  \468  = \155  & \77 ,
  \469  = \468  | \467 ,
  \470  = \469  & \74 ,
  \471  = \128  & \75 ,
  \472  = \337  & \78 ,
  \473  = \183  & \79 ,
  \474  = \473  | \472 ,
  \475  = \474  & \76 ,
  \476  = \156  & \77 ,
  \477  = \476  | \475 ,
  \478  = \477  & \74 ,
  \479  = \129  & \75 ,
  \480  = \338  & \78 ,
  \481  = \184  & \79 ,
  \482  = \481  | \480 ,
  \483  = \482  & \76 ,
  \484  = \157  & \77 ,
  \485  = \484  | \483 ,
  \486  = \485  & \74 ,
  \487  = \130  & \75 ,
  \488  = \339  & \78 ,
  \489  = \185  & \79 ,
  \490  = \489  | \488 ,
  \491  = \490  & \76 ,
  \492  = \158  & \77 ,
  \493  = \492  | \491 ,
  \494  = \493  & \74 ,
  \495  = \131  & \75 ,
  \496  = \340  & \78 ,
  \497  = \186  & \79 ,
  \498  = \497  | \496 ,
  \499  = \498  & \76 ,
  \[50]  = \63 ,
  \[51]  = \64 ,
  \[52]  = \65 ,
  \[53]  = \66 ,
  \[54]  = \67 ,
  \500  = \159  & \77 ,
  \501  = \500  | \499 ,
  \502  = \501  & \74 ,
  \503  = \132  & \75 ,
  \504  = \341  & \78 ,
  \505  = \187  & \79 ,
  \506  = \505  | \504 ,
  \507  = \506  & \76 ,
  \508  = \160  & \77 ,
  \509  = \508  | \507 ,
  \[55]  = \68 ,
  \510  = \509  & \74 ,
  \511  = \133  & \75 ,
  \512  = \342  & \78 ,
  \513  = \188  & \79 ,
  \514  = \513  | \512 ,
  \515  = \514  & \76 ,
  \516  = \161  & \77 ,
  \517  = \516  | \515 ,
  \518  = \517  & \74 ,
  \519  = \134  & \75 ,
  \[56]  = \69 ,
  \520  = \334  & \78 ,
  \521  = \189  & \79 ,
  \522  = \521  | \520 ,
  \523  = \522  & \76 ,
  \524  = \162  & \77 ,
  \525  = \524  | \523 ,
  \526  = \525  & \74 ,
  \527  = \135  & \75 ,
  \528  = \145  & \76 ,
  \529  = \216  & \77 ,
  \[57]  = \70 ,
  \530  = \529  | \528 ,
  \531  = \530  & \74 ,
  \532  = \136  & \75 ,
  \533  = \146  & \76 ,
  \534  = \217  & \77 ,
  \535  = \534  | \533 ,
  \536  = \535  & \74 ,
  \537  = \137  & \75 ,
  \538  = \147  & \76 ,
  \539  = \218  & \77 ,
  \[58]  = \71 ,
  \540  = \539  | \538 ,
  \541  = \540  & \74 ,
  \542  = \138  & \75 ,
  \543  = \148  & \76 ,
  \544  = \219  & \77 ,
  \545  = \544  | \543 ,
  \546  = \545  & \74 ,
  \547  = \139  & \75 ,
  \548  = \149  & \76 ,
  \549  = \220  & \77 ,
  \[59]  = \72 ,
  \550  = \549  | \548 ,
  \551  = \550  & \74 ,
  \552  = \140  & \75 ,
  \553  = \150  & \76 ,
  \554  = \221  & \77 ,
  \555  = \554  | \553 ,
  \556  = \555  & \74 ,
  \557  = \141  & \75 ,
  \558  = \151  & \76 ,
  \559  = \222  & \77 ,
  \560  = \559  | \558 ,
  \561  = \560  & \74 ,
  \562  = \142  & \75 ,
  \563  = \152  & \76 ,
  \564  = \223  & \77 ,
  \565  = \564  | \563 ,
  \566  = \565  & \74 ,
  \567  = \143  & \75 ,
  \568  = \153  & \76 ,
  \569  = \224  & \77 ,
  \570  = \569  | \568 ,
  \571  = \570  & \74 ,
  \572  = \144  & \75 ,
  \573  = \351  & \78 ,
  \574  = \225  & \79 ,
  \575  = \574  | \573 ,
  \576  = \575  & \76 ,
  \577  = \199  & \77 ,
  \578  = \577  | \576 ,
  \579  = \578  & \74 ,
  \580  = \163  & \75 ,
  \581  = \352  & \78 ,
  \582  = \226  & \79 ,
  \583  = \582  | \581 ,
  \584  = \583  & \76 ,
  \585  = \200  & \77 ,
  \586  = \585  | \584 ,
  \587  = \586  & \74 ,
  \588  = \164  & \75 ,
  \589  = \353  & \78 ,
  \590  = \227  & \79 ,
  \591  = \590  | \589 ,
  \592  = \591  & \76 ,
  \593  = \201  & \77 ,
  \594  = \593  | \592 ,
  \595  = \594  & \74 ,
  \596  = \165  & \75 ,
  \597  = \354  & \78 ,
  \598  = \228  & \79 ,
  \599  = \598  | \597 ,
  \[60]  = \73 ,
  \600  = \599  & \76 ,
  \601  = \202  & \77 ,
  \602  = \601  | \600 ,
  \603  = \602  & \74 ,
  \604  = \166  & \75 ,
  \605  = \355  & \78 ,
  \606  = \229  & \79 ,
  \607  = \606  | \605 ,
  \608  = \607  & \76 ,
  \609  = \203  & \77 ,
  \610  = \609  | \608 ,
  \611  = \610  & \74 ,
  \612  = \167  & \75 ,
  \613  = \356  & \78 ,
  \614  = \230  & \79 ,
  \615  = \614  | \613 ,
  \616  = \615  & \76 ,
  \617  = \204  & \77 ,
  \618  = \617  | \616 ,
  \619  = \618  & \74 ,
  \620  = \168  & \75 ,
  \621  = \357  & \78 ,
  \622  = \231  & \79 ,
  \623  = \622  | \621 ,
  \624  = \623  & \76 ,
  \625  = \205  & \77 ,
  \626  = \625  | \624 ,
  \627  = \626  & \74 ,
  \628  = \169  & \75 ,
  \629  = \358  & \78 ,
  \630  = \232  & \79 ,
  \631  = \630  | \629 ,
  \632  = \631  & \76 ,
  \633  = \206  & \77 ,
  \634  = \633  | \632 ,
  \635  = \634  & \74 ,
  \636  = \170  & \75 ,
  \637  = \343  & \78 ,
  \638  = \208  & \79 ,
  \639  = \638  | \637 ,
  \640  = \639  & \76 ,
  \641  = \190  & \77 ,
  \642  = \641  | \640 ,
  \643  = \642  & \74 ,
  \644  = \171  & \75 ,
  \645  = \344  & \78 ,
  \646  = \209  & \79 ,
  \647  = \646  | \645 ,
  \648  = \647  & \76 ,
  \649  = \191  & \77 ,
  \650  = \649  | \648 ,
  \651  = \650  & \74 ,
  \652  = \172  & \75 ,
  \653  = \345  & \78 ,
  \654  = \210  & \79 ,
  \655  = \654  | \653 ,
  \656  = \655  & \76 ,
  \657  = \192  & \77 ,
  \658  = \657  | \656 ,
  \659  = \658  & \74 ,
  \660  = \173  & \75 ,
  \661  = \346  & \78 ,
  \662  = \211  & \79 ,
  \663  = \662  | \661 ,
  \664  = \663  & \76 ,
  \665  = \193  & \77 ,
  \666  = \665  | \664 ,
  \667  = \666  & \74 ,
  \668  = \174  & \75 ,
  \669  = \347  & \78 ,
  \670  = \212  & \79 ,
  \671  = \670  | \669 ,
  \672  = \671  & \76 ,
  \673  = \194  & \77 ,
  \674  = \673  | \672 ,
  \675  = \674  & \74 ,
  \676  = \175  & \75 ,
  \677  = \348  & \78 ,
  \678  = \213  & \79 ,
  \679  = \678  | \677 ,
  \680  = \679  & \76 ,
  \681  = \195  & \77 ,
  \682  = \681  | \680 ,
  \683  = \682  & \74 ,
  \684  = \176  & \75 ,
  \685  = \349  & \78 ,
  \686  = \214  & \79 ,
  \687  = \686  | \685 ,
  \688  = \687  & \76 ,
  \689  = \196  & \77 ,
  \690  = \689  | \688 ,
  \691  = \690  & \74 ,
  \692  = \177  & \75 ,
  \693  = \350  & \78 ,
  \694  = \215  & \79 ,
  \695  = \694  | \693 ,
  \696  = \695  & \76 ,
  \697  = \197  & \77 ,
  \698  = \697  | \696 ,
  \699  = \698  & \74 ,
  \700  = \178  & \75 ,
  \701  = \359  & \124 ,
  \702  = \360  & \125 ,
  \703  = \702  | \701 ,
  \704  = \703  & \78 ,
  \705  = \198  & \79 ,
  \706  = \705  | \704 ,
  \707  = \706  & \76 ,
  \708  = \180  & \77 ,
  \709  = \708  | \707 ,
  \710  = \709  & \74 ,
  \711  = \179  & \75 ,
  \712  = \315  & \122 ,
  \713  = \324  & \123 ,
  \714  = \713  | \712 ,
  \715  = \78  & \76 ,
  \716  = \715  & \74 ,
  \717  = \287  & \102 ,
  \718  = \296  & \103 ,
  \719  = \718  | \717 ,
  \720  = \78  & \76 ,
  \721  = \720  & \74 ,
  \722  = \314  & \122 ,
  \723  = \323  & \123 ,
  \724  = \723  | \722 ,
  \725  = \78  & \76 ,
  \726  = \725  & \74 ,
  \727  = \286  & \102 ,
  \728  = \295  & \103 ,
  \729  = \728  | \727 ,
  \730  = \78  & \76 ,
  \731  = \730  & \74 ,
  \732  = \313  & \122 ,
  \733  = \322  & \123 ,
  \734  = \733  | \732 ,
  \735  = \78  & \76 ,
  \736  = \735  & \74 ,
  \737  = \285  & \102 ,
  \738  = \294  & \103 ,
  \739  = \738  | \737 ,
  \740  = \78  & \76 ,
  \741  = \740  & \74 ,
  \742  = \312  & \122 ,
  \743  = \321  & \123 ,
  \744  = \743  | \742 ,
  \745  = \78  & \76 ,
  \746  = \745  & \74 ,
  \747  = \284  & \102 ,
  \748  = \293  & \103 ,
  \749  = \748  | \747 ,
  \750  = \78  & \76 ,
  \751  = \750  & \74 ,
  \752  = \311  & \122 ,
  \753  = \320  & \123 ,
  \754  = \753  | \752 ,
  \755  = \78  & \76 ,
  \756  = \755  & \74 ,
  \757  = \283  & \102 ,
  \758  = \292  & \103 ,
  \759  = \758  | \757 ,
  \760  = \78  & \76 ,
  \761  = \760  & \74 ,
  \762  = \310  & \122 ,
  \763  = \319  & \123 ,
  \764  = \763  | \762 ,
  \765  = \78  & \76 ,
  \766  = \765  & \74 ,
  \767  = \282  & \102 ,
  \768  = \291  & \103 ,
  \769  = \768  | \767 ,
  \770  = \78  & \76 ,
  \771  = \770  & \74 ,
  \772  = \309  & \122 ,
  \773  = \318  & \123 ,
  \774  = \773  | \772 ,
  \775  = \78  & \76 ,
  \776  = \775  & \74 ,
  \777  = \281  & \102 ,
  \778  = \290  & \103 ,
  \779  = \778  | \777 ,
  \780  = \78  & \76 ,
  \781  = \780  & \74 ,
  \782  = \308  & \122 ,
  \783  = \317  & \123 ,
  \784  = \783  | \782 ,
  \785  = \78  & \76 ,
  \786  = \785  & \74 ,
  \787  = \280  & \102 ,
  \788  = \289  & \103 ,
  \789  = \788  | \787 ,
  \790  = \78  & \76 ,
  \791  = \790  & \74 ,
  \792  = \307  & \122 ,
  \793  = \316  & \123 ,
  \794  = \793  | \792 ,
  \795  = \78  & \76 ,
  \796  = \795  & \74 ,
  \797  = \279  & \102 ,
  \798  = \288  & \103 ,
  \799  = \798  | \797 ,
  \800  = \78  & \76 ,
  \801  = \800  & \74 ,
  \802  = \305  & \120 ,
  \803  = \306  & \121 ,
  \804  = \803  | \802 ,
  \805  = \804  & \118 ,
  \806  = \304  & \119 ,
  \807  = \806  | \805 ,
  \808  = \807  & \116 ,
  \809  = \303  & \117 ,
  \810  = \809  | \808 ,
  \811  = \810  & \114 ,
  \812  = \302  & \115 ,
  \813  = \812  | \811 ,
  \814  = \813  & \112 ,
  \815  = \301  & \113 ,
  \816  = \815  | \814 ,
  \817  = \816  & \110 ,
  \818  = \300  & \111 ,
  \819  = \818  | \817 ,
  \820  = \819  & \108 ,
  \821  = \299  & \109 ,
  \822  = \821  | \820 ,
  \823  = \822  & \106 ,
  \824  = \298  & \107 ,
  \825  = \824  | \823 ,
  \826  = \825  & \104 ,
  \827  = \297  & \105 ,
  \828  = \827  | \826 ,
  \829  = \78  & \76 ,
  \830  = \829  & \74 ,
  \831  = \243  & \82 ,
  \832  = \234  & \83 ,
  \833  = \832  | \831 ,
  \834  = \78  & \76 ,
  \835  = \834  & \74 ,
  \836  = \244  & \82 ,
  \837  = \235  & \83 ,
  \838  = \837  | \836 ,
  \839  = \78  & \76 ,
  \840  = \839  & \74 ,
  \841  = \245  & \82 ,
  \842  = \236  & \83 ,
  \843  = \842  | \841 ,
  \844  = \78  & \76 ,
  \845  = \844  & \74 ,
  \846  = \246  & \82 ,
  \847  = \237  & \83 ,
  \848  = \847  | \846 ,
  \849  = \78  & \76 ,
  \850  = \849  & \74 ,
  \851  = \247  & \82 ,
  \852  = \238  & \83 ,
  \853  = \852  | \851 ,
  \854  = \78  & \76 ,
  \855  = \854  & \74 ,
  \856  = \248  & \82 ,
  \857  = \239  & \83 ,
  \858  = \857  | \856 ,
  \859  = \78  & \76 ,
  \860  = \859  & \74 ,
  \861  = \249  & \82 ,
  \862  = \240  & \83 ,
  \863  = \862  | \861 ,
  \864  = \78  & \76 ,
  \865  = \864  & \74 ,
  \866  = \250  & \82 ,
  \867  = \241  & \83 ,
  \868  = \867  | \866 ,
  \869  = \78  & \76 ,
  \870  = \869  & \74 ,
  \871  = \233  & \82 ,
  \872  = \242  & \83 ,
  \873  = \872  | \871 ,
  \874  = \78  & \76 ,
  \875  = \874  & \74 ,
  \876  = \277  & \100 ,
  \877  = \278  & \101 ,
  \878  = \877  | \876 ,
  \879  = \878  & \98 ,
  \880  = \276  & \99 ,
  \881  = \880  | \879 ,
  \882  = \881  & \96 ,
  \883  = \275  & \97 ,
  \884  = \883  | \882 ,
  \885  = \884  & \94 ,
  \886  = \274  & \95 ,
  \887  = \886  | \885 ,
  \888  = \887  & \92 ,
  \889  = \273  & \93 ,
  \890  = \889  | \888 ,
  \891  = \890  & \90 ,
  \892  = \272  & \91 ,
  \893  = \892  | \891 ,
  \894  = \893  & \88 ,
  \895  = \271  & \89 ,
  \896  = \895  | \894 ,
  \897  = \896  & \86 ,
  \898  = \270  & \87 ,
  \899  = \898  | \897 ,
  \900  = \899  & \84 ,
  \901  = \269  & \85 ,
  \902  = \901  | \900 ,
  \903  = \78  & \76 ,
  \904  = \903  & \74 ,
  \905  = \261  & \82 ,
  \906  = \251  & \83 ,
  \907  = \906  | \905 ,
  \908  = \78  & \76 ,
  \909  = \908  & \74 ,
  \910  = \262  & \82 ,
  \911  = \252  & \83 ,
  \912  = \911  | \910 ,
  \913  = \78  & \76 ,
  \914  = \913  & \74 ,
  \915  = \263  & \82 ,
  \916  = \253  & \83 ,
  \917  = \916  | \915 ,
  \918  = \78  & \76 ,
  \919  = \918  & \74 ,
  \920  = \264  & \82 ,
  \921  = \254  & \83 ,
  \922  = \921  | \920 ,
  \923  = \78  & \76 ,
  \924  = \923  & \74 ,
  \925  = \265  & \82 ,
  \926  = \255  & \83 ,
  \927  = \926  | \925 ,
  \928  = \78  & \76 ,
  \929  = \928  & \74 ,
  \930  = \266  & \82 ,
  \931  = \256  & \83 ,
  \932  = \931  | \930 ,
  \933  = \78  & \76 ,
  \934  = \933  & \74 ,
  \935  = \267  & \82 ,
  \936  = \257  & \83 ,
  \937  = \936  | \935 ,
  \938  = \78  & \76 ,
  \939  = \938  & \74 ,
  \940  = \268  & \82 ,
  \941  = \258  & \83 ,
  \942  = \941  | \940 ,
  \943  = \78  & \76 ,
  \944  = \943  & \74 ,
  \945  = \260  & \82 ,
  \946  = \259  & \83 ,
  \947  = \946  | \945 ,
  \948  = \78  & \76 ,
  \949  = \948  & \74 ,
  \950  = \126  & \80 ,
  \951  = \207  & \81 ,
  \952  = \951  | \950 ,
  \953  = \78  & \76 ,
  \954  = \953  & \74 ;
always begin
  \13  = \[35] ;
  \14  = \[36] ;
  \15  = \[37] ;
  \16  = \[38] ;
  \17  = \[39] ;
  \18  = \[40] ;
  \19  = \[41] ;
  \20  = \[42] ;
  \21  = \[43] ;
  \22  = \[44] ;
  \23  = \[45] ;
  \24  = \[46] ;
  \25  = \[47] ;
  \26  = \[48] ;
  \27  = \[49] ;
  \28  = \[50] ;
  \29  = \[51] ;
  \30  = \[52] ;
  \31  = \[53] ;
  \32  = \[54] ;
  \33  = \[55] ;
  \34  = \[56] ;
  \35  = \[57] ;
  \36  = \[58] ;
  \37  = \[59] ;
  \38  = \[60] ;
end
initial begin
  \13  = 0;
  \14  = 0;
  \15  = 0;
  \16  = 0;
  \17  = 0;
  \18  = 0;
  \19  = 0;
  \20  = 0;
  \21  = 0;
  \22  = 1;
  \23  = 1;
  \24  = 1;
  \25  = 1;
  \26  = 1;
  \27  = 1;
  \28  = 1;
  \29  = 1;
  \30  = 0;
  \31  = 0;
  \32  = 0;
  \33  = 0;
  \34  = 0;
  \35  = 0;
  \36  = 0;
  \37  = 0;
  \38  = 0;
end
endmodule

