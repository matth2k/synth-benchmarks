// IWLS benchmark module "MinMax30" printed on Wed May 29 22:06:07 2002
module mm30a(\1 , \2 , \3 , \4 , \5 , \6 , \7 , \8 , \9 , \10 , \11 , \12 , \13 , \14 , \15 , \16 , \17 , \18 , \19 , \20 , \21 , \22 , \23 , \24 , \25 , \26 , \27 , \28 , \29 , \30 , \31 , \32 , \33 , \124 , \125 , \126 , \127 , \128 , \129 , \130 , \131 , \132 , \133 , \134 , \135 , \136 , \137 , \138 , \139 , \140 , \141 , \142 , \143 , \144 , \145 , \146 , \147 , \148 , \149 , \150 , \151 , \152 , \153 );
input
  \1 ,
  \2 ,
  \3 ,
  \4 ,
  \5 ,
  \6 ,
  \7 ,
  \8 ,
  \9 ,
  \10 ,
  \11 ,
  \12 ,
  \13 ,
  \14 ,
  \15 ,
  \16 ,
  \17 ,
  \18 ,
  \19 ,
  \20 ,
  \21 ,
  \22 ,
  \23 ,
  \24 ,
  \25 ,
  \26 ,
  \27 ,
  \28 ,
  \29 ,
  \30 ,
  \31 ,
  \32 ,
  \33 ;
output
  \124 ,
  \125 ,
  \126 ,
  \127 ,
  \128 ,
  \129 ,
  \130 ,
  \131 ,
  \132 ,
  \133 ,
  \134 ,
  \135 ,
  \136 ,
  \137 ,
  \138 ,
  \139 ,
  \140 ,
  \141 ,
  \142 ,
  \143 ,
  \144 ,
  \145 ,
  \146 ,
  \147 ,
  \148 ,
  \149 ,
  \150 ,
  \151 ,
  \152 ,
  \153 ;
reg
  \34 ,
  \35 ,
  \36 ,
  \37 ,
  \38 ,
  \39 ,
  \40 ,
  \41 ,
  \42 ,
  \43 ,
  \44 ,
  \45 ,
  \46 ,
  \47 ,
  \48 ,
  \49 ,
  \50 ,
  \51 ,
  \52 ,
  \53 ,
  \54 ,
  \55 ,
  \56 ,
  \57 ,
  \58 ,
  \59 ,
  \60 ,
  \61 ,
  \62 ,
  \63 ,
  \64 ,
  \65 ,
  \66 ,
  \67 ,
  \68 ,
  \69 ,
  \70 ,
  \71 ,
  \72 ,
  \73 ,
  \74 ,
  \75 ,
  \76 ,
  \77 ,
  \78 ,
  \79 ,
  \80 ,
  \81 ,
  \82 ,
  \83 ,
  \84 ,
  \85 ,
  \86 ,
  \87 ,
  \88 ,
  \89 ,
  \90 ,
  \91 ,
  \92 ,
  \93 ,
  \94 ,
  \95 ,
  \96 ,
  \97 ,
  \98 ,
  \99 ,
  \100 ,
  \101 ,
  \102 ,
  \103 ,
  \104 ,
  \105 ,
  \106 ,
  \107 ,
  \108 ,
  \109 ,
  \110 ,
  \111 ,
  \112 ,
  \113 ,
  \114 ,
  \115 ,
  \116 ,
  \117 ,
  \118 ,
  \119 ,
  \120 ,
  \121 ,
  \122 ,
  \123 ;
wire
  \650 ,
  \651 ,
  \652 ,
  \653 ,
  \654 ,
  \655 ,
  \656 ,
  \657 ,
  \658 ,
  \659 ,
  \660 ,
  \661 ,
  \662 ,
  \663 ,
  \664 ,
  \665 ,
  \666 ,
  \667 ,
  \668 ,
  \669 ,
  \670 ,
  \671 ,
  \672 ,
  \673 ,
  \674 ,
  \675 ,
  \676 ,
  \677 ,
  \678 ,
  \679 ,
  \680 ,
  \681 ,
  \682 ,
  \683 ,
  \684 ,
  \685 ,
  \686 ,
  \687 ,
  \688 ,
  \689 ,
  \690 ,
  \691 ,
  \692 ,
  \693 ,
  \694 ,
  \695 ,
  \696 ,
  \697 ,
  \698 ,
  \699 ,
  \700 ,
  \701 ,
  \702 ,
  \703 ,
  \704 ,
  \705 ,
  \706 ,
  \707 ,
  \708 ,
  \709 ,
  \710 ,
  \711 ,
  \712 ,
  \713 ,
  \714 ,
  \715 ,
  \716 ,
  \717 ,
  \718 ,
  \719 ,
  \720 ,
  \721 ,
  \722 ,
  \723 ,
  \724 ,
  \725 ,
  \726 ,
  \727 ,
  \728 ,
  \729 ,
  \730 ,
  \731 ,
  \732 ,
  \733 ,
  \734 ,
  \735 ,
  \736 ,
  \737 ,
  \738 ,
  \739 ,
  \740 ,
  \741 ,
  \742 ,
  \743 ,
  \744 ,
  \745 ,
  \746 ,
  \747 ,
  \748 ,
  \749 ,
  \750 ,
  \751 ,
  \752 ,
  \753 ,
  \754 ,
  \755 ,
  \756 ,
  \757 ,
  \758 ,
  \759 ,
  \760 ,
  \761 ,
  \762 ,
  \763 ,
  \764 ,
  \765 ,
  \766 ,
  \767 ,
  \768 ,
  \769 ,
  \770 ,
  \771 ,
  \772 ,
  \773 ,
  \774 ,
  \775 ,
  \776 ,
  \777 ,
  \778 ,
  \779 ,
  \780 ,
  \781 ,
  \782 ,
  \783 ,
  \784 ,
  \785 ,
  \786 ,
  \787 ,
  \788 ,
  \789 ,
  \790 ,
  \791 ,
  \792 ,
  \793 ,
  \794 ,
  \795 ,
  \796 ,
  \797 ,
  \798 ,
  \799 ,
  \800 ,
  \801 ,
  \802 ,
  \803 ,
  \804 ,
  \805 ,
  \806 ,
  \807 ,
  \808 ,
  \809 ,
  \810 ,
  \811 ,
  \812 ,
  \813 ,
  \814 ,
  \815 ,
  \816 ,
  \817 ,
  \818 ,
  \819 ,
  \820 ,
  \821 ,
  \822 ,
  \823 ,
  \824 ,
  \825 ,
  \826 ,
  \827 ,
  \828 ,
  \829 ,
  \830 ,
  \831 ,
  \832 ,
  \833 ,
  \834 ,
  \835 ,
  \836 ,
  \837 ,
  \838 ,
  \839 ,
  \840 ,
  \841 ,
  \842 ,
  \843 ,
  \844 ,
  \845 ,
  \846 ,
  \847 ,
  \848 ,
  \849 ,
  \850 ,
  \851 ,
  \852 ,
  \853 ,
  \854 ,
  \855 ,
  \856 ,
  \857 ,
  \858 ,
  \859 ,
  \860 ,
  \861 ,
  \862 ,
  \863 ,
  \864 ,
  \865 ,
  \866 ,
  \867 ,
  \868 ,
  \869 ,
  \870 ,
  \871 ,
  \872 ,
  \873 ,
  \874 ,
  \875 ,
  \876 ,
  \877 ,
  \878 ,
  \879 ,
  \880 ,
  \881 ,
  \882 ,
  \883 ,
  \884 ,
  \885 ,
  \886 ,
  \887 ,
  \888 ,
  \889 ,
  \890 ,
  \891 ,
  \892 ,
  \893 ,
  \894 ,
  \895 ,
  \896 ,
  \[200] ,
  \897 ,
  \898 ,
  \899 ,
  \[201] ,
  \[202] ,
  \[203] ,
  \[204] ,
  \[205] ,
  \[206] ,
  \900 ,
  \901 ,
  \902 ,
  \903 ,
  \904 ,
  \905 ,
  \906 ,
  \[207] ,
  \907 ,
  \908 ,
  \909 ,
  \910 ,
  \911 ,
  \912 ,
  \913 ,
  \914 ,
  \915 ,
  \916 ,
  \[208] ,
  \917 ,
  \918 ,
  \919 ,
  \920 ,
  \921 ,
  \922 ,
  \923 ,
  \924 ,
  \925 ,
  \926 ,
  \[209] ,
  \927 ,
  \928 ,
  \929 ,
  \930 ,
  \931 ,
  \932 ,
  \933 ,
  \934 ,
  \935 ,
  \936 ,
  \937 ,
  \938 ,
  \939 ,
  \940 ,
  \941 ,
  \942 ,
  \943 ,
  \944 ,
  \945 ,
  \946 ,
  \947 ,
  \948 ,
  \949 ,
  \950 ,
  \951 ,
  \952 ,
  \953 ,
  \954 ,
  \955 ,
  \956 ,
  \957 ,
  \958 ,
  \959 ,
  \960 ,
  \961 ,
  \962 ,
  \963 ,
  \964 ,
  \965 ,
  \966 ,
  \967 ,
  \968 ,
  \969 ,
  \970 ,
  \971 ,
  \972 ,
  \973 ,
  \974 ,
  \975 ,
  \976 ,
  \977 ,
  \978 ,
  \979 ,
  \980 ,
  \981 ,
  \982 ,
  \983 ,
  \984 ,
  \985 ,
  \986 ,
  \987 ,
  \988 ,
  \989 ,
  \990 ,
  \991 ,
  \992 ,
  \993 ,
  \994 ,
  \995 ,
  \996 ,
  \997 ,
  \998 ,
  \999 ,
  \[90] ,
  \[91] ,
  \[92] ,
  \[93] ,
  \[94] ,
  \[95] ,
  \[96] ,
  \[97] ,
  \[98] ,
  \[99] ,
  \1000 ,
  \1001 ,
  \1002 ,
  \1003 ,
  \1004 ,
  \1005 ,
  \1006 ,
  \1007 ,
  \1008 ,
  \1009 ,
  \1010 ,
  \1011 ,
  \1012 ,
  \1013 ,
  \1014 ,
  \1015 ,
  \1016 ,
  \1017 ,
  \1018 ,
  \1019 ,
  \1020 ,
  \1021 ,
  \1022 ,
  \1023 ,
  \1024 ,
  \1025 ,
  \1026 ,
  \1027 ,
  \1028 ,
  \1029 ,
  \1030 ,
  \1031 ,
  \1032 ,
  \1033 ,
  \1034 ,
  \1035 ,
  \1036 ,
  \1037 ,
  \1038 ,
  \1039 ,
  \1040 ,
  \1041 ,
  \1042 ,
  \1043 ,
  \1044 ,
  \1045 ,
  \1046 ,
  \1047 ,
  \1048 ,
  \1049 ,
  \1050 ,
  \1051 ,
  \1052 ,
  \1053 ,
  \1054 ,
  \1055 ,
  \1056 ,
  \1057 ,
  \1058 ,
  \1059 ,
  \1060 ,
  \1061 ,
  \1062 ,
  \1063 ,
  \1064 ,
  \1065 ,
  \1066 ,
  \1067 ,
  \1068 ,
  \1069 ,
  \1070 ,
  \1071 ,
  \1072 ,
  \1073 ,
  \1074 ,
  \1075 ,
  \1076 ,
  \1077 ,
  \1078 ,
  \1079 ,
  \1080 ,
  \1081 ,
  \1082 ,
  \1083 ,
  \1084 ,
  \1085 ,
  \1086 ,
  \1087 ,
  \1088 ,
  \1089 ,
  \1090 ,
  \1091 ,
  \1092 ,
  \1093 ,
  \1094 ,
  \1095 ,
  \1096 ,
  \1097 ,
  \1098 ,
  \1099 ,
  \1100 ,
  \1101 ,
  \1102 ,
  \1103 ,
  \1104 ,
  \1105 ,
  \1106 ,
  \1107 ,
  \1108 ,
  \1109 ,
  \1110 ,
  \1111 ,
  \1112 ,
  \1113 ,
  \1114 ,
  \1115 ,
  \1116 ,
  \1117 ,
  \1118 ,
  \1119 ,
  \1120 ,
  \1121 ,
  \1122 ,
  \1123 ,
  \1124 ,
  \1125 ,
  \1126 ,
  \1127 ,
  \1128 ,
  \1129 ,
  \1130 ,
  \1131 ,
  \1132 ,
  \1133 ,
  \1134 ,
  \1135 ,
  \1136 ,
  \1137 ,
  \1138 ,
  \1139 ,
  \1140 ,
  \1141 ,
  \1142 ,
  \1143 ,
  \1144 ,
  \1145 ,
  \1146 ,
  \1147 ,
  \1148 ,
  \1149 ,
  \1150 ,
  \1151 ,
  \1152 ,
  \1153 ,
  \1154 ,
  \1155 ,
  \1156 ,
  \1157 ,
  \1158 ,
  \1159 ,
  \1160 ,
  \1161 ,
  \1162 ,
  \1163 ,
  \1164 ,
  \1165 ,
  \1166 ,
  \1167 ,
  \1168 ,
  \1169 ,
  \1170 ,
  \1171 ,
  \1172 ,
  \1173 ,
  \1174 ,
  \1175 ,
  \1176 ,
  \1177 ,
  \1178 ,
  \1179 ,
  \1180 ,
  \1181 ,
  \1182 ,
  \1183 ,
  \1184 ,
  \1185 ,
  \1186 ,
  \1187 ,
  \1188 ,
  \1189 ,
  \1190 ,
  \1191 ,
  \1192 ,
  \1193 ,
  \1194 ,
  \1195 ,
  \1196 ,
  \1197 ,
  \1198 ,
  \1199 ,
  \1200 ,
  \1201 ,
  \1202 ,
  \1203 ,
  \1204 ,
  \1205 ,
  \1206 ,
  \1207 ,
  \1208 ,
  \1209 ,
  \1210 ,
  \1211 ,
  \1212 ,
  \1213 ,
  \1214 ,
  \1215 ,
  \1216 ,
  \1217 ,
  \1218 ,
  \1219 ,
  \1220 ,
  \1221 ,
  \1222 ,
  \1223 ,
  \1224 ,
  \1225 ,
  \1226 ,
  \1227 ,
  \1228 ,
  \1229 ,
  \1230 ,
  \1231 ,
  \1232 ,
  \1233 ,
  \1234 ,
  \1235 ,
  \1236 ,
  \1237 ,
  \1238 ,
  \1239 ,
  \1240 ,
  \1241 ,
  \1242 ,
  \1243 ,
  \1244 ,
  \1245 ,
  \1246 ,
  \1247 ,
  \1248 ,
  \1249 ,
  \1250 ,
  \1251 ,
  \1252 ,
  \1253 ,
  \1254 ,
  \1255 ,
  \1256 ,
  \1257 ,
  \1258 ,
  \1259 ,
  \1260 ,
  \1261 ,
  \1262 ,
  \1263 ,
  \1264 ,
  \1265 ,
  \1266 ,
  \1267 ,
  \1268 ,
  \1269 ,
  \1270 ,
  \1271 ,
  \1272 ,
  \1273 ,
  \1274 ,
  \1275 ,
  \1276 ,
  \1277 ,
  \1278 ,
  \1279 ,
  \1280 ,
  \1281 ,
  \1282 ,
  \1283 ,
  \1284 ,
  \1285 ,
  \1286 ,
  \1287 ,
  \1288 ,
  \1289 ,
  \1290 ,
  \1291 ,
  \1292 ,
  \1293 ,
  \1294 ,
  \1295 ,
  \1296 ,
  \1297 ,
  \1298 ,
  \1299 ,
  \1300 ,
  \1301 ,
  \1302 ,
  \1303 ,
  \1304 ,
  \1305 ,
  \1306 ,
  \1307 ,
  \1308 ,
  \1309 ,
  \1310 ,
  \1311 ,
  \1312 ,
  \1313 ,
  \1314 ,
  \1315 ,
  \1316 ,
  \1317 ,
  \1318 ,
  \1319 ,
  \1320 ,
  \1321 ,
  \1322 ,
  \1323 ,
  \1324 ,
  \1325 ,
  \1326 ,
  \1327 ,
  \1328 ,
  \1329 ,
  \1330 ,
  \1331 ,
  \1332 ,
  \1333 ,
  \1334 ,
  \1335 ,
  \1336 ,
  \1337 ,
  \1338 ,
  \1339 ,
  \1340 ,
  \1341 ,
  \1342 ,
  \1343 ,
  \1344 ,
  \1345 ,
  \1346 ,
  \1347 ,
  \1348 ,
  \1349 ,
  \1350 ,
  \1351 ,
  \1352 ,
  \1353 ,
  \1354 ,
  \1355 ,
  \1356 ,
  \1357 ,
  \1358 ,
  \1359 ,
  \1360 ,
  \1361 ,
  \1362 ,
  \1363 ,
  \1364 ,
  \1365 ,
  \1366 ,
  \1367 ,
  \1368 ,
  \1369 ,
  \1370 ,
  \1371 ,
  \1372 ,
  \1373 ,
  \1374 ,
  \1375 ,
  \1376 ,
  \1377 ,
  \1378 ,
  \1379 ,
  \1380 ,
  \1381 ,
  \1382 ,
  \1383 ,
  \1384 ,
  \1385 ,
  \1386 ,
  \1387 ,
  \1388 ,
  \1389 ,
  \1390 ,
  \1391 ,
  \1392 ,
  \1393 ,
  \1394 ,
  \1395 ,
  \1396 ,
  \1397 ,
  \1398 ,
  \1399 ,
  \1400 ,
  \1401 ,
  \1402 ,
  \1403 ,
  \1404 ,
  \1405 ,
  \1406 ,
  \1407 ,
  \1408 ,
  \1409 ,
  \1410 ,
  \1411 ,
  \1412 ,
  \1413 ,
  \1414 ,
  \1415 ,
  \1416 ,
  \1417 ,
  \1418 ,
  \1419 ,
  \1420 ,
  \1421 ,
  \1422 ,
  \1423 ,
  \1424 ,
  \1425 ,
  \1426 ,
  \1427 ,
  \1428 ,
  \1429 ,
  \1430 ,
  \1431 ,
  \1432 ,
  \1433 ,
  \1434 ,
  \1435 ,
  \1436 ,
  \1437 ,
  \1438 ,
  \1439 ,
  \1440 ,
  \1441 ,
  \1442 ,
  \1443 ,
  \1444 ,
  \1445 ,
  \1446 ,
  \1447 ,
  \1448 ,
  \1449 ,
  \1450 ,
  \1451 ,
  \1452 ,
  \1453 ,
  \1454 ,
  \1455 ,
  \1456 ,
  \1457 ,
  \1458 ,
  \1459 ,
  \1460 ,
  \1461 ,
  \1462 ,
  \1463 ,
  \1464 ,
  \1465 ,
  \1466 ,
  \1467 ,
  \1468 ,
  \1469 ,
  \1470 ,
  \1471 ,
  \1472 ,
  \1473 ,
  \1474 ,
  \1475 ,
  \1476 ,
  \1477 ,
  \1478 ,
  \1479 ,
  \1480 ,
  \1481 ,
  \1482 ,
  \1483 ,
  \1484 ,
  \1485 ,
  \1486 ,
  \1487 ,
  \1488 ,
  \1489 ,
  \1490 ,
  \1491 ,
  \1492 ,
  \1493 ,
  \1494 ,
  \1495 ,
  \1496 ,
  \1497 ,
  \1498 ,
  \1499 ,
  \1500 ,
  \1501 ,
  \1502 ,
  \1503 ,
  \1504 ,
  \1505 ,
  \1506 ,
  \1507 ,
  \1508 ,
  \1509 ,
  \1510 ,
  \1511 ,
  \1512 ,
  \1513 ,
  \1514 ,
  \1515 ,
  \1516 ,
  \1517 ,
  \1518 ,
  \1519 ,
  \1520 ,
  \1521 ,
  \1522 ,
  \1523 ,
  \1524 ,
  \1525 ,
  \1526 ,
  \1527 ,
  \1528 ,
  \1529 ,
  \1530 ,
  \1531 ,
  \1532 ,
  \1533 ,
  \1534 ,
  \1535 ,
  \1536 ,
  \1537 ,
  \1538 ,
  \1539 ,
  \1540 ,
  \1541 ,
  \1542 ,
  \1543 ,
  \1544 ,
  \1545 ,
  \1546 ,
  \1547 ,
  \1548 ,
  \1549 ,
  \1550 ,
  \1551 ,
  \1552 ,
  \1553 ,
  \1554 ,
  \1555 ,
  \1556 ,
  \1557 ,
  \1558 ,
  \1559 ,
  \1560 ,
  \1561 ,
  \1562 ,
  \1563 ,
  \1564 ,
  \1565 ,
  \1566 ,
  \1567 ,
  \1568 ,
  \1569 ,
  \1570 ,
  \1571 ,
  \1572 ,
  \1573 ,
  \1574 ,
  \1575 ,
  \1576 ,
  \1577 ,
  \1578 ,
  \1579 ,
  \1580 ,
  \1581 ,
  \1582 ,
  \1583 ,
  \1584 ,
  \1585 ,
  \1586 ,
  \1587 ,
  \1588 ,
  \1589 ,
  \1590 ,
  \1591 ,
  \1592 ,
  \1593 ,
  \1594 ,
  \1595 ,
  \1596 ,
  \1597 ,
  \1598 ,
  \1599 ,
  \1600 ,
  \1601 ,
  \1602 ,
  \1603 ,
  \1604 ,
  \1605 ,
  \1606 ,
  \1607 ,
  \1608 ,
  \1609 ,
  \1610 ,
  \1611 ,
  \1612 ,
  \1613 ,
  \1614 ,
  \1615 ,
  \1616 ,
  \1617 ,
  \1618 ,
  \1619 ,
  \1620 ,
  \1621 ,
  \1622 ,
  \1623 ,
  \1624 ,
  \1625 ,
  \1626 ,
  \1627 ,
  \1628 ,
  \1629 ,
  \1630 ,
  \1631 ,
  \1632 ,
  \1633 ,
  \1634 ,
  \1635 ,
  \1636 ,
  \1637 ,
  \1638 ,
  \1639 ,
  \1640 ,
  \1641 ,
  \1642 ,
  \1643 ,
  \1644 ,
  \1645 ,
  \1646 ,
  \1647 ,
  \1648 ,
  \1649 ,
  \1650 ,
  \1651 ,
  \1652 ,
  \1653 ,
  \1654 ,
  \1655 ,
  \1656 ,
  \1657 ,
  \1658 ,
  \1659 ,
  \1660 ,
  \1661 ,
  \1662 ,
  \1663 ,
  \1664 ,
  \1665 ,
  \1666 ,
  \1667 ,
  \1668 ,
  \1669 ,
  \1670 ,
  \1671 ,
  \1672 ,
  \1673 ,
  \1674 ,
  \1675 ,
  \1676 ,
  \1677 ,
  \1678 ,
  \1679 ,
  \1680 ,
  \1681 ,
  \1682 ,
  \1683 ,
  \1684 ,
  \1685 ,
  \1686 ,
  \1687 ,
  \1688 ,
  \1689 ,
  \1690 ,
  \1691 ,
  \1692 ,
  \1693 ,
  \1694 ,
  \1695 ,
  \1696 ,
  \1697 ,
  \1698 ,
  \1699 ,
  \1700 ,
  \1701 ,
  \1702 ,
  \1703 ,
  \1704 ,
  \1705 ,
  \1706 ,
  \1707 ,
  \1708 ,
  \1709 ,
  \1710 ,
  \1711 ,
  \1712 ,
  \1713 ,
  \1714 ,
  \1715 ,
  \1716 ,
  \1717 ,
  \1718 ,
  \1719 ,
  \1720 ,
  \1721 ,
  \1722 ,
  \1723 ,
  \1724 ,
  \1725 ,
  \1726 ,
  \1727 ,
  \1728 ,
  \1729 ,
  \1730 ,
  \1731 ,
  \1732 ,
  \1733 ,
  \1734 ,
  \1735 ,
  \1736 ,
  \1737 ,
  \1738 ,
  \1739 ,
  \1740 ,
  \1741 ,
  \1742 ,
  \1743 ,
  \1744 ,
  \1745 ,
  \1746 ,
  \1747 ,
  \1748 ,
  \1749 ,
  \1750 ,
  \1751 ,
  \1752 ,
  \1753 ,
  \1754 ,
  \1755 ,
  \1756 ,
  \1757 ,
  \1758 ,
  \1759 ,
  \1760 ,
  \1761 ,
  \1762 ,
  \1763 ,
  \1764 ,
  \1765 ,
  \1766 ,
  \1767 ,
  \1768 ,
  \1769 ,
  \1770 ,
  \1771 ,
  \1772 ,
  \1773 ,
  \1774 ,
  \1775 ,
  \1776 ,
  \1777 ,
  \1778 ,
  \1779 ,
  \1780 ,
  \1781 ,
  \1782 ,
  \1783 ,
  \1784 ,
  \1785 ,
  \1786 ,
  \1787 ,
  \1788 ,
  \1789 ,
  \1790 ,
  \1791 ,
  \1792 ,
  \1793 ,
  \1794 ,
  \1795 ,
  \1796 ,
  \1797 ,
  \1798 ,
  \1799 ,
  \1800 ,
  \1801 ,
  \1802 ,
  \1803 ,
  \1804 ,
  \1805 ,
  \1806 ,
  \1807 ,
  \1808 ,
  \1809 ,
  \1810 ,
  \1811 ,
  \1812 ,
  \1813 ,
  \1814 ,
  \1815 ,
  \1816 ,
  \1817 ,
  \1818 ,
  \1819 ,
  \1820 ,
  \1821 ,
  \1822 ,
  \1823 ,
  \1824 ,
  \1825 ,
  \1826 ,
  \1827 ,
  \1828 ,
  \1829 ,
  \1830 ,
  \1831 ,
  \1832 ,
  \1833 ,
  \1834 ,
  \1835 ,
  \1836 ,
  \1837 ,
  \1838 ,
  \1839 ,
  \1840 ,
  \1841 ,
  \1842 ,
  \1843 ,
  \1844 ,
  \1845 ,
  \1846 ,
  \1847 ,
  \1848 ,
  \1849 ,
  \1850 ,
  \1851 ,
  \1852 ,
  \1853 ,
  \1854 ,
  \1855 ,
  \1856 ,
  \1857 ,
  \1858 ,
  \1859 ,
  \1860 ,
  \1861 ,
  \1862 ,
  \1863 ,
  \1864 ,
  \1865 ,
  \1866 ,
  \1867 ,
  \1868 ,
  \1869 ,
  \1870 ,
  \1871 ,
  \1872 ,
  \1873 ,
  \1874 ,
  \1875 ,
  \1876 ,
  \1877 ,
  \1878 ,
  \1879 ,
  \1880 ,
  \1881 ,
  \1882 ,
  \1883 ,
  \1884 ,
  \1885 ,
  \1886 ,
  \1887 ,
  \1888 ,
  \1889 ,
  \1890 ,
  \1891 ,
  \1892 ,
  \1893 ,
  \1894 ,
  \1895 ,
  \1896 ,
  \1897 ,
  \1898 ,
  \1899 ,
  \1900 ,
  \1901 ,
  \1902 ,
  \1903 ,
  \1904 ,
  \1905 ,
  \1906 ,
  \1907 ,
  \1908 ,
  \1909 ,
  \1910 ,
  \1911 ,
  \1912 ,
  \1913 ,
  \1914 ,
  \1915 ,
  \1916 ,
  \1917 ,
  \1918 ,
  \1919 ,
  \1920 ,
  \1921 ,
  \1922 ,
  \1923 ,
  \1924 ,
  \1925 ,
  \1926 ,
  \1927 ,
  \1928 ,
  \1929 ,
  \1930 ,
  \1931 ,
  \1932 ,
  \1933 ,
  \1934 ,
  \1935 ,
  \1936 ,
  \1937 ,
  \1938 ,
  \1939 ,
  \1940 ,
  \1941 ,
  \1942 ,
  \1943 ,
  \1944 ,
  \1945 ,
  \1946 ,
  \1947 ,
  \1948 ,
  \1949 ,
  \1950 ,
  \1951 ,
  \1952 ,
  \1953 ,
  \1954 ,
  \1955 ,
  \1956 ,
  \1957 ,
  \1958 ,
  \1959 ,
  \1960 ,
  \1961 ,
  \1962 ,
  \1963 ,
  \1964 ,
  \1965 ,
  \1966 ,
  \1967 ,
  \1968 ,
  \1969 ,
  \1970 ,
  \1971 ,
  \1972 ,
  \1973 ,
  \1974 ,
  \1975 ,
  \1976 ,
  \1977 ,
  \1978 ,
  \1979 ,
  \1980 ,
  \1981 ,
  \1982 ,
  \1983 ,
  \1984 ,
  \1985 ,
  \1986 ,
  \1987 ,
  \1988 ,
  \1989 ,
  \1990 ,
  \1991 ,
  \1992 ,
  \1993 ,
  \1994 ,
  \1995 ,
  \1996 ,
  \1997 ,
  \1998 ,
  \1999 ,
  \[100] ,
  \[101] ,
  \[102] ,
  \[103] ,
  \[104] ,
  \[105] ,
  \[106] ,
  \[107] ,
  \[108] ,
  \[109] ,
  \[110] ,
  \[111] ,
  \[112] ,
  \[113] ,
  \[114] ,
  \[115] ,
  \[116] ,
  \[117] ,
  \[118] ,
  \[119] ,
  \[120] ,
  \[121] ,
  \[122] ,
  \[123] ,
  \[124] ,
  \[125] ,
  \[126] ,
  \[127] ,
  \[128] ,
  \[129] ,
  \2000 ,
  \2001 ,
  \2002 ,
  \2003 ,
  \2004 ,
  \2005 ,
  \2006 ,
  \2007 ,
  \2008 ,
  \2009 ,
  \2010 ,
  \2011 ,
  \2012 ,
  \2013 ,
  \2014 ,
  \2015 ,
  \2016 ,
  \2017 ,
  \2018 ,
  \2019 ,
  \2020 ,
  \2021 ,
  \2022 ,
  \2023 ,
  \2024 ,
  \2025 ,
  \2026 ,
  \2027 ,
  \2028 ,
  \2029 ,
  \2030 ,
  \2031 ,
  \2032 ,
  \2033 ,
  \2034 ,
  \2035 ,
  \2036 ,
  \2037 ,
  \2038 ,
  \2039 ,
  \2040 ,
  \2041 ,
  \2042 ,
  \2043 ,
  \2044 ,
  \2045 ,
  \2046 ,
  \2047 ,
  \2048 ,
  \2049 ,
  \2050 ,
  \2051 ,
  \2052 ,
  \2053 ,
  \2054 ,
  \2055 ,
  \2056 ,
  \2057 ,
  \2058 ,
  \2059 ,
  \2060 ,
  \2061 ,
  \2062 ,
  \2063 ,
  \2064 ,
  \2065 ,
  \2066 ,
  \2067 ,
  \2068 ,
  \2069 ,
  \[130] ,
  \2070 ,
  \2071 ,
  \2072 ,
  \2073 ,
  \2074 ,
  \2075 ,
  \2076 ,
  \2077 ,
  \2078 ,
  \2079 ,
  \[131] ,
  \2080 ,
  \2081 ,
  \2082 ,
  \2083 ,
  \2084 ,
  \2085 ,
  \2086 ,
  \2087 ,
  \2088 ,
  \2089 ,
  \[132] ,
  \2090 ,
  \2091 ,
  \2092 ,
  \2093 ,
  \2094 ,
  \2095 ,
  \2096 ,
  \2097 ,
  \2098 ,
  \2099 ,
  \[133] ,
  \[134] ,
  \[135] ,
  \[136] ,
  \[137] ,
  \[138] ,
  \[139] ,
  \2100 ,
  \2101 ,
  \2102 ,
  \2103 ,
  \2104 ,
  \2105 ,
  \2106 ,
  \2107 ,
  \2108 ,
  \2109 ,
  \2110 ,
  \2111 ,
  \2112 ,
  \2113 ,
  \2114 ,
  \2115 ,
  \2116 ,
  \2117 ,
  \2118 ,
  \2119 ,
  \2120 ,
  \2121 ,
  \2122 ,
  \2123 ,
  \2124 ,
  \2125 ,
  \2126 ,
  \2127 ,
  \2128 ,
  \2129 ,
  \2130 ,
  \2131 ,
  \2132 ,
  \2133 ,
  \2134 ,
  \2135 ,
  \2136 ,
  \2137 ,
  \2138 ,
  \2139 ,
  \2140 ,
  \2141 ,
  \2142 ,
  \2143 ,
  \2144 ,
  \2145 ,
  \2146 ,
  \2147 ,
  \2148 ,
  \2149 ,
  \2150 ,
  \2151 ,
  \2152 ,
  \2153 ,
  \2154 ,
  \2155 ,
  \2156 ,
  \2157 ,
  \2158 ,
  \2159 ,
  \2160 ,
  \2161 ,
  \2162 ,
  \2163 ,
  \2164 ,
  \2165 ,
  \2166 ,
  \2167 ,
  \2168 ,
  \2169 ,
  \[140] ,
  \2170 ,
  \2171 ,
  \2172 ,
  \2173 ,
  \2174 ,
  \2175 ,
  \2176 ,
  \2177 ,
  \2178 ,
  \2179 ,
  \[141] ,
  \2180 ,
  \2181 ,
  \2182 ,
  \2183 ,
  \2184 ,
  \2185 ,
  \2186 ,
  \2187 ,
  \2188 ,
  \2189 ,
  \[142] ,
  \2190 ,
  \2191 ,
  \2192 ,
  \2193 ,
  \2194 ,
  \2195 ,
  \2196 ,
  \2197 ,
  \2198 ,
  \2199 ,
  \[143] ,
  \[144] ,
  \[145] ,
  \[146] ,
  \[147] ,
  \[148] ,
  \[149] ,
  \2200 ,
  \2201 ,
  \2202 ,
  \2203 ,
  \2204 ,
  \2205 ,
  \2206 ,
  \2207 ,
  \2208 ,
  \2209 ,
  \2210 ,
  \2211 ,
  \2212 ,
  \2213 ,
  \2214 ,
  \2215 ,
  \2216 ,
  \2217 ,
  \2218 ,
  \2219 ,
  \2220 ,
  \2221 ,
  \2222 ,
  \2223 ,
  \2224 ,
  \2225 ,
  \2226 ,
  \2227 ,
  \2228 ,
  \2229 ,
  \2230 ,
  \2231 ,
  \2232 ,
  \2233 ,
  \2234 ,
  \2235 ,
  \2236 ,
  \2237 ,
  \2238 ,
  \2239 ,
  \2240 ,
  \2241 ,
  \2242 ,
  \2243 ,
  \2244 ,
  \2245 ,
  \2246 ,
  \2247 ,
  \2248 ,
  \2249 ,
  \2250 ,
  \2251 ,
  \2252 ,
  \2253 ,
  \2254 ,
  \2255 ,
  \2256 ,
  \2257 ,
  \2258 ,
  \2259 ,
  \2260 ,
  \2261 ,
  \2262 ,
  \2263 ,
  \2264 ,
  \2265 ,
  \2266 ,
  \2267 ,
  \2268 ,
  \2269 ,
  \[150] ,
  \2270 ,
  \2271 ,
  \2272 ,
  \2273 ,
  \2274 ,
  \2275 ,
  \2276 ,
  \2277 ,
  \2278 ,
  \2279 ,
  \[151] ,
  \2280 ,
  \2281 ,
  \2282 ,
  \2283 ,
  \2284 ,
  \2285 ,
  \2286 ,
  \2287 ,
  \2288 ,
  \2289 ,
  \[152] ,
  \2290 ,
  \2291 ,
  \2292 ,
  \2293 ,
  \2294 ,
  \2295 ,
  \2296 ,
  \2297 ,
  \2298 ,
  \2299 ,
  \[153] ,
  \[154] ,
  \[155] ,
  \[156] ,
  \[157] ,
  \[158] ,
  \[159] ,
  \2300 ,
  \2301 ,
  \2302 ,
  \2303 ,
  \2304 ,
  \2305 ,
  \2306 ,
  \2307 ,
  \2308 ,
  \2309 ,
  \2310 ,
  \2311 ,
  \2312 ,
  \2313 ,
  \2314 ,
  \2315 ,
  \2316 ,
  \2317 ,
  \2318 ,
  \2319 ,
  \2320 ,
  \2321 ,
  \2322 ,
  \2323 ,
  \2324 ,
  \2325 ,
  \2326 ,
  \2327 ,
  \2328 ,
  \2329 ,
  \2330 ,
  \2331 ,
  \2332 ,
  \2333 ,
  \2334 ,
  \2335 ,
  \2336 ,
  \2337 ,
  \2338 ,
  \2339 ,
  \2340 ,
  \2341 ,
  \2342 ,
  \2343 ,
  \2344 ,
  \2345 ,
  \2346 ,
  \2347 ,
  \2348 ,
  \2349 ,
  \2350 ,
  \2351 ,
  \2352 ,
  \2353 ,
  \2354 ,
  \2355 ,
  \2356 ,
  \2357 ,
  \2358 ,
  \2359 ,
  \2360 ,
  \2361 ,
  \2362 ,
  \2363 ,
  \2364 ,
  \2365 ,
  \2366 ,
  \2367 ,
  \2368 ,
  \2369 ,
  \[160] ,
  \2370 ,
  \2371 ,
  \2372 ,
  \2373 ,
  \2374 ,
  \2375 ,
  \2376 ,
  \2377 ,
  \2378 ,
  \2379 ,
  \[161] ,
  \2380 ,
  \2381 ,
  \2382 ,
  \2383 ,
  \2384 ,
  \2385 ,
  \2386 ,
  \2387 ,
  \2388 ,
  \2389 ,
  \[162] ,
  \2390 ,
  \2391 ,
  \2392 ,
  \2393 ,
  \2394 ,
  \2395 ,
  \2396 ,
  \2397 ,
  \2398 ,
  \2399 ,
  \[163] ,
  \[164] ,
  \[165] ,
  \[166] ,
  \[167] ,
  \[168] ,
  \[169] ,
  \2400 ,
  \2401 ,
  \2402 ,
  \2403 ,
  \2404 ,
  \2405 ,
  \2406 ,
  \2407 ,
  \2408 ,
  \2409 ,
  \2410 ,
  \2411 ,
  \2412 ,
  \2413 ,
  \2414 ,
  \2415 ,
  \2416 ,
  \2417 ,
  \2418 ,
  \2419 ,
  \2420 ,
  \2421 ,
  \2422 ,
  \2423 ,
  \2424 ,
  \2425 ,
  \2426 ,
  \2427 ,
  \2428 ,
  \2429 ,
  \2430 ,
  \2431 ,
  \2432 ,
  \2433 ,
  \2434 ,
  \2435 ,
  \2436 ,
  \2437 ,
  \2438 ,
  \2439 ,
  \2440 ,
  \2441 ,
  \2442 ,
  \2443 ,
  \2444 ,
  \2445 ,
  \2446 ,
  \2447 ,
  \2448 ,
  \2449 ,
  \2450 ,
  \2451 ,
  \2452 ,
  \2453 ,
  \2454 ,
  \2455 ,
  \2456 ,
  \2457 ,
  \2458 ,
  \2459 ,
  \2460 ,
  \2461 ,
  \2462 ,
  \2463 ,
  \2464 ,
  \2465 ,
  \2466 ,
  \2467 ,
  \2468 ,
  \2469 ,
  \[170] ,
  \2470 ,
  \2471 ,
  \2472 ,
  \2473 ,
  \2474 ,
  \2475 ,
  \2476 ,
  \2477 ,
  \2478 ,
  \2479 ,
  \[171] ,
  \2480 ,
  \2481 ,
  \[172] ,
  \[173] ,
  \[174] ,
  \[175] ,
  \[176] ,
  \[177] ,
  \[178] ,
  \[179] ,
  \[180] ,
  \[181] ,
  \[182] ,
  \[183] ,
  \[184] ,
  \[185] ,
  \[186] ,
  \[187] ,
  \[188] ,
  \[189] ,
  \154 ,
  \155 ,
  \156 ,
  \157 ,
  \158 ,
  \159 ,
  \160 ,
  \161 ,
  \162 ,
  \163 ,
  \164 ,
  \165 ,
  \166 ,
  \167 ,
  \168 ,
  \169 ,
  \170 ,
  \171 ,
  \172 ,
  \173 ,
  \174 ,
  \175 ,
  \176 ,
  \177 ,
  \178 ,
  \179 ,
  \180 ,
  \181 ,
  \182 ,
  \183 ,
  \184 ,
  \185 ,
  \186 ,
  \187 ,
  \188 ,
  \189 ,
  \190 ,
  \191 ,
  \192 ,
  \193 ,
  \194 ,
  \195 ,
  \196 ,
  \[190] ,
  \197 ,
  \198 ,
  \199 ,
  \[191] ,
  \[192] ,
  \[193] ,
  \[194] ,
  \[195] ,
  \[196] ,
  \200 ,
  \201 ,
  \202 ,
  \203 ,
  \204 ,
  \205 ,
  \206 ,
  \[197] ,
  \207 ,
  \208 ,
  \209 ,
  \210 ,
  \211 ,
  \212 ,
  \213 ,
  \214 ,
  \215 ,
  \216 ,
  \[198] ,
  \217 ,
  \218 ,
  \219 ,
  \220 ,
  \221 ,
  \222 ,
  \223 ,
  \224 ,
  \225 ,
  \226 ,
  \[199] ,
  \227 ,
  \228 ,
  \229 ,
  \230 ,
  \231 ,
  \232 ,
  \233 ,
  \234 ,
  \235 ,
  \236 ,
  \237 ,
  \238 ,
  \239 ,
  \240 ,
  \241 ,
  \242 ,
  \243 ,
  \244 ,
  \245 ,
  \246 ,
  \247 ,
  \248 ,
  \249 ,
  \250 ,
  \251 ,
  \252 ,
  \253 ,
  \254 ,
  \255 ,
  \256 ,
  \257 ,
  \258 ,
  \259 ,
  \260 ,
  \261 ,
  \262 ,
  \263 ,
  \264 ,
  \265 ,
  \266 ,
  \267 ,
  \268 ,
  \269 ,
  \270 ,
  \271 ,
  \272 ,
  \273 ,
  \274 ,
  \275 ,
  \276 ,
  \277 ,
  \278 ,
  \279 ,
  \280 ,
  \281 ,
  \282 ,
  \283 ,
  \284 ,
  \285 ,
  \286 ,
  \287 ,
  \288 ,
  \289 ,
  \290 ,
  \291 ,
  \292 ,
  \293 ,
  \294 ,
  \295 ,
  \296 ,
  \297 ,
  \298 ,
  \299 ,
  \300 ,
  \301 ,
  \302 ,
  \303 ,
  \304 ,
  \305 ,
  \306 ,
  \307 ,
  \308 ,
  \309 ,
  \310 ,
  \311 ,
  \312 ,
  \313 ,
  \314 ,
  \315 ,
  \316 ,
  \317 ,
  \318 ,
  \319 ,
  \320 ,
  \321 ,
  \322 ,
  \323 ,
  \324 ,
  \325 ,
  \326 ,
  \327 ,
  \328 ,
  \329 ,
  \330 ,
  \331 ,
  \332 ,
  \333 ,
  \334 ,
  \335 ,
  \336 ,
  \337 ,
  \338 ,
  \339 ,
  \340 ,
  \341 ,
  \342 ,
  \343 ,
  \344 ,
  \345 ,
  \346 ,
  \347 ,
  \348 ,
  \349 ,
  \350 ,
  \351 ,
  \352 ,
  \353 ,
  \354 ,
  \355 ,
  \356 ,
  \357 ,
  \358 ,
  \359 ,
  \360 ,
  \361 ,
  \362 ,
  \363 ,
  \364 ,
  \365 ,
  \366 ,
  \367 ,
  \368 ,
  \369 ,
  \370 ,
  \371 ,
  \372 ,
  \373 ,
  \374 ,
  \375 ,
  \376 ,
  \377 ,
  \378 ,
  \379 ,
  \380 ,
  \381 ,
  \382 ,
  \383 ,
  \384 ,
  \385 ,
  \386 ,
  \387 ,
  \388 ,
  \389 ,
  \390 ,
  \391 ,
  \392 ,
  \393 ,
  \394 ,
  \395 ,
  \396 ,
  \397 ,
  \398 ,
  \399 ,
  \400 ,
  \401 ,
  \402 ,
  \403 ,
  \404 ,
  \405 ,
  \406 ,
  \407 ,
  \408 ,
  \409 ,
  \410 ,
  \411 ,
  \412 ,
  \413 ,
  \414 ,
  \415 ,
  \416 ,
  \417 ,
  \418 ,
  \419 ,
  \420 ,
  \421 ,
  \422 ,
  \423 ,
  \424 ,
  \425 ,
  \426 ,
  \427 ,
  \428 ,
  \429 ,
  \430 ,
  \431 ,
  \432 ,
  \433 ,
  \434 ,
  \435 ,
  \436 ,
  \437 ,
  \438 ,
  \439 ,
  \440 ,
  \441 ,
  \442 ,
  \443 ,
  \444 ,
  \445 ,
  \446 ,
  \447 ,
  \448 ,
  \449 ,
  \450 ,
  \451 ,
  \452 ,
  \453 ,
  \454 ,
  \455 ,
  \456 ,
  \457 ,
  \458 ,
  \459 ,
  \460 ,
  \461 ,
  \462 ,
  \463 ,
  \464 ,
  \465 ,
  \466 ,
  \467 ,
  \468 ,
  \469 ,
  \470 ,
  \471 ,
  \472 ,
  \473 ,
  \474 ,
  \475 ,
  \476 ,
  \477 ,
  \478 ,
  \479 ,
  \480 ,
  \481 ,
  \482 ,
  \483 ,
  \484 ,
  \485 ,
  \486 ,
  \487 ,
  \488 ,
  \489 ,
  \490 ,
  \491 ,
  \492 ,
  \493 ,
  \494 ,
  \495 ,
  \496 ,
  \497 ,
  \498 ,
  \499 ,
  \500 ,
  \501 ,
  \502 ,
  \503 ,
  \504 ,
  \505 ,
  \506 ,
  \507 ,
  \508 ,
  \509 ,
  \510 ,
  \511 ,
  \512 ,
  \513 ,
  \514 ,
  \515 ,
  \516 ,
  \517 ,
  \518 ,
  \519 ,
  \520 ,
  \521 ,
  \522 ,
  \523 ,
  \524 ,
  \525 ,
  \526 ,
  \527 ,
  \528 ,
  \529 ,
  \530 ,
  \531 ,
  \532 ,
  \533 ,
  \534 ,
  \535 ,
  \536 ,
  \537 ,
  \538 ,
  \539 ,
  \540 ,
  \541 ,
  \542 ,
  \543 ,
  \544 ,
  \545 ,
  \546 ,
  \547 ,
  \548 ,
  \549 ,
  \550 ,
  \551 ,
  \552 ,
  \553 ,
  \554 ,
  \555 ,
  \556 ,
  \557 ,
  \558 ,
  \559 ,
  \560 ,
  \561 ,
  \562 ,
  \563 ,
  \564 ,
  \565 ,
  \566 ,
  \567 ,
  \568 ,
  \569 ,
  \570 ,
  \571 ,
  \572 ,
  \573 ,
  \574 ,
  \575 ,
  \576 ,
  \577 ,
  \578 ,
  \579 ,
  \580 ,
  \581 ,
  \582 ,
  \583 ,
  \584 ,
  \585 ,
  \586 ,
  \587 ,
  \588 ,
  \589 ,
  \590 ,
  \591 ,
  \592 ,
  \593 ,
  \594 ,
  \595 ,
  \596 ,
  \597 ,
  \598 ,
  \599 ,
  \600 ,
  \601 ,
  \602 ,
  \603 ,
  \604 ,
  \605 ,
  \606 ,
  \607 ,
  \608 ,
  \609 ,
  \610 ,
  \611 ,
  \612 ,
  \613 ,
  \614 ,
  \615 ,
  \616 ,
  \617 ,
  \618 ,
  \619 ,
  \620 ,
  \621 ,
  \622 ,
  \623 ,
  \624 ,
  \625 ,
  \626 ,
  \627 ,
  \628 ,
  \629 ,
  \630 ,
  \631 ,
  \632 ,
  \633 ,
  \634 ,
  \635 ,
  \636 ,
  \637 ,
  \638 ,
  \639 ,
  \640 ,
  \641 ,
  \642 ,
  \643 ,
  \644 ,
  \645 ,
  \646 ,
  \647 ,
  \648 ,
  \649 ;
assign
  \650  = 0,
  \651  = 0,
  \652  = 0,
  \653  = 0,
  \654  = 0,
  \655  = 0,
  \656  = 0,
  \657  = 0,
  \658  = 0,
  \659  = 0,
  \660  = 0,
  \661  = 0,
  \662  = 0,
  \663  = 0,
  \664  = 0,
  \665  = 0,
  \666  = 0,
  \667  = 0,
  \668  = 0,
  \669  = 0,
  \670  = 0,
  \671  = 0,
  \672  = 0,
  \673  = 0,
  \674  = 1,
  \675  = 1,
  \676  = 1,
  \677  = 1,
  \678  = 1,
  \679  = 1,
  \680  = 1,
  \681  = 1,
  \682  = 1,
  \683  = 1,
  \684  = 1,
  \685  = 1,
  \686  = 1,
  \687  = 1,
  \688  = 1,
  \689  = 1,
  \690  = 1,
  \691  = 1,
  \692  = 1,
  \693  = 1,
  \694  = 1,
  \695  = 1,
  \696  = 1,
  \697  = 1,
  \698  = 1,
  \699  = 1,
  \700  = 1,
  \701  = 1,
  \702  = 1,
  \703  = 1,
  \704  = \33 ,
  \705  = 1,
  \706  = 1,
  \707  = 1,
  \708  = 1,
  \709  = 1,
  \710  = 1,
  \711  = 1,
  \712  = 1,
  \713  = 1,
  \714  = 1,
  \715  = 1,
  \716  = 1,
  \717  = 1,
  \718  = 1,
  \719  = 1,
  \720  = 1,
  \721  = 1,
  \722  = 1,
  \723  = 1,
  \724  = 1,
  \725  = 1,
  \726  = 1,
  \727  = 1,
  \728  = 1,
  \729  = 1,
  \730  = 1,
  \731  = 1,
  \732  = 1,
  \733  = 1,
  \734  = 1,
  \735  = \32 ,
  \736  = \31 ,
  \737  = \30 ,
  \738  = \29 ,
  \739  = \28 ,
  \740  = \27 ,
  \741  = \26 ,
  \742  = \25 ,
  \743  = \24 ,
  \744  = \23 ,
  \745  = \22 ,
  \746  = \21 ,
  \747  = \20 ,
  \748  = \19 ,
  \749  = \18 ,
  \750  = \17 ,
  \751  = \16 ,
  \752  = \15 ,
  \753  = \14 ,
  \754  = \13 ,
  \755  = \12 ,
  \756  = \11 ,
  \757  = \10 ,
  \758  = \9 ,
  \759  = \8 ,
  \760  = \7 ,
  \761  = \6 ,
  \762  = \5 ,
  \763  = 0,
  \764  = \4 ,
  \765  = \94 ,
  \766  = \95 ,
  \767  = \96 ,
  \768  = \97 ,
  \769  = \98 ,
  \770  = \99 ,
  \771  = \100 ,
  \772  = \101 ,
  \773  = \102 ,
  \774  = \103 ,
  \775  = \104 ,
  \776  = \105 ,
  \777  = \106 ,
  \778  = \107 ,
  \779  = \108 ,
  \780  = \109 ,
  \781  = \110 ,
  \782  = \111 ,
  \783  = \112 ,
  \784  = \113 ,
  \785  = \114 ,
  \786  = \115 ,
  \787  = \116 ,
  \788  = \117 ,
  \789  = \118 ,
  \790  = \119 ,
  \791  = \120 ,
  \792  = \121 ,
  \793  = \122 ,
  \794  = \123 ,
  \795  = \4 ,
  \796  = \5 ,
  \797  = \6 ,
  \798  = \7 ,
  \799  = \8 ,
  \800  = \9 ,
  \801  = \10 ,
  \802  = \11 ,
  \803  = \12 ,
  \804  = \13 ,
  \805  = \14 ,
  \806  = \15 ,
  \807  = \16 ,
  \808  = \17 ,
  \809  = \18 ,
  \810  = \19 ,
  \811  = \20 ,
  \812  = \21 ,
  \813  = \22 ,
  \814  = \23 ,
  \815  = \24 ,
  \816  = \25 ,
  \817  = \26 ,
  \818  = \27 ,
  \819  = \28 ,
  \820  = \29 ,
  \821  = \30 ,
  \822  = \31 ,
  \823  = \32 ,
  \824  = \33 ,
  \825  = \33 ,
  \826  = \32 ,
  \827  = \31 ,
  \828  = \30 ,
  \829  = \29 ,
  \830  = \28 ,
  \831  = \27 ,
  \832  = \26 ,
  \833  = \25 ,
  \834  = \24 ,
  \835  = \23 ,
  \836  = \22 ,
  \837  = \21 ,
  \838  = \20 ,
  \839  = \19 ,
  \840  = \18 ,
  \841  = \17 ,
  \842  = \16 ,
  \843  = \15 ,
  \844  = \14 ,
  \845  = \13 ,
  \846  = \12 ,
  \847  = \11 ,
  \848  = \10 ,
  \849  = \9 ,
  \850  = \8 ,
  \851  = \7 ,
  \852  = \6 ,
  \853  = \5 ,
  \854  = 0,
  \855  = \4 ,
  \856  = \64 ,
  \857  = \65 ,
  \858  = \66 ,
  \859  = \67 ,
  \860  = \68 ,
  \861  = \69 ,
  \862  = \70 ,
  \863  = \71 ,
  \864  = \72 ,
  \865  = \73 ,
  \866  = \74 ,
  \867  = \75 ,
  \868  = \76 ,
  \869  = \77 ,
  \870  = \78 ,
  \871  = \79 ,
  \872  = \80 ,
  \873  = \81 ,
  \874  = \82 ,
  \875  = \83 ,
  \876  = \84 ,
  \877  = \85 ,
  \878  = \86 ,
  \879  = \87 ,
  \880  = \88 ,
  \881  = \89 ,
  \882  = \90 ,
  \883  = \91 ,
  \884  = \92 ,
  \885  = \93 ,
  \886  = \4 ,
  \887  = \5 ,
  \888  = \6 ,
  \889  = \7 ,
  \890  = \8 ,
  \891  = \9 ,
  \892  = \10 ,
  \893  = \11 ,
  \894  = \12 ,
  \895  = \13 ,
  \896  = \14 ,
  \[200]  = \234 ,
  \897  = \15 ,
  \898  = \16 ,
  \899  = \17 ,
  \[201]  = \235 ,
  \[202]  = \236 ,
  \[203]  = \237 ,
  \[204]  = \238 ,
  \[205]  = \239 ,
  \[206]  = \240 ,
  \900  = \18 ,
  \901  = \19 ,
  \902  = \20 ,
  \903  = \21 ,
  \904  = \22 ,
  \905  = \23 ,
  \906  = \24 ,
  \[207]  = \241 ,
  \907  = \25 ,
  \908  = \26 ,
  \909  = \27 ,
  \910  = \28 ,
  \911  = \29 ,
  \912  = \30 ,
  \913  = \31 ,
  \914  = \32 ,
  \915  = \33 ,
  \916  = (\1127  & \1126 ) | ((\1127  & \1125 ) | (\1126  & \1125 )),
  \[208]  = \242 ,
  \917  = (~\1043  & (~\1042  & \1041 )) | ((~\1043  & (\1042  & ~\1041 )) | ((\1043  & (~\1042  & ~\1041 )) | (\1043  & (\1042  & \1041 )))),
  \918  = (~\1046  & (~\1045  & \1044 )) | ((~\1046  & (\1045  & ~\1044 )) | ((\1046  & (~\1045  & ~\1044 )) | (\1046  & (\1045  & \1044 )))),
  \919  = (~\1049  & (~\1048  & \1047 )) | ((~\1049  & (\1048  & ~\1047 )) | ((\1049  & (~\1048  & ~\1047 )) | (\1049  & (\1048  & \1047 )))),
  \920  = (~\1052  & (~\1051  & \1050 )) | ((~\1052  & (\1051  & ~\1050 )) | ((\1052  & (~\1051  & ~\1050 )) | (\1052  & (\1051  & \1050 )))),
  \921  = (~\1055  & (~\1054  & \1053 )) | ((~\1055  & (\1054  & ~\1053 )) | ((\1055  & (~\1054  & ~\1053 )) | (\1055  & (\1054  & \1053 )))),
  \922  = (~\1058  & (~\1057  & \1056 )) | ((~\1058  & (\1057  & ~\1056 )) | ((\1058  & (~\1057  & ~\1056 )) | (\1058  & (\1057  & \1056 )))),
  \923  = (~\1061  & (~\1060  & \1059 )) | ((~\1061  & (\1060  & ~\1059 )) | ((\1061  & (~\1060  & ~\1059 )) | (\1061  & (\1060  & \1059 )))),
  \924  = (~\1064  & (~\1063  & \1062 )) | ((~\1064  & (\1063  & ~\1062 )) | ((\1064  & (~\1063  & ~\1062 )) | (\1064  & (\1063  & \1062 )))),
  \925  = (~\1067  & (~\1066  & \1065 )) | ((~\1067  & (\1066  & ~\1065 )) | ((\1067  & (~\1066  & ~\1065 )) | (\1067  & (\1066  & \1065 )))),
  \926  = (~\1070  & (~\1069  & \1068 )) | ((~\1070  & (\1069  & ~\1068 )) | ((\1070  & (~\1069  & ~\1068 )) | (\1070  & (\1069  & \1068 )))),
  \[209]  = \243 ,
  \927  = (~\1073  & (~\1072  & \1071 )) | ((~\1073  & (\1072  & ~\1071 )) | ((\1073  & (~\1072  & ~\1071 )) | (\1073  & (\1072  & \1071 )))),
  \928  = (~\1076  & (~\1075  & \1074 )) | ((~\1076  & (\1075  & ~\1074 )) | ((\1076  & (~\1075  & ~\1074 )) | (\1076  & (\1075  & \1074 )))),
  \929  = (~\1079  & (~\1078  & \1077 )) | ((~\1079  & (\1078  & ~\1077 )) | ((\1079  & (~\1078  & ~\1077 )) | (\1079  & (\1078  & \1077 )))),
  \930  = (~\1082  & (~\1081  & \1080 )) | ((~\1082  & (\1081  & ~\1080 )) | ((\1082  & (~\1081  & ~\1080 )) | (\1082  & (\1081  & \1080 )))),
  \931  = (~\1085  & (~\1084  & \1083 )) | ((~\1085  & (\1084  & ~\1083 )) | ((\1085  & (~\1084  & ~\1083 )) | (\1085  & (\1084  & \1083 )))),
  \932  = (~\1088  & (~\1087  & \1086 )) | ((~\1088  & (\1087  & ~\1086 )) | ((\1088  & (~\1087  & ~\1086 )) | (\1088  & (\1087  & \1086 )))),
  \933  = (~\1091  & (~\1090  & \1089 )) | ((~\1091  & (\1090  & ~\1089 )) | ((\1091  & (~\1090  & ~\1089 )) | (\1091  & (\1090  & \1089 )))),
  \934  = (~\1094  & (~\1093  & \1092 )) | ((~\1094  & (\1093  & ~\1092 )) | ((\1094  & (~\1093  & ~\1092 )) | (\1094  & (\1093  & \1092 )))),
  \935  = (~\1097  & (~\1096  & \1095 )) | ((~\1097  & (\1096  & ~\1095 )) | ((\1097  & (~\1096  & ~\1095 )) | (\1097  & (\1096  & \1095 )))),
  \936  = (~\1100  & (~\1099  & \1098 )) | ((~\1100  & (\1099  & ~\1098 )) | ((\1100  & (~\1099  & ~\1098 )) | (\1100  & (\1099  & \1098 )))),
  \937  = (~\1103  & (~\1102  & \1101 )) | ((~\1103  & (\1102  & ~\1101 )) | ((\1103  & (~\1102  & ~\1101 )) | (\1103  & (\1102  & \1101 )))),
  \938  = (~\1106  & (~\1105  & \1104 )) | ((~\1106  & (\1105  & ~\1104 )) | ((\1106  & (~\1105  & ~\1104 )) | (\1106  & (\1105  & \1104 )))),
  \939  = (~\1109  & (~\1108  & \1107 )) | ((~\1109  & (\1108  & ~\1107 )) | ((\1109  & (~\1108  & ~\1107 )) | (\1109  & (\1108  & \1107 )))),
  \940  = (~\1112  & (~\1111  & \1110 )) | ((~\1112  & (\1111  & ~\1110 )) | ((\1112  & (~\1111  & ~\1110 )) | (\1112  & (\1111  & \1110 )))),
  \941  = (~\1115  & (~\1114  & \1113 )) | ((~\1115  & (\1114  & ~\1113 )) | ((\1115  & (~\1114  & ~\1113 )) | (\1115  & (\1114  & \1113 )))),
  \942  = (~\1118  & (~\1117  & \1116 )) | ((~\1118  & (\1117  & ~\1116 )) | ((\1118  & (~\1117  & ~\1116 )) | (\1118  & (\1117  & \1116 )))),
  \943  = (~\1121  & (~\1120  & \1119 )) | ((~\1121  & (\1120  & ~\1119 )) | ((\1121  & (~\1120  & ~\1119 )) | (\1121  & (\1120  & \1119 )))),
  \944  = (~\1124  & (~\1123  & \1122 )) | ((~\1124  & (\1123  & ~\1122 )) | ((\1124  & (~\1123  & ~\1122 )) | (\1124  & (\1123  & \1122 )))),
  \945  = (~\1127  & (~\1126  & \1125 )) | ((~\1127  & (\1126  & ~\1125 )) | ((\1127  & (~\1126  & ~\1125 )) | (\1127  & (\1126  & \1125 )))),
  \946  = \916 ,
  \947  = \917 ,
  \948  = \918 ,
  \949  = \919 ,
  \950  = \920 ,
  \951  = \921 ,
  \952  = \922 ,
  \953  = \923 ,
  \954  = \924 ,
  \955  = \925 ,
  \956  = \926 ,
  \957  = \927 ,
  \958  = \928 ,
  \959  = \929 ,
  \960  = \930 ,
  \961  = \931 ,
  \962  = \932 ,
  \963  = \933 ,
  \964  = \934 ,
  \965  = \935 ,
  \966  = \936 ,
  \967  = \937 ,
  \968  = \938 ,
  \969  = \939 ,
  \970  = \940 ,
  \971  = \941 ,
  \972  = \942 ,
  \973  = \943 ,
  \974  = \944 ,
  \975  = \945 ,
  \976  = \1039 ,
  \977  = \1042 ,
  \978  = \1045 ,
  \979  = \1048 ,
  \980  = \1051 ,
  \981  = \1054 ,
  \982  = \1057 ,
  \983  = \1060 ,
  \984  = \1063 ,
  \985  = \1066 ,
  \986  = \1069 ,
  \987  = \1072 ,
  \988  = \1075 ,
  \989  = \1078 ,
  \990  = \1081 ,
  \991  = \1084 ,
  \992  = \1087 ,
  \993  = \1090 ,
  \994  = \1093 ,
  \995  = \1096 ,
  \996  = \1099 ,
  \997  = \1102 ,
  \998  = \1105 ,
  \999  = \1108 ,
  \[90]  = \1135  | \1134 ,
  \[91]  = \1143  | \1142 ,
  \[92]  = \1151  | \1150 ,
  \[93]  = \1159  | \1158 ,
  \[94]  = \1167  | \1166 ,
  \[95]  = \1175  | \1174 ,
  \[96]  = \1183  | \1182 ,
  \[97]  = \1191  | \1190 ,
  \[98]  = \1199  | \1198 ,
  \[99]  = \1207  | \1206 ,
  \1000  = \1111 ,
  \1001  = \1114 ,
  \1002  = \1117 ,
  \1003  = \1120 ,
  \1004  = \1123 ,
  \1005  = \1126 ,
  \1006  = \1040 ,
  \1007  = \1043 ,
  \1008  = \1046 ,
  \1009  = \1049 ,
  \1010  = \1052 ,
  \1011  = \1055 ,
  \1012  = \1058 ,
  \1013  = \1061 ,
  \1014  = \1064 ,
  \1015  = \1067 ,
  \1016  = \1070 ,
  \1017  = \1073 ,
  \1018  = \1076 ,
  \1019  = \1079 ,
  \1020  = \1082 ,
  \1021  = \1085 ,
  \1022  = \1088 ,
  \1023  = \1091 ,
  \1024  = \1094 ,
  \1025  = \1097 ,
  \1026  = \1100 ,
  \1027  = \1103 ,
  \1028  = \1106 ,
  \1029  = \1109 ,
  \1030  = \1112 ,
  \1031  = \1115 ,
  \1032  = \1118 ,
  \1033  = \1121 ,
  \1034  = \1124 ,
  \1035  = \1127 ,
  \1036  = \2481  & \2479 ,
  \1037  = \2389  & \2387 ,
  \1038  = 0,
  \1039  = \2297  & \2295 ,
  \1040  = \2292  & \2290 ,
  \1041  = (\1040  & \1039 ) | ((\1040  & \1038 ) | (\1039  & \1038 )),
  \1042  = \2287  & \2285 ,
  \1043  = \2282  & \2280 ,
  \1044  = (\1043  & \1042 ) | ((\1043  & \1041 ) | (\1042  & \1041 )),
  \1045  = \2277  & \2275 ,
  \1046  = \2272  & \2270 ,
  \1047  = (\1046  & \1045 ) | ((\1046  & \1044 ) | (\1045  & \1044 )),
  \1048  = \2267  & \2265 ,
  \1049  = \2262  & \2260 ,
  \1050  = (\1049  & \1048 ) | ((\1049  & \1047 ) | (\1048  & \1047 )),
  \1051  = \2257  & \2255 ,
  \1052  = \2252  & \2250 ,
  \1053  = (\1052  & \1051 ) | ((\1052  & \1050 ) | (\1051  & \1050 )),
  \1054  = \2247  & \2245 ,
  \1055  = \2242  & \2240 ,
  \1056  = (\1055  & \1054 ) | ((\1055  & \1053 ) | (\1054  & \1053 )),
  \1057  = \2237  & \2235 ,
  \1058  = \2232  & \2230 ,
  \1059  = (\1058  & \1057 ) | ((\1058  & \1056 ) | (\1057  & \1056 )),
  \1060  = \2227  & \2225 ,
  \1061  = \2222  & \2220 ,
  \1062  = (\1061  & \1060 ) | ((\1061  & \1059 ) | (\1060  & \1059 )),
  \1063  = \2217  & \2215 ,
  \1064  = \2212  & \2210 ,
  \1065  = (\1064  & \1063 ) | ((\1064  & \1062 ) | (\1063  & \1062 )),
  \1066  = \2207  & \2205 ,
  \1067  = \2202  & \2200 ,
  \1068  = (\1067  & \1066 ) | ((\1067  & \1065 ) | (\1066  & \1065 )),
  \1069  = \2197  & \2195 ,
  \1070  = \2192  & \2190 ,
  \1071  = (\1070  & \1069 ) | ((\1070  & \1068 ) | (\1069  & \1068 )),
  \1072  = \2187  & \2185 ,
  \1073  = \2182  & \2180 ,
  \1074  = (\1073  & \1072 ) | ((\1073  & \1071 ) | (\1072  & \1071 )),
  \1075  = \2177  & \2175 ,
  \1076  = \2172  & \2170 ,
  \1077  = (\1076  & \1075 ) | ((\1076  & \1074 ) | (\1075  & \1074 )),
  \1078  = \2167  & \2165 ,
  \1079  = \2162  & \2160 ,
  \1080  = (\1079  & \1078 ) | ((\1079  & \1077 ) | (\1078  & \1077 )),
  \1081  = \2157  & \2155 ,
  \1082  = \2152  & \2150 ,
  \1083  = (\1082  & \1081 ) | ((\1082  & \1080 ) | (\1081  & \1080 )),
  \1084  = \2147  & \2145 ,
  \1085  = \2142  & \2140 ,
  \1086  = (\1085  & \1084 ) | ((\1085  & \1083 ) | (\1084  & \1083 )),
  \1087  = \2137  & \2135 ,
  \1088  = \2132  & \2130 ,
  \1089  = (\1088  & \1087 ) | ((\1088  & \1086 ) | (\1087  & \1086 )),
  \1090  = \2127  & \2125 ,
  \1091  = \2122  & \2120 ,
  \1092  = (\1091  & \1090 ) | ((\1091  & \1089 ) | (\1090  & \1089 )),
  \1093  = \2117  & \2115 ,
  \1094  = \2112  & \2110 ,
  \1095  = (\1094  & \1093 ) | ((\1094  & \1092 ) | (\1093  & \1092 )),
  \1096  = \2107  & \2105 ,
  \1097  = \2102  & \2100 ,
  \1098  = (\1097  & \1096 ) | ((\1097  & \1095 ) | (\1096  & \1095 )),
  \1099  = \2097  & \2095 ,
  \1100  = \2092  & \2090 ,
  \1101  = (\1100  & \1099 ) | ((\1100  & \1098 ) | (\1099  & \1098 )),
  \1102  = \2087  & \2085 ,
  \1103  = \2082  & \2080 ,
  \1104  = (\1103  & \1102 ) | ((\1103  & \1101 ) | (\1102  & \1101 )),
  \1105  = \2077  & \2075 ,
  \1106  = \2072  & \2070 ,
  \1107  = (\1106  & \1105 ) | ((\1106  & \1104 ) | (\1105  & \1104 )),
  \1108  = \2067  & \2065 ,
  \1109  = \2062  & \2060 ,
  \1110  = (\1109  & \1108 ) | ((\1109  & \1107 ) | (\1108  & \1107 )),
  \1111  = \2057  & \2055 ,
  \1112  = \2052  & \2050 ,
  \1113  = (\1112  & \1111 ) | ((\1112  & \1110 ) | (\1111  & \1110 )),
  \1114  = \2047  & \2045 ,
  \1115  = \2042  & \2040 ,
  \1116  = (\1115  & \1114 ) | ((\1115  & \1113 ) | (\1114  & \1113 )),
  \1117  = \2037  & \2035 ,
  \1118  = \2032  & \2030 ,
  \1119  = (\1118  & \1117 ) | ((\1118  & \1116 ) | (\1117  & \1116 )),
  \1120  = \2027  & \2025 ,
  \1121  = \2022  & \2020 ,
  \1122  = (\1121  & \1120 ) | ((\1121  & \1119 ) | (\1120  & \1119 )),
  \1123  = \2017  & \2015 ,
  \1124  = \2012  & \2010 ,
  \1125  = (\1124  & \1123 ) | ((\1124  & \1122 ) | (\1123  & \1122 )),
  \1126  = \2007  & \2005 ,
  \1127  = \2002  & \2000 ,
  \1128  = \947  & \248 ,
  \1129  = \584  & \249 ,
  \1130  = \1129  | \1128 ,
  \1131  = \1130  & \246 ,
  \1132  = \464  & \247 ,
  \1133  = \1132  | \1131 ,
  \1134  = \1133  & \244 ,
  \1135  = \374  & \245 ,
  \1136  = \948  & \248 ,
  \1137  = \585  & \249 ,
  \1138  = \1137  | \1136 ,
  \1139  = \1138  & \246 ,
  \1140  = \465  & \247 ,
  \1141  = \1140  | \1139 ,
  \1142  = \1141  & \244 ,
  \1143  = \375  & \245 ,
  \1144  = \949  & \248 ,
  \1145  = \586  & \249 ,
  \1146  = \1145  | \1144 ,
  \1147  = \1146  & \246 ,
  \1148  = \466  & \247 ,
  \1149  = \1148  | \1147 ,
  \1150  = \1149  & \244 ,
  \1151  = \376  & \245 ,
  \1152  = \950  & \248 ,
  \1153  = \587  & \249 ,
  \1154  = \1153  | \1152 ,
  \1155  = \1154  & \246 ,
  \1156  = \467  & \247 ,
  \1157  = \1156  | \1155 ,
  \1158  = \1157  & \244 ,
  \1159  = \377  & \245 ,
  \1160  = \951  & \248 ,
  \1161  = \588  & \249 ,
  \1162  = \1161  | \1160 ,
  \1163  = \1162  & \246 ,
  \1164  = \468  & \247 ,
  \1165  = \1164  | \1163 ,
  \1166  = \1165  & \244 ,
  \1167  = \378  & \245 ,
  \1168  = \952  & \248 ,
  \1169  = \589  & \249 ,
  \1170  = \1169  | \1168 ,
  \1171  = \1170  & \246 ,
  \1172  = \469  & \247 ,
  \1173  = \1172  | \1171 ,
  \1174  = \1173  & \244 ,
  \1175  = \379  & \245 ,
  \1176  = \953  & \248 ,
  \1177  = \590  & \249 ,
  \1178  = \1177  | \1176 ,
  \1179  = \1178  & \246 ,
  \1180  = \470  & \247 ,
  \1181  = \1180  | \1179 ,
  \1182  = \1181  & \244 ,
  \1183  = \380  & \245 ,
  \1184  = \954  & \248 ,
  \1185  = \591  & \249 ,
  \1186  = \1185  | \1184 ,
  \1187  = \1186  & \246 ,
  \1188  = \471  & \247 ,
  \1189  = \1188  | \1187 ,
  \1190  = \1189  & \244 ,
  \1191  = \381  & \245 ,
  \1192  = \955  & \248 ,
  \1193  = \592  & \249 ,
  \1194  = \1193  | \1192 ,
  \1195  = \1194  & \246 ,
  \1196  = \472  & \247 ,
  \1197  = \1196  | \1195 ,
  \1198  = \1197  & \244 ,
  \1199  = \382  & \245 ,
  \1200  = \956  & \248 ,
  \1201  = \593  & \249 ,
  \1202  = \1201  | \1200 ,
  \1203  = \1202  & \246 ,
  \1204  = \473  & \247 ,
  \1205  = \1204  | \1203 ,
  \1206  = \1205  & \244 ,
  \1207  = \383  & \245 ,
  \1208  = \957  & \248 ,
  \1209  = \594  & \249 ,
  \1210  = \1209  | \1208 ,
  \1211  = \1210  & \246 ,
  \1212  = \474  & \247 ,
  \1213  = \1212  | \1211 ,
  \1214  = \1213  & \244 ,
  \1215  = \384  & \245 ,
  \1216  = \958  & \248 ,
  \1217  = \595  & \249 ,
  \1218  = \1217  | \1216 ,
  \1219  = \1218  & \246 ,
  \1220  = \475  & \247 ,
  \1221  = \1220  | \1219 ,
  \1222  = \1221  & \244 ,
  \1223  = \385  & \245 ,
  \1224  = \959  & \248 ,
  \1225  = \596  & \249 ,
  \1226  = \1225  | \1224 ,
  \1227  = \1226  & \246 ,
  \1228  = \476  & \247 ,
  \1229  = \1228  | \1227 ,
  \1230  = \1229  & \244 ,
  \1231  = \386  & \245 ,
  \1232  = \960  & \248 ,
  \1233  = \597  & \249 ,
  \1234  = \1233  | \1232 ,
  \1235  = \1234  & \246 ,
  \1236  = \477  & \247 ,
  \1237  = \1236  | \1235 ,
  \1238  = \1237  & \244 ,
  \1239  = \387  & \245 ,
  \1240  = \961  & \248 ,
  \1241  = \598  & \249 ,
  \1242  = \1241  | \1240 ,
  \1243  = \1242  & \246 ,
  \1244  = \478  & \247 ,
  \1245  = \1244  | \1243 ,
  \1246  = \1245  & \244 ,
  \1247  = \388  & \245 ,
  \1248  = \962  & \248 ,
  \1249  = \599  & \249 ,
  \1250  = \1249  | \1248 ,
  \1251  = \1250  & \246 ,
  \1252  = \479  & \247 ,
  \1253  = \1252  | \1251 ,
  \1254  = \1253  & \244 ,
  \1255  = \389  & \245 ,
  \1256  = \963  & \248 ,
  \1257  = \600  & \249 ,
  \1258  = \1257  | \1256 ,
  \1259  = \1258  & \246 ,
  \1260  = \480  & \247 ,
  \1261  = \1260  | \1259 ,
  \1262  = \1261  & \244 ,
  \1263  = \390  & \245 ,
  \1264  = \964  & \248 ,
  \1265  = \601  & \249 ,
  \1266  = \1265  | \1264 ,
  \1267  = \1266  & \246 ,
  \1268  = \481  & \247 ,
  \1269  = \1268  | \1267 ,
  \1270  = \1269  & \244 ,
  \1271  = \391  & \245 ,
  \1272  = \965  & \248 ,
  \1273  = \602  & \249 ,
  \1274  = \1273  | \1272 ,
  \1275  = \1274  & \246 ,
  \1276  = \482  & \247 ,
  \1277  = \1276  | \1275 ,
  \1278  = \1277  & \244 ,
  \1279  = \392  & \245 ,
  \1280  = \966  & \248 ,
  \1281  = \603  & \249 ,
  \1282  = \1281  | \1280 ,
  \1283  = \1282  & \246 ,
  \1284  = \483  & \247 ,
  \1285  = \1284  | \1283 ,
  \1286  = \1285  & \244 ,
  \1287  = \393  & \245 ,
  \1288  = \967  & \248 ,
  \1289  = \604  & \249 ,
  \1290  = \1289  | \1288 ,
  \1291  = \1290  & \246 ,
  \1292  = \484  & \247 ,
  \1293  = \1292  | \1291 ,
  \1294  = \1293  & \244 ,
  \1295  = \394  & \245 ,
  \1296  = \968  & \248 ,
  \1297  = \605  & \249 ,
  \1298  = \1297  | \1296 ,
  \1299  = \1298  & \246 ,
  \1300  = \485  & \247 ,
  \1301  = \1300  | \1299 ,
  \1302  = \1301  & \244 ,
  \1303  = \395  & \245 ,
  \1304  = \969  & \248 ,
  \1305  = \606  & \249 ,
  \1306  = \1305  | \1304 ,
  \1307  = \1306  & \246 ,
  \1308  = \486  & \247 ,
  \1309  = \1308  | \1307 ,
  \1310  = \1309  & \244 ,
  \1311  = \396  & \245 ,
  \1312  = \970  & \248 ,
  \1313  = \607  & \249 ,
  \1314  = \1313  | \1312 ,
  \1315  = \1314  & \246 ,
  \1316  = \487  & \247 ,
  \1317  = \1316  | \1315 ,
  \1318  = \1317  & \244 ,
  \1319  = \397  & \245 ,
  \1320  = \971  & \248 ,
  \1321  = \608  & \249 ,
  \1322  = \1321  | \1320 ,
  \1323  = \1322  & \246 ,
  \1324  = \488  & \247 ,
  \1325  = \1324  | \1323 ,
  \1326  = \1325  & \244 ,
  \1327  = \398  & \245 ,
  \1328  = \972  & \248 ,
  \1329  = \609  & \249 ,
  \1330  = \1329  | \1328 ,
  \1331  = \1330  & \246 ,
  \1332  = \489  & \247 ,
  \1333  = \1332  | \1331 ,
  \1334  = \1333  & \244 ,
  \1335  = \399  & \245 ,
  \1336  = \973  & \248 ,
  \1337  = \610  & \249 ,
  \1338  = \1337  | \1336 ,
  \1339  = \1338  & \246 ,
  \1340  = \490  & \247 ,
  \1341  = \1340  | \1339 ,
  \1342  = \1341  & \244 ,
  \1343  = \400  & \245 ,
  \1344  = \974  & \248 ,
  \1345  = \611  & \249 ,
  \1346  = \1345  | \1344 ,
  \1347  = \1346  & \246 ,
  \1348  = \491  & \247 ,
  \1349  = \1348  | \1347 ,
  \1350  = \1349  & \244 ,
  \1351  = \401  & \245 ,
  \1352  = \975  & \248 ,
  \1353  = \612  & \249 ,
  \1354  = \1353  | \1352 ,
  \1355  = \1354  & \246 ,
  \1356  = \492  & \247 ,
  \1357  = \1356  | \1355 ,
  \1358  = \1357  & \244 ,
  \1359  = \402  & \245 ,
  \1360  = \946  & \248 ,
  \1361  = \613  & \249 ,
  \1362  = \1361  | \1360 ,
  \1363  = \1362  & \246 ,
  \1364  = \493  & \247 ,
  \1365  = \1364  | \1363 ,
  \1366  = \1365  & \244 ,
  \1367  = \403  & \245 ,
  \1368  = \434  & \246 ,
  \1369  = \614  & \247 ,
  \1370  = \1369  | \1368 ,
  \1371  = \1370  & \244 ,
  \1372  = \404  & \245 ,
  \1373  = \435  & \246 ,
  \1374  = \615  & \247 ,
  \1375  = \1374  | \1373 ,
  \1376  = \1375  & \244 ,
  \1377  = \405  & \245 ,
  \1378  = \436  & \246 ,
  \1379  = \616  & \247 ,
  \1380  = \1379  | \1378 ,
  \1381  = \1380  & \244 ,
  \1382  = \406  & \245 ,
  \1383  = \437  & \246 ,
  \1384  = \617  & \247 ,
  \1385  = \1384  | \1383 ,
  \1386  = \1385  & \244 ,
  \1387  = \407  & \245 ,
  \1388  = \438  & \246 ,
  \1389  = \618  & \247 ,
  \1390  = \1389  | \1388 ,
  \1391  = \1390  & \244 ,
  \1392  = \408  & \245 ,
  \1393  = \439  & \246 ,
  \1394  = \619  & \247 ,
  \1395  = \1394  | \1393 ,
  \1396  = \1395  & \244 ,
  \1397  = \409  & \245 ,
  \1398  = \440  & \246 ,
  \1399  = \620  & \247 ,
  \1400  = \1399  | \1398 ,
  \1401  = \1400  & \244 ,
  \1402  = \410  & \245 ,
  \1403  = \441  & \246 ,
  \1404  = \621  & \247 ,
  \1405  = \1404  | \1403 ,
  \1406  = \1405  & \244 ,
  \1407  = \411  & \245 ,
  \1408  = \442  & \246 ,
  \1409  = \622  & \247 ,
  \1410  = \1409  | \1408 ,
  \1411  = \1410  & \244 ,
  \1412  = \412  & \245 ,
  \1413  = \443  & \246 ,
  \1414  = \623  & \247 ,
  \1415  = \1414  | \1413 ,
  \1416  = \1415  & \244 ,
  \1417  = \413  & \245 ,
  \1418  = \444  & \246 ,
  \1419  = \624  & \247 ,
  \1420  = \1419  | \1418 ,
  \1421  = \1420  & \244 ,
  \1422  = \414  & \245 ,
  \1423  = \445  & \246 ,
  \1424  = \625  & \247 ,
  \1425  = \1424  | \1423 ,
  \1426  = \1425  & \244 ,
  \1427  = \415  & \245 ,
  \1428  = \446  & \246 ,
  \1429  = \626  & \247 ,
  \1430  = \1429  | \1428 ,
  \1431  = \1430  & \244 ,
  \1432  = \416  & \245 ,
  \1433  = \447  & \246 ,
  \1434  = \627  & \247 ,
  \1435  = \1434  | \1433 ,
  \1436  = \1435  & \244 ,
  \1437  = \417  & \245 ,
  \1438  = \448  & \246 ,
  \1439  = \628  & \247 ,
  \1440  = \1439  | \1438 ,
  \1441  = \1440  & \244 ,
  \1442  = \418  & \245 ,
  \1443  = \449  & \246 ,
  \1444  = \629  & \247 ,
  \1445  = \1444  | \1443 ,
  \1446  = \1445  & \244 ,
  \1447  = \419  & \245 ,
  \1448  = \450  & \246 ,
  \1449  = \630  & \247 ,
  \1450  = \1449  | \1448 ,
  \1451  = \1450  & \244 ,
  \1452  = \420  & \245 ,
  \1453  = \451  & \246 ,
  \1454  = \631  & \247 ,
  \1455  = \1454  | \1453 ,
  \1456  = \1455  & \244 ,
  \1457  = \421  & \245 ,
  \1458  = \452  & \246 ,
  \1459  = \632  & \247 ,
  \1460  = \1459  | \1458 ,
  \1461  = \1460  & \244 ,
  \1462  = \422  & \245 ,
  \1463  = \453  & \246 ,
  \1464  = \633  & \247 ,
  \1465  = \1464  | \1463 ,
  \1466  = \1465  & \244 ,
  \1467  = \423  & \245 ,
  \1468  = \454  & \246 ,
  \1469  = \634  & \247 ,
  \1470  = \1469  | \1468 ,
  \1471  = \1470  & \244 ,
  \1472  = \424  & \245 ,
  \1473  = \455  & \246 ,
  \1474  = \635  & \247 ,
  \1475  = \1474  | \1473 ,
  \1476  = \1475  & \244 ,
  \1477  = \425  & \245 ,
  \1478  = \456  & \246 ,
  \1479  = \636  & \247 ,
  \1480  = \1479  | \1478 ,
  \1481  = \1480  & \244 ,
  \1482  = \426  & \245 ,
  \1483  = \457  & \246 ,
  \1484  = \637  & \247 ,
  \1485  = \1484  | \1483 ,
  \1486  = \1485  & \244 ,
  \1487  = \427  & \245 ,
  \1488  = \458  & \246 ,
  \1489  = \638  & \247 ,
  \1490  = \1489  | \1488 ,
  \1491  = \1490  & \244 ,
  \1492  = \428  & \245 ,
  \1493  = \459  & \246 ,
  \1494  = \639  & \247 ,
  \1495  = \1494  | \1493 ,
  \1496  = \1495  & \244 ,
  \1497  = \429  & \245 ,
  \1498  = \460  & \246 ,
  \1499  = \640  & \247 ,
  \1500  = \1499  | \1498 ,
  \1501  = \1500  & \244 ,
  \1502  = \430  & \245 ,
  \1503  = \461  & \246 ,
  \1504  = \641  & \247 ,
  \1505  = \1504  | \1503 ,
  \1506  = \1505  & \244 ,
  \1507  = \431  & \245 ,
  \1508  = \462  & \246 ,
  \1509  = \642  & \247 ,
  \1510  = \1509  | \1508 ,
  \1511  = \1510  & \244 ,
  \1512  = \432  & \245 ,
  \1513  = \463  & \246 ,
  \1514  = \643  & \247 ,
  \1515  = \1514  | \1513 ,
  \1516  = \1515  & \244 ,
  \1517  = \433  & \245 ,
  \1518  = \1006  & \248 ,
  \1519  = \705  & \249 ,
  \1520  = \1519  | \1518 ,
  \1521  = \1520  & \246 ,
  \1522  = \674  & \247 ,
  \1523  = \1522  | \1521 ,
  \1524  = \1523  & \244 ,
  \1525  = \554  & \245 ,
  \1526  = \1007  & \248 ,
  \1527  = \706  & \249 ,
  \1528  = \1527  | \1526 ,
  \1529  = \1528  & \246 ,
  \1530  = \675  & \247 ,
  \1531  = \1530  | \1529 ,
  \1532  = \1531  & \244 ,
  \1533  = \555  & \245 ,
  \1534  = \1008  & \248 ,
  \1535  = \707  & \249 ,
  \1536  = \1535  | \1534 ,
  \1537  = \1536  & \246 ,
  \1538  = \676  & \247 ,
  \1539  = \1538  | \1537 ,
  \1540  = \1539  & \244 ,
  \1541  = \556  & \245 ,
  \1542  = \1009  & \248 ,
  \1543  = \708  & \249 ,
  \1544  = \1543  | \1542 ,
  \1545  = \1544  & \246 ,
  \1546  = \677  & \247 ,
  \1547  = \1546  | \1545 ,
  \1548  = \1547  & \244 ,
  \1549  = \557  & \245 ,
  \1550  = \1010  & \248 ,
  \1551  = \709  & \249 ,
  \1552  = \1551  | \1550 ,
  \1553  = \1552  & \246 ,
  \1554  = \678  & \247 ,
  \1555  = \1554  | \1553 ,
  \1556  = \1555  & \244 ,
  \1557  = \558  & \245 ,
  \1558  = \1011  & \248 ,
  \1559  = \710  & \249 ,
  \1560  = \1559  | \1558 ,
  \1561  = \1560  & \246 ,
  \1562  = \679  & \247 ,
  \1563  = \1562  | \1561 ,
  \1564  = \1563  & \244 ,
  \1565  = \559  & \245 ,
  \1566  = \1012  & \248 ,
  \1567  = \711  & \249 ,
  \1568  = \1567  | \1566 ,
  \1569  = \1568  & \246 ,
  \1570  = \680  & \247 ,
  \1571  = \1570  | \1569 ,
  \1572  = \1571  & \244 ,
  \1573  = \560  & \245 ,
  \1574  = \1013  & \248 ,
  \1575  = \712  & \249 ,
  \1576  = \1575  | \1574 ,
  \1577  = \1576  & \246 ,
  \1578  = \681  & \247 ,
  \1579  = \1578  | \1577 ,
  \1580  = \1579  & \244 ,
  \1581  = \561  & \245 ,
  \1582  = \1014  & \248 ,
  \1583  = \713  & \249 ,
  \1584  = \1583  | \1582 ,
  \1585  = \1584  & \246 ,
  \1586  = \682  & \247 ,
  \1587  = \1586  | \1585 ,
  \1588  = \1587  & \244 ,
  \1589  = \562  & \245 ,
  \1590  = \1015  & \248 ,
  \1591  = \714  & \249 ,
  \1592  = \1591  | \1590 ,
  \1593  = \1592  & \246 ,
  \1594  = \683  & \247 ,
  \1595  = \1594  | \1593 ,
  \1596  = \1595  & \244 ,
  \1597  = \563  & \245 ,
  \1598  = \1016  & \248 ,
  \1599  = \715  & \249 ,
  \1600  = \1599  | \1598 ,
  \1601  = \1600  & \246 ,
  \1602  = \684  & \247 ,
  \1603  = \1602  | \1601 ,
  \1604  = \1603  & \244 ,
  \1605  = \564  & \245 ,
  \1606  = \1017  & \248 ,
  \1607  = \716  & \249 ,
  \1608  = \1607  | \1606 ,
  \1609  = \1608  & \246 ,
  \1610  = \685  & \247 ,
  \1611  = \1610  | \1609 ,
  \1612  = \1611  & \244 ,
  \1613  = \565  & \245 ,
  \1614  = \1018  & \248 ,
  \1615  = \717  & \249 ,
  \1616  = \1615  | \1614 ,
  \1617  = \1616  & \246 ,
  \1618  = \686  & \247 ,
  \1619  = \1618  | \1617 ,
  \1620  = \1619  & \244 ,
  \1621  = \566  & \245 ,
  \1622  = \1019  & \248 ,
  \1623  = \718  & \249 ,
  \1624  = \1623  | \1622 ,
  \1625  = \1624  & \246 ,
  \1626  = \687  & \247 ,
  \1627  = \1626  | \1625 ,
  \1628  = \1627  & \244 ,
  \1629  = \567  & \245 ,
  \1630  = \1020  & \248 ,
  \1631  = \719  & \249 ,
  \1632  = \1631  | \1630 ,
  \1633  = \1632  & \246 ,
  \1634  = \688  & \247 ,
  \1635  = \1634  | \1633 ,
  \1636  = \1635  & \244 ,
  \1637  = \568  & \245 ,
  \1638  = \1021  & \248 ,
  \1639  = \720  & \249 ,
  \1640  = \1639  | \1638 ,
  \1641  = \1640  & \246 ,
  \1642  = \689  & \247 ,
  \1643  = \1642  | \1641 ,
  \1644  = \1643  & \244 ,
  \1645  = \569  & \245 ,
  \1646  = \1022  & \248 ,
  \1647  = \721  & \249 ,
  \1648  = \1647  | \1646 ,
  \1649  = \1648  & \246 ,
  \1650  = \690  & \247 ,
  \1651  = \1650  | \1649 ,
  \1652  = \1651  & \244 ,
  \1653  = \570  & \245 ,
  \1654  = \1023  & \248 ,
  \1655  = \722  & \249 ,
  \1656  = \1655  | \1654 ,
  \1657  = \1656  & \246 ,
  \1658  = \691  & \247 ,
  \1659  = \1658  | \1657 ,
  \1660  = \1659  & \244 ,
  \1661  = \571  & \245 ,
  \1662  = \1024  & \248 ,
  \1663  = \723  & \249 ,
  \1664  = \1663  | \1662 ,
  \1665  = \1664  & \246 ,
  \1666  = \692  & \247 ,
  \1667  = \1666  | \1665 ,
  \1668  = \1667  & \244 ,
  \1669  = \572  & \245 ,
  \1670  = \1025  & \248 ,
  \1671  = \724  & \249 ,
  \1672  = \1671  | \1670 ,
  \1673  = \1672  & \246 ,
  \1674  = \693  & \247 ,
  \1675  = \1674  | \1673 ,
  \1676  = \1675  & \244 ,
  \1677  = \573  & \245 ,
  \1678  = \1026  & \248 ,
  \1679  = \725  & \249 ,
  \1680  = \1679  | \1678 ,
  \1681  = \1680  & \246 ,
  \1682  = \694  & \247 ,
  \1683  = \1682  | \1681 ,
  \1684  = \1683  & \244 ,
  \1685  = \574  & \245 ,
  \1686  = \1027  & \248 ,
  \1687  = \726  & \249 ,
  \1688  = \1687  | \1686 ,
  \1689  = \1688  & \246 ,
  \1690  = \695  & \247 ,
  \1691  = \1690  | \1689 ,
  \1692  = \1691  & \244 ,
  \1693  = \575  & \245 ,
  \1694  = \1028  & \248 ,
  \1695  = \727  & \249 ,
  \1696  = \1695  | \1694 ,
  \1697  = \1696  & \246 ,
  \1698  = \696  & \247 ,
  \1699  = \1698  | \1697 ,
  \1700  = \1699  & \244 ,
  \1701  = \576  & \245 ,
  \1702  = \1029  & \248 ,
  \1703  = \728  & \249 ,
  \1704  = \1703  | \1702 ,
  \1705  = \1704  & \246 ,
  \1706  = \697  & \247 ,
  \1707  = \1706  | \1705 ,
  \1708  = \1707  & \244 ,
  \1709  = \577  & \245 ,
  \1710  = \1030  & \248 ,
  \1711  = \729  & \249 ,
  \1712  = \1711  | \1710 ,
  \1713  = \1712  & \246 ,
  \1714  = \698  & \247 ,
  \1715  = \1714  | \1713 ,
  \1716  = \1715  & \244 ,
  \1717  = \578  & \245 ,
  \1718  = \1031  & \248 ,
  \1719  = \730  & \249 ,
  \1720  = \1719  | \1718 ,
  \1721  = \1720  & \246 ,
  \1722  = \699  & \247 ,
  \1723  = \1722  | \1721 ,
  \1724  = \1723  & \244 ,
  \1725  = \579  & \245 ,
  \1726  = \1032  & \248 ,
  \1727  = \731  & \249 ,
  \1728  = \1727  | \1726 ,
  \1729  = \1728  & \246 ,
  \1730  = \700  & \247 ,
  \1731  = \1730  | \1729 ,
  \1732  = \1731  & \244 ,
  \1733  = \580  & \245 ,
  \1734  = \1033  & \248 ,
  \1735  = \732  & \249 ,
  \1736  = \1735  | \1734 ,
  \1737  = \1736  & \246 ,
  \1738  = \701  & \247 ,
  \1739  = \1738  | \1737 ,
  \1740  = \1739  & \244 ,
  \1741  = \581  & \245 ,
  \1742  = \1034  & \248 ,
  \1743  = \733  & \249 ,
  \1744  = \1743  | \1742 ,
  \1745  = \1744  & \246 ,
  \1746  = \702  & \247 ,
  \1747  = \1746  | \1745 ,
  \1748  = \1747  & \244 ,
  \1749  = \582  & \245 ,
  \1750  = \1035  & \248 ,
  \1751  = \734  & \249 ,
  \1752  = \1751  | \1750 ,
  \1753  = \1752  & \246 ,
  \1754  = \703  & \247 ,
  \1755  = \1754  | \1753 ,
  \1756  = \1755  & \244 ,
  \1757  = \583  & \245 ,
  \1758  = \976  & \248 ,
  \1759  = \644  & \249 ,
  \1760  = \1759  | \1758 ,
  \1761  = \1760  & \246 ,
  \1762  = \524  & \247 ,
  \1763  = \1762  | \1761 ,
  \1764  = \1763  & \244 ,
  \1765  = \494  & \245 ,
  \1766  = \977  & \248 ,
  \1767  = \645  & \249 ,
  \1768  = \1767  | \1766 ,
  \1769  = \1768  & \246 ,
  \1770  = \525  & \247 ,
  \1771  = \1770  | \1769 ,
  \1772  = \1771  & \244 ,
  \1773  = \495  & \245 ,
  \1774  = \978  & \248 ,
  \1775  = \646  & \249 ,
  \1776  = \1775  | \1774 ,
  \1777  = \1776  & \246 ,
  \1778  = \526  & \247 ,
  \1779  = \1778  | \1777 ,
  \1780  = \1779  & \244 ,
  \1781  = \496  & \245 ,
  \1782  = \979  & \248 ,
  \1783  = \647  & \249 ,
  \1784  = \1783  | \1782 ,
  \1785  = \1784  & \246 ,
  \1786  = \527  & \247 ,
  \1787  = \1786  | \1785 ,
  \1788  = \1787  & \244 ,
  \1789  = \497  & \245 ,
  \1790  = \980  & \248 ,
  \1791  = \648  & \249 ,
  \1792  = \1791  | \1790 ,
  \1793  = \1792  & \246 ,
  \1794  = \528  & \247 ,
  \1795  = \1794  | \1793 ,
  \1796  = \1795  & \244 ,
  \1797  = \498  & \245 ,
  \1798  = \981  & \248 ,
  \1799  = \649  & \249 ,
  \1800  = \1799  | \1798 ,
  \1801  = \1800  & \246 ,
  \1802  = \529  & \247 ,
  \1803  = \1802  | \1801 ,
  \1804  = \1803  & \244 ,
  \1805  = \499  & \245 ,
  \1806  = \982  & \248 ,
  \1807  = \650  & \249 ,
  \1808  = \1807  | \1806 ,
  \1809  = \1808  & \246 ,
  \1810  = \530  & \247 ,
  \1811  = \1810  | \1809 ,
  \1812  = \1811  & \244 ,
  \1813  = \500  & \245 ,
  \1814  = \983  & \248 ,
  \1815  = \651  & \249 ,
  \1816  = \1815  | \1814 ,
  \1817  = \1816  & \246 ,
  \1818  = \531  & \247 ,
  \1819  = \1818  | \1817 ,
  \1820  = \1819  & \244 ,
  \1821  = \501  & \245 ,
  \1822  = \984  & \248 ,
  \1823  = \652  & \249 ,
  \1824  = \1823  | \1822 ,
  \1825  = \1824  & \246 ,
  \1826  = \532  & \247 ,
  \1827  = \1826  | \1825 ,
  \1828  = \1827  & \244 ,
  \1829  = \502  & \245 ,
  \1830  = \985  & \248 ,
  \1831  = \653  & \249 ,
  \1832  = \1831  | \1830 ,
  \1833  = \1832  & \246 ,
  \1834  = \533  & \247 ,
  \1835  = \1834  | \1833 ,
  \1836  = \1835  & \244 ,
  \1837  = \503  & \245 ,
  \1838  = \986  & \248 ,
  \1839  = \654  & \249 ,
  \1840  = \1839  | \1838 ,
  \1841  = \1840  & \246 ,
  \1842  = \534  & \247 ,
  \1843  = \1842  | \1841 ,
  \1844  = \1843  & \244 ,
  \1845  = \504  & \245 ,
  \1846  = \987  & \248 ,
  \1847  = \655  & \249 ,
  \1848  = \1847  | \1846 ,
  \1849  = \1848  & \246 ,
  \1850  = \535  & \247 ,
  \1851  = \1850  | \1849 ,
  \1852  = \1851  & \244 ,
  \1853  = \505  & \245 ,
  \1854  = \988  & \248 ,
  \1855  = \656  & \249 ,
  \1856  = \1855  | \1854 ,
  \1857  = \1856  & \246 ,
  \1858  = \536  & \247 ,
  \1859  = \1858  | \1857 ,
  \1860  = \1859  & \244 ,
  \1861  = \506  & \245 ,
  \1862  = \989  & \248 ,
  \1863  = \657  & \249 ,
  \1864  = \1863  | \1862 ,
  \1865  = \1864  & \246 ,
  \1866  = \537  & \247 ,
  \1867  = \1866  | \1865 ,
  \1868  = \1867  & \244 ,
  \1869  = \507  & \245 ,
  \1870  = \990  & \248 ,
  \1871  = \658  & \249 ,
  \1872  = \1871  | \1870 ,
  \1873  = \1872  & \246 ,
  \1874  = \538  & \247 ,
  \1875  = \1874  | \1873 ,
  \1876  = \1875  & \244 ,
  \1877  = \508  & \245 ,
  \1878  = \991  & \248 ,
  \1879  = \659  & \249 ,
  \1880  = \1879  | \1878 ,
  \1881  = \1880  & \246 ,
  \1882  = \539  & \247 ,
  \1883  = \1882  | \1881 ,
  \1884  = \1883  & \244 ,
  \1885  = \509  & \245 ,
  \1886  = \992  & \248 ,
  \1887  = \660  & \249 ,
  \1888  = \1887  | \1886 ,
  \1889  = \1888  & \246 ,
  \1890  = \540  & \247 ,
  \1891  = \1890  | \1889 ,
  \1892  = \1891  & \244 ,
  \1893  = \510  & \245 ,
  \1894  = \993  & \248 ,
  \1895  = \661  & \249 ,
  \1896  = \1895  | \1894 ,
  \1897  = \1896  & \246 ,
  \1898  = \541  & \247 ,
  \1899  = \1898  | \1897 ,
  \1900  = \1899  & \244 ,
  \1901  = \511  & \245 ,
  \1902  = \994  & \248 ,
  \1903  = \662  & \249 ,
  \1904  = \1903  | \1902 ,
  \1905  = \1904  & \246 ,
  \1906  = \542  & \247 ,
  \1907  = \1906  | \1905 ,
  \1908  = \1907  & \244 ,
  \1909  = \512  & \245 ,
  \1910  = \995  & \248 ,
  \1911  = \663  & \249 ,
  \1912  = \1911  | \1910 ,
  \1913  = \1912  & \246 ,
  \1914  = \543  & \247 ,
  \1915  = \1914  | \1913 ,
  \1916  = \1915  & \244 ,
  \1917  = \513  & \245 ,
  \1918  = \996  & \248 ,
  \1919  = \664  & \249 ,
  \1920  = \1919  | \1918 ,
  \1921  = \1920  & \246 ,
  \1922  = \544  & \247 ,
  \1923  = \1922  | \1921 ,
  \1924  = \1923  & \244 ,
  \1925  = \514  & \245 ,
  \1926  = \997  & \248 ,
  \1927  = \665  & \249 ,
  \1928  = \1927  | \1926 ,
  \1929  = \1928  & \246 ,
  \1930  = \545  & \247 ,
  \1931  = \1930  | \1929 ,
  \1932  = \1931  & \244 ,
  \1933  = \515  & \245 ,
  \1934  = \998  & \248 ,
  \1935  = \666  & \249 ,
  \1936  = \1935  | \1934 ,
  \1937  = \1936  & \246 ,
  \1938  = \546  & \247 ,
  \1939  = \1938  | \1937 ,
  \1940  = \1939  & \244 ,
  \1941  = \516  & \245 ,
  \1942  = \999  & \248 ,
  \1943  = \667  & \249 ,
  \1944  = \1943  | \1942 ,
  \1945  = \1944  & \246 ,
  \1946  = \547  & \247 ,
  \1947  = \1946  | \1945 ,
  \1948  = \1947  & \244 ,
  \1949  = \517  & \245 ,
  \1950  = \1000  & \248 ,
  \1951  = \668  & \249 ,
  \1952  = \1951  | \1950 ,
  \1953  = \1952  & \246 ,
  \1954  = \548  & \247 ,
  \1955  = \1954  | \1953 ,
  \1956  = \1955  & \244 ,
  \1957  = \518  & \245 ,
  \1958  = \1001  & \248 ,
  \1959  = \669  & \249 ,
  \1960  = \1959  | \1958 ,
  \1961  = \1960  & \246 ,
  \1962  = \549  & \247 ,
  \1963  = \1962  | \1961 ,
  \1964  = \1963  & \244 ,
  \1965  = \519  & \245 ,
  \1966  = \1002  & \248 ,
  \1967  = \670  & \249 ,
  \1968  = \1967  | \1966 ,
  \1969  = \1968  & \246 ,
  \1970  = \550  & \247 ,
  \1971  = \1970  | \1969 ,
  \1972  = \1971  & \244 ,
  \1973  = \520  & \245 ,
  \1974  = \1003  & \248 ,
  \1975  = \671  & \249 ,
  \1976  = \1975  | \1974 ,
  \1977  = \1976  & \246 ,
  \1978  = \551  & \247 ,
  \1979  = \1978  | \1977 ,
  \1980  = \1979  & \244 ,
  \1981  = \521  & \245 ,
  \1982  = \1004  & \248 ,
  \1983  = \672  & \249 ,
  \1984  = \1983  | \1982 ,
  \1985  = \1984  & \246 ,
  \1986  = \552  & \247 ,
  \1987  = \1986  | \1985 ,
  \1988  = \1987  & \244 ,
  \1989  = \522  & \245 ,
  \1990  = \1005  & \248 ,
  \1991  = \673  & \249 ,
  \1992  = \1991  | \1990 ,
  \1993  = \1992  & \246 ,
  \1994  = \553  & \247 ,
  \1995  = \1994  | \1993 ,
  \1996  = \1995  & \244 ,
  \1997  = \523  & \245 ,
  \1998  = \885  & \372 ,
  \1999  = \915  & \373 ,
  \[100]  = \1215  | \1214 ,
  \[101]  = \1223  | \1222 ,
  \[102]  = \1231  | \1230 ,
  \[103]  = \1239  | \1238 ,
  \[104]  = \1247  | \1246 ,
  \[105]  = \1255  | \1254 ,
  \[106]  = \1263  | \1262 ,
  \[107]  = \1271  | \1270 ,
  \[108]  = \1279  | \1278 ,
  \[109]  = \1287  | \1286 ,
  \[110]  = \1295  | \1294 ,
  \[111]  = \1303  | \1302 ,
  \[112]  = \1311  | \1310 ,
  \[113]  = \1319  | \1318 ,
  \[114]  = \1327  | \1326 ,
  \[115]  = \1335  | \1334 ,
  \[116]  = \1343  | \1342 ,
  \[117]  = \1351  | \1350 ,
  \[118]  = \1359  | \1358 ,
  \[119]  = \1367  | \1366 ,
  \[120]  = \154 ,
  \[121]  = \155 ,
  \[122]  = \156 ,
  \[123]  = \157 ,
  \[124]  = \158 ,
  \[125]  = \159 ,
  \[126]  = \160 ,
  \[127]  = \161 ,
  \[128]  = \162 ,
  \[129]  = \163 ,
  \2000  = \1999  | \1998 ,
  \2001  = \248  & \246 ,
  \2002  = \2001  & \244 ,
  \2003  = \794  & \310 ,
  \2004  = \824  & \311 ,
  \2005  = \2004  | \2003 ,
  \2006  = \248  & \246 ,
  \2007  = \2006  & \244 ,
  \2008  = \884  & \372 ,
  \2009  = \914  & \373 ,
  \2010  = \2009  | \2008 ,
  \2011  = \248  & \246 ,
  \2012  = \2011  & \244 ,
  \2013  = \793  & \310 ,
  \2014  = \823  & \311 ,
  \2015  = \2014  | \2013 ,
  \2016  = \248  & \246 ,
  \2017  = \2016  & \244 ,
  \2018  = \883  & \372 ,
  \2019  = \913  & \373 ,
  \2020  = \2019  | \2018 ,
  \2021  = \248  & \246 ,
  \2022  = \2021  & \244 ,
  \2023  = \792  & \310 ,
  \2024  = \822  & \311 ,
  \2025  = \2024  | \2023 ,
  \2026  = \248  & \246 ,
  \2027  = \2026  & \244 ,
  \2028  = \882  & \372 ,
  \2029  = \912  & \373 ,
  \2030  = \2029  | \2028 ,
  \2031  = \248  & \246 ,
  \2032  = \2031  & \244 ,
  \2033  = \791  & \310 ,
  \2034  = \821  & \311 ,
  \2035  = \2034  | \2033 ,
  \2036  = \248  & \246 ,
  \2037  = \2036  & \244 ,
  \2038  = \881  & \372 ,
  \2039  = \911  & \373 ,
  \2040  = \2039  | \2038 ,
  \2041  = \248  & \246 ,
  \2042  = \2041  & \244 ,
  \2043  = \790  & \310 ,
  \2044  = \820  & \311 ,
  \2045  = \2044  | \2043 ,
  \2046  = \248  & \246 ,
  \2047  = \2046  & \244 ,
  \2048  = \880  & \372 ,
  \2049  = \910  & \373 ,
  \2050  = \2049  | \2048 ,
  \2051  = \248  & \246 ,
  \2052  = \2051  & \244 ,
  \2053  = \789  & \310 ,
  \2054  = \819  & \311 ,
  \2055  = \2054  | \2053 ,
  \2056  = \248  & \246 ,
  \2057  = \2056  & \244 ,
  \2058  = \879  & \372 ,
  \2059  = \909  & \373 ,
  \2060  = \2059  | \2058 ,
  \2061  = \248  & \246 ,
  \2062  = \2061  & \244 ,
  \2063  = \788  & \310 ,
  \2064  = \818  & \311 ,
  \2065  = \2064  | \2063 ,
  \2066  = \248  & \246 ,
  \2067  = \2066  & \244 ,
  \2068  = \878  & \372 ,
  \2069  = \908  & \373 ,
  \[130]  = \164 ,
  \2070  = \2069  | \2068 ,
  \2071  = \248  & \246 ,
  \2072  = \2071  & \244 ,
  \2073  = \787  & \310 ,
  \2074  = \817  & \311 ,
  \2075  = \2074  | \2073 ,
  \2076  = \248  & \246 ,
  \2077  = \2076  & \244 ,
  \2078  = \877  & \372 ,
  \2079  = \907  & \373 ,
  \[131]  = \165 ,
  \2080  = \2079  | \2078 ,
  \2081  = \248  & \246 ,
  \2082  = \2081  & \244 ,
  \2083  = \786  & \310 ,
  \2084  = \816  & \311 ,
  \2085  = \2084  | \2083 ,
  \2086  = \248  & \246 ,
  \2087  = \2086  & \244 ,
  \2088  = \876  & \372 ,
  \2089  = \906  & \373 ,
  \[132]  = \166 ,
  \2090  = \2089  | \2088 ,
  \2091  = \248  & \246 ,
  \2092  = \2091  & \244 ,
  \2093  = \785  & \310 ,
  \2094  = \815  & \311 ,
  \2095  = \2094  | \2093 ,
  \2096  = \248  & \246 ,
  \2097  = \2096  & \244 ,
  \2098  = \875  & \372 ,
  \2099  = \905  & \373 ,
  \[133]  = \167 ,
  \[134]  = \168 ,
  \[135]  = \169 ,
  \[136]  = \170 ,
  \[137]  = \171 ,
  \[138]  = \172 ,
  \[139]  = \173 ,
  \2100  = \2099  | \2098 ,
  \2101  = \248  & \246 ,
  \2102  = \2101  & \244 ,
  \2103  = \784  & \310 ,
  \2104  = \814  & \311 ,
  \2105  = \2104  | \2103 ,
  \2106  = \248  & \246 ,
  \2107  = \2106  & \244 ,
  \2108  = \874  & \372 ,
  \2109  = \904  & \373 ,
  \2110  = \2109  | \2108 ,
  \2111  = \248  & \246 ,
  \2112  = \2111  & \244 ,
  \2113  = \783  & \310 ,
  \2114  = \813  & \311 ,
  \2115  = \2114  | \2113 ,
  \2116  = \248  & \246 ,
  \2117  = \2116  & \244 ,
  \2118  = \873  & \372 ,
  \2119  = \903  & \373 ,
  \2120  = \2119  | \2118 ,
  \2121  = \248  & \246 ,
  \2122  = \2121  & \244 ,
  \2123  = \782  & \310 ,
  \2124  = \812  & \311 ,
  \2125  = \2124  | \2123 ,
  \2126  = \248  & \246 ,
  \2127  = \2126  & \244 ,
  \2128  = \872  & \372 ,
  \2129  = \902  & \373 ,
  \2130  = \2129  | \2128 ,
  \2131  = \248  & \246 ,
  \2132  = \2131  & \244 ,
  \2133  = \781  & \310 ,
  \2134  = \811  & \311 ,
  \2135  = \2134  | \2133 ,
  \2136  = \248  & \246 ,
  \2137  = \2136  & \244 ,
  \2138  = \871  & \372 ,
  \2139  = \901  & \373 ,
  \2140  = \2139  | \2138 ,
  \2141  = \248  & \246 ,
  \2142  = \2141  & \244 ,
  \2143  = \780  & \310 ,
  \2144  = \810  & \311 ,
  \2145  = \2144  | \2143 ,
  \2146  = \248  & \246 ,
  \2147  = \2146  & \244 ,
  \2148  = \870  & \372 ,
  \2149  = \900  & \373 ,
  \2150  = \2149  | \2148 ,
  \2151  = \248  & \246 ,
  \2152  = \2151  & \244 ,
  \2153  = \779  & \310 ,
  \2154  = \809  & \311 ,
  \2155  = \2154  | \2153 ,
  \2156  = \248  & \246 ,
  \2157  = \2156  & \244 ,
  \2158  = \869  & \372 ,
  \2159  = \899  & \373 ,
  \2160  = \2159  | \2158 ,
  \2161  = \248  & \246 ,
  \2162  = \2161  & \244 ,
  \2163  = \778  & \310 ,
  \2164  = \808  & \311 ,
  \2165  = \2164  | \2163 ,
  \2166  = \248  & \246 ,
  \2167  = \2166  & \244 ,
  \2168  = \868  & \372 ,
  \2169  = \898  & \373 ,
  \[140]  = \174 ,
  \2170  = \2169  | \2168 ,
  \2171  = \248  & \246 ,
  \2172  = \2171  & \244 ,
  \2173  = \777  & \310 ,
  \2174  = \807  & \311 ,
  \2175  = \2174  | \2173 ,
  \2176  = \248  & \246 ,
  \2177  = \2176  & \244 ,
  \2178  = \867  & \372 ,
  \2179  = \897  & \373 ,
  \[141]  = \175 ,
  \2180  = \2179  | \2178 ,
  \2181  = \248  & \246 ,
  \2182  = \2181  & \244 ,
  \2183  = \776  & \310 ,
  \2184  = \806  & \311 ,
  \2185  = \2184  | \2183 ,
  \2186  = \248  & \246 ,
  \2187  = \2186  & \244 ,
  \2188  = \866  & \372 ,
  \2189  = \896  & \373 ,
  \[142]  = \176 ,
  \2190  = \2189  | \2188 ,
  \2191  = \248  & \246 ,
  \2192  = \2191  & \244 ,
  \2193  = \775  & \310 ,
  \2194  = \805  & \311 ,
  \2195  = \2194  | \2193 ,
  \2196  = \248  & \246 ,
  \2197  = \2196  & \244 ,
  \2198  = \865  & \372 ,
  \2199  = \895  & \373 ,
  \[143]  = \177 ,
  \[144]  = \178 ,
  \[145]  = \179 ,
  \[146]  = \180 ,
  \[147]  = \181 ,
  \[148]  = \182 ,
  \[149]  = \183 ,
  \2200  = \2199  | \2198 ,
  \2201  = \248  & \246 ,
  \2202  = \2201  & \244 ,
  \2203  = \774  & \310 ,
  \2204  = \804  & \311 ,
  \2205  = \2204  | \2203 ,
  \2206  = \248  & \246 ,
  \2207  = \2206  & \244 ,
  \2208  = \864  & \372 ,
  \2209  = \894  & \373 ,
  \2210  = \2209  | \2208 ,
  \2211  = \248  & \246 ,
  \2212  = \2211  & \244 ,
  \2213  = \773  & \310 ,
  \2214  = \803  & \311 ,
  \2215  = \2214  | \2213 ,
  \2216  = \248  & \246 ,
  \2217  = \2216  & \244 ,
  \2218  = \863  & \372 ,
  \2219  = \893  & \373 ,
  \2220  = \2219  | \2218 ,
  \2221  = \248  & \246 ,
  \2222  = \2221  & \244 ,
  \2223  = \772  & \310 ,
  \2224  = \802  & \311 ,
  \2225  = \2224  | \2223 ,
  \2226  = \248  & \246 ,
  \2227  = \2226  & \244 ,
  \2228  = \862  & \372 ,
  \2229  = \892  & \373 ,
  \2230  = \2229  | \2228 ,
  \2231  = \248  & \246 ,
  \2232  = \2231  & \244 ,
  \2233  = \771  & \310 ,
  \2234  = \801  & \311 ,
  \2235  = \2234  | \2233 ,
  \2236  = \248  & \246 ,
  \2237  = \2236  & \244 ,
  \2238  = \861  & \372 ,
  \2239  = \891  & \373 ,
  \2240  = \2239  | \2238 ,
  \2241  = \248  & \246 ,
  \2242  = \2241  & \244 ,
  \2243  = \770  & \310 ,
  \2244  = \800  & \311 ,
  \2245  = \2244  | \2243 ,
  \2246  = \248  & \246 ,
  \2247  = \2246  & \244 ,
  \2248  = \860  & \372 ,
  \2249  = \890  & \373 ,
  \2250  = \2249  | \2248 ,
  \2251  = \248  & \246 ,
  \2252  = \2251  & \244 ,
  \2253  = \769  & \310 ,
  \2254  = \799  & \311 ,
  \2255  = \2254  | \2253 ,
  \2256  = \248  & \246 ,
  \2257  = \2256  & \244 ,
  \2258  = \859  & \372 ,
  \2259  = \889  & \373 ,
  \2260  = \2259  | \2258 ,
  \2261  = \248  & \246 ,
  \2262  = \2261  & \244 ,
  \2263  = \768  & \310 ,
  \2264  = \798  & \311 ,
  \2265  = \2264  | \2263 ,
  \2266  = \248  & \246 ,
  \2267  = \2266  & \244 ,
  \2268  = \858  & \372 ,
  \2269  = \888  & \373 ,
  \[150]  = \184 ,
  \2270  = \2269  | \2268 ,
  \2271  = \248  & \246 ,
  \2272  = \2271  & \244 ,
  \2273  = \767  & \310 ,
  \2274  = \797  & \311 ,
  \2275  = \2274  | \2273 ,
  \2276  = \248  & \246 ,
  \2277  = \2276  & \244 ,
  \2278  = \857  & \372 ,
  \2279  = \887  & \373 ,
  \[151]  = \185 ,
  \2280  = \2279  | \2278 ,
  \2281  = \248  & \246 ,
  \2282  = \2281  & \244 ,
  \2283  = \766  & \310 ,
  \2284  = \796  & \311 ,
  \2285  = \2284  | \2283 ,
  \2286  = \248  & \246 ,
  \2287  = \2286  & \244 ,
  \2288  = \856  & \372 ,
  \2289  = \886  & \373 ,
  \[152]  = \186 ,
  \2290  = \2289  | \2288 ,
  \2291  = \248  & \246 ,
  \2292  = \2291  & \244 ,
  \2293  = \765  & \310 ,
  \2294  = \795  & \311 ,
  \2295  = \2294  | \2293 ,
  \2296  = \248  & \246 ,
  \2297  = \2296  & \244 ,
  \2298  = \854  & \370 ,
  \2299  = \855  & \371 ,
  \[153]  = \187 ,
  \[154]  = \188 ,
  \[155]  = \189 ,
  \[156]  = \190 ,
  \[157]  = \191 ,
  \[158]  = \192 ,
  \[159]  = \193 ,
  \2300  = \2299  | \2298 ,
  \2301  = \2300  & \368 ,
  \2302  = \853  & \369 ,
  \2303  = \2302  | \2301 ,
  \2304  = \2303  & \366 ,
  \2305  = \852  & \367 ,
  \2306  = \2305  | \2304 ,
  \2307  = \2306  & \364 ,
  \2308  = \851  & \365 ,
  \2309  = \2308  | \2307 ,
  \2310  = \2309  & \362 ,
  \2311  = \850  & \363 ,
  \2312  = \2311  | \2310 ,
  \2313  = \2312  & \360 ,
  \2314  = \849  & \361 ,
  \2315  = \2314  | \2313 ,
  \2316  = \2315  & \358 ,
  \2317  = \848  & \359 ,
  \2318  = \2317  | \2316 ,
  \2319  = \2318  & \356 ,
  \2320  = \847  & \357 ,
  \2321  = \2320  | \2319 ,
  \2322  = \2321  & \354 ,
  \2323  = \846  & \355 ,
  \2324  = \2323  | \2322 ,
  \2325  = \2324  & \352 ,
  \2326  = \845  & \353 ,
  \2327  = \2326  | \2325 ,
  \2328  = \2327  & \350 ,
  \2329  = \844  & \351 ,
  \2330  = \2329  | \2328 ,
  \2331  = \2330  & \348 ,
  \2332  = \843  & \349 ,
  \2333  = \2332  | \2331 ,
  \2334  = \2333  & \346 ,
  \2335  = \842  & \347 ,
  \2336  = \2335  | \2334 ,
  \2337  = \2336  & \344 ,
  \2338  = \841  & \345 ,
  \2339  = \2338  | \2337 ,
  \2340  = \2339  & \342 ,
  \2341  = \840  & \343 ,
  \2342  = \2341  | \2340 ,
  \2343  = \2342  & \340 ,
  \2344  = \839  & \341 ,
  \2345  = \2344  | \2343 ,
  \2346  = \2345  & \338 ,
  \2347  = \838  & \339 ,
  \2348  = \2347  | \2346 ,
  \2349  = \2348  & \336 ,
  \2350  = \837  & \337 ,
  \2351  = \2350  | \2349 ,
  \2352  = \2351  & \334 ,
  \2353  = \836  & \335 ,
  \2354  = \2353  | \2352 ,
  \2355  = \2354  & \332 ,
  \2356  = \835  & \333 ,
  \2357  = \2356  | \2355 ,
  \2358  = \2357  & \330 ,
  \2359  = \834  & \331 ,
  \2360  = \2359  | \2358 ,
  \2361  = \2360  & \328 ,
  \2362  = \833  & \329 ,
  \2363  = \2362  | \2361 ,
  \2364  = \2363  & \326 ,
  \2365  = \832  & \327 ,
  \2366  = \2365  | \2364 ,
  \2367  = \2366  & \324 ,
  \2368  = \831  & \325 ,
  \2369  = \2368  | \2367 ,
  \[160]  = \194 ,
  \2370  = \2369  & \322 ,
  \2371  = \830  & \323 ,
  \2372  = \2371  | \2370 ,
  \2373  = \2372  & \320 ,
  \2374  = \829  & \321 ,
  \2375  = \2374  | \2373 ,
  \2376  = \2375  & \318 ,
  \2377  = \828  & \319 ,
  \2378  = \2377  | \2376 ,
  \2379  = \2378  & \316 ,
  \[161]  = \195 ,
  \2380  = \827  & \317 ,
  \2381  = \2380  | \2379 ,
  \2382  = \2381  & \314 ,
  \2383  = \826  & \315 ,
  \2384  = \2383  | \2382 ,
  \2385  = \2384  & \312 ,
  \2386  = \825  & \313 ,
  \2387  = \2386  | \2385 ,
  \2388  = \248  & \246 ,
  \2389  = \2388  & \244 ,
  \[162]  = \196 ,
  \2390  = \763  & \308 ,
  \2391  = \764  & \309 ,
  \2392  = \2391  | \2390 ,
  \2393  = \2392  & \306 ,
  \2394  = \762  & \307 ,
  \2395  = \2394  | \2393 ,
  \2396  = \2395  & \304 ,
  \2397  = \761  & \305 ,
  \2398  = \2397  | \2396 ,
  \2399  = \2398  & \302 ,
  \[163]  = \197 ,
  \[164]  = \198 ,
  \[165]  = \199 ,
  \[166]  = \200 ,
  \[167]  = \201 ,
  \[168]  = \202 ,
  \[169]  = \203 ,
  \2400  = \760  & \303 ,
  \2401  = \2400  | \2399 ,
  \2402  = \2401  & \300 ,
  \2403  = \759  & \301 ,
  \2404  = \2403  | \2402 ,
  \2405  = \2404  & \298 ,
  \2406  = \758  & \299 ,
  \2407  = \2406  | \2405 ,
  \2408  = \2407  & \296 ,
  \2409  = \757  & \297 ,
  \2410  = \2409  | \2408 ,
  \2411  = \2410  & \294 ,
  \2412  = \756  & \295 ,
  \2413  = \2412  | \2411 ,
  \2414  = \2413  & \292 ,
  \2415  = \755  & \293 ,
  \2416  = \2415  | \2414 ,
  \2417  = \2416  & \290 ,
  \2418  = \754  & \291 ,
  \2419  = \2418  | \2417 ,
  \2420  = \2419  & \288 ,
  \2421  = \753  & \289 ,
  \2422  = \2421  | \2420 ,
  \2423  = \2422  & \286 ,
  \2424  = \752  & \287 ,
  \2425  = \2424  | \2423 ,
  \2426  = \2425  & \284 ,
  \2427  = \751  & \285 ,
  \2428  = \2427  | \2426 ,
  \2429  = \2428  & \282 ,
  \2430  = \750  & \283 ,
  \2431  = \2430  | \2429 ,
  \2432  = \2431  & \280 ,
  \2433  = \749  & \281 ,
  \2434  = \2433  | \2432 ,
  \2435  = \2434  & \278 ,
  \2436  = \748  & \279 ,
  \2437  = \2436  | \2435 ,
  \2438  = \2437  & \276 ,
  \2439  = \747  & \277 ,
  \2440  = \2439  | \2438 ,
  \2441  = \2440  & \274 ,
  \2442  = \746  & \275 ,
  \2443  = \2442  | \2441 ,
  \2444  = \2443  & \272 ,
  \2445  = \745  & \273 ,
  \2446  = \2445  | \2444 ,
  \2447  = \2446  & \270 ,
  \2448  = \744  & \271 ,
  \2449  = \2448  | \2447 ,
  \2450  = \2449  & \268 ,
  \2451  = \743  & \269 ,
  \2452  = \2451  | \2450 ,
  \2453  = \2452  & \266 ,
  \2454  = \742  & \267 ,
  \2455  = \2454  | \2453 ,
  \2456  = \2455  & \264 ,
  \2457  = \741  & \265 ,
  \2458  = \2457  | \2456 ,
  \2459  = \2458  & \262 ,
  \2460  = \740  & \263 ,
  \2461  = \2460  | \2459 ,
  \2462  = \2461  & \260 ,
  \2463  = \739  & \261 ,
  \2464  = \2463  | \2462 ,
  \2465  = \2464  & \258 ,
  \2466  = \738  & \259 ,
  \2467  = \2466  | \2465 ,
  \2468  = \2467  & \256 ,
  \2469  = \737  & \257 ,
  \[170]  = \204 ,
  \2470  = \2469  | \2468 ,
  \2471  = \2470  & \254 ,
  \2472  = \736  & \255 ,
  \2473  = \2472  | \2471 ,
  \2474  = \2473  & \252 ,
  \2475  = \735  & \253 ,
  \2476  = \2475  | \2474 ,
  \2477  = \2476  & \250 ,
  \2478  = \704  & \251 ,
  \2479  = \2478  | \2477 ,
  \[171]  = \205 ,
  \2480  = \248  & \246 ,
  \2481  = \2480  & \244 ,
  \[172]  = \206 ,
  \[173]  = \207 ,
  \[174]  = \208 ,
  \[175]  = \209 ,
  \[176]  = \210 ,
  \[177]  = \211 ,
  \[178]  = \212 ,
  \[179]  = \213 ,
  \[180]  = \214 ,
  \[181]  = \215 ,
  \[182]  = \216 ,
  \[183]  = \217 ,
  \[184]  = \218 ,
  \[185]  = \219 ,
  \[186]  = \220 ,
  \[187]  = \221 ,
  \[188]  = \222 ,
  \124  = \[90] ,
  \125  = \[91] ,
  \126  = \[92] ,
  \[189]  = \223 ,
  \127  = \[93] ,
  \128  = \[94] ,
  \129  = \[95] ,
  \130  = \[96] ,
  \131  = \[97] ,
  \132  = \[98] ,
  \133  = \[99] ,
  \134  = \[100] ,
  \135  = \[101] ,
  \136  = \[102] ,
  \137  = \[103] ,
  \138  = \[104] ,
  \139  = \[105] ,
  \140  = \[106] ,
  \141  = \[107] ,
  \142  = \[108] ,
  \143  = \[109] ,
  \144  = \[110] ,
  \145  = \[111] ,
  \146  = \[112] ,
  \147  = \[113] ,
  \148  = \[114] ,
  \149  = \[115] ,
  \150  = \[116] ,
  \151  = \[117] ,
  \152  = \[118] ,
  \153  = \[119] ,
  \154  = \1372  | \1371 ,
  \155  = \1377  | \1376 ,
  \156  = \1382  | \1381 ,
  \157  = \1387  | \1386 ,
  \158  = \1392  | \1391 ,
  \159  = \1397  | \1396 ,
  \160  = \1402  | \1401 ,
  \161  = \1407  | \1406 ,
  \162  = \1412  | \1411 ,
  \163  = \1417  | \1416 ,
  \164  = \1422  | \1421 ,
  \165  = \1427  | \1426 ,
  \166  = \1432  | \1431 ,
  \167  = \1437  | \1436 ,
  \168  = \1442  | \1441 ,
  \169  = \1447  | \1446 ,
  \170  = \1452  | \1451 ,
  \171  = \1457  | \1456 ,
  \172  = \1462  | \1461 ,
  \173  = \1467  | \1466 ,
  \174  = \1472  | \1471 ,
  \175  = \1477  | \1476 ,
  \176  = \1482  | \1481 ,
  \177  = \1487  | \1486 ,
  \178  = \1492  | \1491 ,
  \179  = \1497  | \1496 ,
  \180  = \1502  | \1501 ,
  \181  = \1507  | \1506 ,
  \182  = \1512  | \1511 ,
  \183  = \1517  | \1516 ,
  \184  = \1525  | \1524 ,
  \185  = \1533  | \1532 ,
  \186  = \1541  | \1540 ,
  \187  = \1549  | \1548 ,
  \188  = \1557  | \1556 ,
  \189  = \1565  | \1564 ,
  \190  = \1573  | \1572 ,
  \191  = \1581  | \1580 ,
  \192  = \1589  | \1588 ,
  \193  = \1597  | \1596 ,
  \194  = \1605  | \1604 ,
  \195  = \1613  | \1612 ,
  \196  = \1621  | \1620 ,
  \[190]  = \224 ,
  \197  = \1629  | \1628 ,
  \198  = \1637  | \1636 ,
  \199  = \1645  | \1644 ,
  \[191]  = \225 ,
  \[192]  = \226 ,
  \[193]  = \227 ,
  \[194]  = \228 ,
  \[195]  = \229 ,
  \[196]  = \230 ,
  \200  = \1653  | \1652 ,
  \201  = \1661  | \1660 ,
  \202  = \1669  | \1668 ,
  \203  = \1677  | \1676 ,
  \204  = \1685  | \1684 ,
  \205  = \1693  | \1692 ,
  \206  = \1701  | \1700 ,
  \[197]  = \231 ,
  \207  = \1709  | \1708 ,
  \208  = \1717  | \1716 ,
  \209  = \1725  | \1724 ,
  \210  = \1733  | \1732 ,
  \211  = \1741  | \1740 ,
  \212  = \1749  | \1748 ,
  \213  = \1757  | \1756 ,
  \214  = \1765  | \1764 ,
  \215  = \1773  | \1772 ,
  \216  = \1781  | \1780 ,
  \[198]  = \232 ,
  \217  = \1789  | \1788 ,
  \218  = \1797  | \1796 ,
  \219  = \1805  | \1804 ,
  \220  = \1813  | \1812 ,
  \221  = \1821  | \1820 ,
  \222  = \1829  | \1828 ,
  \223  = \1837  | \1836 ,
  \224  = \1845  | \1844 ,
  \225  = \1853  | \1852 ,
  \226  = \1861  | \1860 ,
  \[199]  = \233 ,
  \227  = \1869  | \1868 ,
  \228  = \1877  | \1876 ,
  \229  = \1885  | \1884 ,
  \230  = \1893  | \1892 ,
  \231  = \1901  | \1900 ,
  \232  = \1909  | \1908 ,
  \233  = \1917  | \1916 ,
  \234  = \1925  | \1924 ,
  \235  = \1933  | \1932 ,
  \236  = \1941  | \1940 ,
  \237  = \1949  | \1948 ,
  \238  = \1957  | \1956 ,
  \239  = \1965  | \1964 ,
  \240  = \1973  | \1972 ,
  \241  = \1981  | \1980 ,
  \242  = \1989  | \1988 ,
  \243  = \1997  | \1996 ,
  \244  = ~\245 ,
  \245  = \1 ,
  \246  = ~\247 ,
  \247  = ~\2 ,
  \248  = ~\249 ,
  \249  = \3 ,
  \250  = ~\251 ,
  \251  = (~\33  & \123 ) | (\33  & ~\123 ),
  \252  = ~\253 ,
  \253  = (~\32  & \122 ) | (\32  & ~\122 ),
  \254  = ~\255 ,
  \255  = (~\31  & \121 ) | (\31  & ~\121 ),
  \256  = ~\257 ,
  \257  = (~\30  & \120 ) | (\30  & ~\120 ),
  \258  = ~\259 ,
  \259  = (~\29  & \119 ) | (\29  & ~\119 ),
  \260  = ~\261 ,
  \261  = (~\28  & \118 ) | (\28  & ~\118 ),
  \262  = ~\263 ,
  \263  = (~\27  & \117 ) | (\27  & ~\117 ),
  \264  = ~\265 ,
  \265  = (~\26  & \116 ) | (\26  & ~\116 ),
  \266  = ~\267 ,
  \267  = (~\25  & \115 ) | (\25  & ~\115 ),
  \268  = ~\269 ,
  \269  = (~\24  & \114 ) | (\24  & ~\114 ),
  \270  = ~\271 ,
  \271  = (~\23  & \113 ) | (\23  & ~\113 ),
  \272  = ~\273 ,
  \273  = (~\22  & \112 ) | (\22  & ~\112 ),
  \274  = ~\275 ,
  \275  = (~\21  & \111 ) | (\21  & ~\111 ),
  \276  = ~\277 ,
  \277  = (~\20  & \110 ) | (\20  & ~\110 ),
  \278  = ~\279 ,
  \279  = (~\19  & \109 ) | (\19  & ~\109 ),
  \280  = ~\281 ,
  \281  = (~\18  & \108 ) | (\18  & ~\108 ),
  \282  = ~\283 ,
  \283  = (~\17  & \107 ) | (\17  & ~\107 ),
  \284  = ~\285 ,
  \285  = (~\16  & \106 ) | (\16  & ~\106 ),
  \286  = ~\287 ,
  \287  = (~\15  & \105 ) | (\15  & ~\105 ),
  \288  = ~\289 ,
  \289  = (~\14  & \104 ) | (\14  & ~\104 ),
  \290  = ~\291 ,
  \291  = (~\13  & \103 ) | (\13  & ~\103 ),
  \292  = ~\293 ,
  \293  = (~\12  & \102 ) | (\12  & ~\102 ),
  \294  = ~\295 ,
  \295  = (~\11  & \101 ) | (\11  & ~\101 ),
  \296  = ~\297 ,
  \297  = (~\10  & \100 ) | (\10  & ~\100 ),
  \298  = ~\299 ,
  \299  = (~\9  & \99 ) | (\9  & ~\99 ),
  \300  = ~\301 ,
  \301  = (~\8  & \98 ) | (\8  & ~\98 ),
  \302  = ~\303 ,
  \303  = (~\7  & \97 ) | (\7  & ~\97 ),
  \304  = ~\305 ,
  \305  = (~\6  & \96 ) | (\6  & ~\96 ),
  \306  = ~\307 ,
  \307  = (~\5  & \95 ) | (\5  & ~\95 ),
  \308  = ~\309 ,
  \309  = (~\4  & \94 ) | (\4  & ~\94 ),
  \310  = ~\311 ,
  \311  = \1036 ,
  \312  = ~\313 ,
  \313  = (~\33  & \93 ) | (\33  & ~\93 ),
  \314  = ~\315 ,
  \315  = (~\32  & \92 ) | (\32  & ~\92 ),
  \316  = ~\317 ,
  \317  = (~\31  & \91 ) | (\31  & ~\91 ),
  \318  = ~\319 ,
  \319  = (~\30  & \90 ) | (\30  & ~\90 ),
  \320  = ~\321 ,
  \321  = (~\29  & \89 ) | (\29  & ~\89 ),
  \322  = ~\323 ,
  \323  = (~\28  & \88 ) | (\28  & ~\88 ),
  \324  = ~\325 ,
  \325  = (~\27  & \87 ) | (\27  & ~\87 ),
  \326  = ~\327 ,
  \327  = (~\26  & \86 ) | (\26  & ~\86 ),
  \328  = ~\329 ,
  \329  = (~\25  & \85 ) | (\25  & ~\85 ),
  \330  = ~\331 ,
  \331  = (~\24  & \84 ) | (\24  & ~\84 ),
  \332  = ~\333 ,
  \333  = (~\23  & \83 ) | (\23  & ~\83 ),
  \334  = ~\335 ,
  \335  = (~\22  & \82 ) | (\22  & ~\82 ),
  \336  = ~\337 ,
  \337  = (~\21  & \81 ) | (\21  & ~\81 ),
  \338  = ~\339 ,
  \339  = (~\20  & \80 ) | (\20  & ~\80 ),
  \340  = ~\341 ,
  \341  = (~\19  & \79 ) | (\19  & ~\79 ),
  \342  = ~\343 ,
  \343  = (~\18  & \78 ) | (\18  & ~\78 ),
  \344  = ~\345 ,
  \345  = (~\17  & \77 ) | (\17  & ~\77 ),
  \346  = ~\347 ,
  \347  = (~\16  & \76 ) | (\16  & ~\76 ),
  \348  = ~\349 ,
  \349  = (~\15  & \75 ) | (\15  & ~\75 ),
  \350  = ~\351 ,
  \351  = (~\14  & \74 ) | (\14  & ~\74 ),
  \352  = ~\353 ,
  \353  = (~\13  & \73 ) | (\13  & ~\73 ),
  \354  = ~\355 ,
  \355  = (~\12  & \72 ) | (\12  & ~\72 ),
  \356  = ~\357 ,
  \357  = (~\11  & \71 ) | (\11  & ~\71 ),
  \358  = ~\359 ,
  \359  = (~\10  & \70 ) | (\10  & ~\70 ),
  \360  = ~\361 ,
  \361  = (~\9  & \69 ) | (\9  & ~\69 ),
  \362  = ~\363 ,
  \363  = (~\8  & \68 ) | (\8  & ~\68 ),
  \364  = ~\365 ,
  \365  = (~\7  & \67 ) | (\7  & ~\67 ),
  \366  = ~\367 ,
  \367  = (~\6  & \66 ) | (\6  & ~\66 ),
  \368  = ~\369 ,
  \369  = (~\5  & \65 ) | (\5  & ~\65 ),
  \370  = ~\371 ,
  \371  = (~\4  & \64 ) | (\4  & ~\64 ),
  \372  = ~\373 ,
  \373  = ~\1037 ,
  \374  = 0,
  \375  = 0,
  \376  = 0,
  \377  = 0,
  \378  = 0,
  \379  = 0,
  \380  = 0,
  \381  = 0,
  \382  = 0,
  \383  = 0,
  \384  = 0,
  \385  = 0,
  \386  = 0,
  \387  = 0,
  \388  = 0,
  \389  = 0,
  \390  = 0,
  \391  = 0,
  \392  = 0,
  \393  = 0,
  \394  = 0,
  \395  = 0,
  \396  = 0,
  \397  = 0,
  \398  = 0,
  \399  = 0,
  \400  = 0,
  \401  = 0,
  \402  = 0,
  \403  = 0,
  \404  = 0,
  \405  = 0,
  \406  = 0,
  \407  = 0,
  \408  = 0,
  \409  = 0,
  \410  = 0,
  \411  = 0,
  \412  = 0,
  \413  = 0,
  \414  = 0,
  \415  = 0,
  \416  = 0,
  \417  = 0,
  \418  = 0,
  \419  = 0,
  \420  = 0,
  \421  = 0,
  \422  = 0,
  \423  = 0,
  \424  = 0,
  \425  = 0,
  \426  = 0,
  \427  = 0,
  \428  = 0,
  \429  = 0,
  \430  = 0,
  \431  = 0,
  \432  = 0,
  \433  = 0,
  \434  = \4 ,
  \435  = \5 ,
  \436  = \6 ,
  \437  = \7 ,
  \438  = \8 ,
  \439  = \9 ,
  \440  = \10 ,
  \441  = \11 ,
  \442  = \12 ,
  \443  = \13 ,
  \444  = \14 ,
  \445  = \15 ,
  \446  = \16 ,
  \447  = \17 ,
  \448  = \18 ,
  \449  = \19 ,
  \450  = \20 ,
  \451  = \21 ,
  \452  = \22 ,
  \453  = \23 ,
  \454  = \24 ,
  \455  = \25 ,
  \456  = \26 ,
  \457  = \27 ,
  \458  = \28 ,
  \459  = \29 ,
  \460  = \30 ,
  \461  = \31 ,
  \462  = \32 ,
  \463  = \33 ,
  \464  = \34 ,
  \465  = \35 ,
  \466  = \36 ,
  \467  = \37 ,
  \468  = \38 ,
  \469  = \39 ,
  \470  = \40 ,
  \471  = \41 ,
  \472  = \42 ,
  \473  = \43 ,
  \474  = \44 ,
  \475  = \45 ,
  \476  = \46 ,
  \477  = \47 ,
  \478  = \48 ,
  \479  = \49 ,
  \480  = \50 ,
  \481  = \51 ,
  \482  = \52 ,
  \483  = \53 ,
  \484  = \54 ,
  \485  = \55 ,
  \486  = \56 ,
  \487  = \57 ,
  \488  = \58 ,
  \489  = \59 ,
  \490  = \60 ,
  \491  = \61 ,
  \492  = \62 ,
  \493  = \63 ,
  \494  = 0,
  \495  = 0,
  \496  = 0,
  \497  = 0,
  \498  = 0,
  \499  = 0,
  \500  = 0,
  \501  = 0,
  \502  = 0,
  \503  = 0,
  \504  = 0,
  \505  = 0,
  \506  = 0,
  \507  = 0,
  \508  = 0,
  \509  = 0,
  \510  = 0,
  \511  = 0,
  \512  = 0,
  \513  = 0,
  \514  = 0,
  \515  = 0,
  \516  = 0,
  \517  = 0,
  \518  = 0,
  \519  = 0,
  \520  = 0,
  \521  = 0,
  \522  = 0,
  \523  = 0,
  \524  = 0,
  \525  = 0,
  \526  = 0,
  \527  = 0,
  \528  = 0,
  \529  = 0,
  \530  = 0,
  \531  = 0,
  \532  = 0,
  \533  = 0,
  \534  = 0,
  \535  = 0,
  \536  = 0,
  \537  = 0,
  \538  = 0,
  \539  = 0,
  \540  = 0,
  \541  = 0,
  \542  = 0,
  \543  = 0,
  \544  = 0,
  \545  = 0,
  \546  = 0,
  \547  = 0,
  \548  = 0,
  \549  = 0,
  \550  = 0,
  \551  = 0,
  \552  = 0,
  \553  = 0,
  \554  = 1,
  \555  = 1,
  \556  = 1,
  \557  = 1,
  \558  = 1,
  \559  = 1,
  \560  = 1,
  \561  = 1,
  \562  = 1,
  \563  = 1,
  \564  = 1,
  \565  = 1,
  \566  = 1,
  \567  = 1,
  \568  = 1,
  \569  = 1,
  \570  = 1,
  \571  = 1,
  \572  = 1,
  \573  = 1,
  \574  = 1,
  \575  = 1,
  \576  = 1,
  \577  = 1,
  \578  = 1,
  \579  = 1,
  \580  = 1,
  \581  = 1,
  \582  = 1,
  \583  = 1,
  \584  = \4 ,
  \585  = \5 ,
  \586  = \6 ,
  \587  = \7 ,
  \588  = \8 ,
  \589  = \9 ,
  \590  = \10 ,
  \591  = \11 ,
  \592  = \12 ,
  \593  = \13 ,
  \594  = \14 ,
  \595  = \15 ,
  \596  = \16 ,
  \597  = \17 ,
  \598  = \18 ,
  \599  = \19 ,
  \600  = \20 ,
  \601  = \21 ,
  \602  = \22 ,
  \603  = \23 ,
  \604  = \24 ,
  \605  = \25 ,
  \606  = \26 ,
  \607  = \27 ,
  \608  = \28 ,
  \609  = \29 ,
  \610  = \30 ,
  \611  = \31 ,
  \612  = \32 ,
  \613  = \33 ,
  \614  = 0,
  \615  = 0,
  \616  = 0,
  \617  = 0,
  \618  = 0,
  \619  = 0,
  \620  = 0,
  \621  = 0,
  \622  = 0,
  \623  = 0,
  \624  = 0,
  \625  = 0,
  \626  = 0,
  \627  = 0,
  \628  = 0,
  \629  = 0,
  \630  = 0,
  \631  = 0,
  \632  = 0,
  \633  = 0,
  \634  = 0,
  \635  = 0,
  \636  = 0,
  \637  = 0,
  \638  = 0,
  \639  = 0,
  \640  = 0,
  \641  = 0,
  \642  = 0,
  \643  = 0,
  \644  = 0,
  \645  = 0,
  \646  = 0,
  \647  = 0,
  \648  = 0,
  \649  = 0;
always begin
  \34  = \[120] ;
  \35  = \[121] ;
  \36  = \[122] ;
  \37  = \[123] ;
  \38  = \[124] ;
  \39  = \[125] ;
  \40  = \[126] ;
  \41  = \[127] ;
  \42  = \[128] ;
  \43  = \[129] ;
  \44  = \[130] ;
  \45  = \[131] ;
  \46  = \[132] ;
  \47  = \[133] ;
  \48  = \[134] ;
  \49  = \[135] ;
  \50  = \[136] ;
  \51  = \[137] ;
  \52  = \[138] ;
  \53  = \[139] ;
  \54  = \[140] ;
  \55  = \[141] ;
  \56  = \[142] ;
  \57  = \[143] ;
  \58  = \[144] ;
  \59  = \[145] ;
  \60  = \[146] ;
  \61  = \[147] ;
  \62  = \[148] ;
  \63  = \[149] ;
  \64  = \[150] ;
  \65  = \[151] ;
  \66  = \[152] ;
  \67  = \[153] ;
  \68  = \[154] ;
  \69  = \[155] ;
  \70  = \[156] ;
  \71  = \[157] ;
  \72  = \[158] ;
  \73  = \[159] ;
  \74  = \[160] ;
  \75  = \[161] ;
  \76  = \[162] ;
  \77  = \[163] ;
  \78  = \[164] ;
  \79  = \[165] ;
  \80  = \[166] ;
  \81  = \[167] ;
  \82  = \[168] ;
  \83  = \[169] ;
  \84  = \[170] ;
  \85  = \[171] ;
  \86  = \[172] ;
  \87  = \[173] ;
  \88  = \[174] ;
  \89  = \[175] ;
  \90  = \[176] ;
  \91  = \[177] ;
  \92  = \[178] ;
  \93  = \[179] ;
  \94  = \[180] ;
  \95  = \[181] ;
  \96  = \[182] ;
  \97  = \[183] ;
  \98  = \[184] ;
  \99  = \[185] ;
  \100  = \[186] ;
  \101  = \[187] ;
  \102  = \[188] ;
  \103  = \[189] ;
  \104  = \[190] ;
  \105  = \[191] ;
  \106  = \[192] ;
  \107  = \[193] ;
  \108  = \[194] ;
  \109  = \[195] ;
  \110  = \[196] ;
  \111  = \[197] ;
  \112  = \[198] ;
  \113  = \[199] ;
  \114  = \[200] ;
  \115  = \[201] ;
  \116  = \[202] ;
  \117  = \[203] ;
  \118  = \[204] ;
  \119  = \[205] ;
  \120  = \[206] ;
  \121  = \[207] ;
  \122  = \[208] ;
  \123  = \[209] ;
end
initial begin
  \64  = 1;
  \65  = 1;
  \66  = 1;
  \67  = 1;
  \68  = 1;
  \69  = 1;
  \70  = 1;
  \71  = 1;
  \72  = 1;
  \73  = 1;
  \74  = 1;
  \75  = 1;
  \76  = 1;
  \77  = 1;
  \78  = 1;
  \79  = 1;
  \80  = 1;
  \81  = 1;
  \82  = 1;
  \83  = 1;
  \84  = 1;
  \85  = 1;
  \86  = 1;
  \87  = 1;
  \88  = 1;
  \89  = 1;
  \90  = 1;
  \91  = 1;
  \92  = 1;
  \93  = 1;
  \94  = 0;
  \95  = 0;
  \96  = 0;
  \97  = 0;
  \98  = 0;
  \99  = 0;
  \100  = 0;
  \101  = 0;
  \102  = 0;
  \103  = 0;
  \104  = 0;
  \105  = 0;
  \106  = 0;
  \107  = 0;
  \108  = 0;
  \109  = 0;
  \110  = 0;
  \111  = 0;
  \112  = 0;
  \113  = 0;
  \114  = 0;
  \115  = 0;
  \116  = 0;
  \117  = 0;
  \118  = 0;
  \119  = 0;
  \120  = 0;
  \121  = 0;
  \122  = 0;
  \123  = 0;
end
endmodule

