module s382 (
  CK,
  CLR,
  FM,
  TEST,
  YLW2,
  RED2,
  GRN1,
  RED1,
  YLW1,
  GRN2
);
  input CK;
  wire CK;
  input CLR;
  wire CLR;
  input FM;
  wire FM;
  input TEST;
  wire TEST;
  output YLW2;
  wire YLW2;
  output RED2;
  wire RED2;
  output GRN1;
  wire GRN1;
  output RED1;
  wire RED1;
  output YLW1;
  wire YLW1;
  output GRN2;
  wire GRN2;
  wire __0__;
  wire __1__;
  wire __2__;
  wire __3__;
  wire __4__;
  wire __5__;
  wire __6__;
  wire __7__;
  wire __8__;
  wire __9__;
  wire __10__;
  wire __11__;
  wire __12__;
  wire __13__;
  wire __14__;
  wire __15__;
  wire __16__;
  wire __17__;
  wire __18__;
  wire __19__;
  wire __20__;
  wire __21__;
  wire __22__;
  wire __25__;
  wire __26__;
  wire __27__;
  wire __28__;
  wire __29__;
  wire __30__;
  wire __31__;
  wire __32__;
  wire __33__;
  wire __34__;
  wire __35__;
  wire __36__;
  wire __37__;
  wire __38__;
  wire __39__;
  wire __40__;
  wire __41__;
  wire __42__;
  wire __43__;
  wire __44__;
  wire __45__;
  wire __46__;
  wire __47__;
  wire __48__;
  wire __49__;
  wire __50__;
  wire __51__;
  wire __52__;
  wire __53__;
  INV __54__ (
    .I(__6__),
    .O(__0__)
  );
  INV __55__ (
    .I(__5__),
    .O(__1__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __56__ (
    .D(__28__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__2__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __57__ (
    .D(__34__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__3__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __58__ (
    .D(__35__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__4__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __59__ (
    .D(__51__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__5__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __60__ (
    .D(__53__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__6__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __61__ (
    .D(__41__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__7__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __62__ (
    .D(__38__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__8__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __63__ (
    .D(__45__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__9__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __64__ (
    .D(__33__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__10__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __65__ (
    .D(__46__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__11__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __66__ (
    .D(__40__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__12__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __67__ (
    .D(__30__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__13__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __68__ (
    .D(__43__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__14__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __69__ (
    .D(__36__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__15__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __70__ (
    .D(__27__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__16__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __71__ (
    .D(__49__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__17__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __72__ (
    .D(__37__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__18__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __73__ (
    .D(__25__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__19__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __74__ (
    .D(__42__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__20__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __75__ (
    .D(__48__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__21__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __76__ (
    .D(__47__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__22__)
  );
  LUT5 #(
    .INIT(32'h10000004)
  ) __79__ (
    .I4(__22__),
    .I3(__21__),
    .I2(__20__),
    .I1(__19__),
    .I0(CLR),
    .O(__25__)
  );
  LUT5 #(
    .INIT(32'h000001ff)
  ) __80__ (
    .I4(__3__),
    .I3(__19__),
    .I2(__22__),
    .I1(__21__),
    .I0(__20__),
    .O(__26__)
  );
  LUT6 #(
    .INIT(64'h0000aabf00000040)
  ) __81__ (
    .I5(__16__),
    .I4(CLR),
    .I3(__15__),
    .I2(__17__),
    .I1(__18__),
    .I0(__26__),
    .O(__27__)
  );
  LUT5 #(
    .INIT(32'h00000020)
  ) __82__ (
    .I4(CLR),
    .I3(__12__),
    .I2(__14__),
    .I1(__10__),
    .I0(__13__),
    .O(__28__)
  );
  LUT4 #(
    .INIT(16'hfe00)
  ) __83__ (
    .I3(__15__),
    .I2(__16__),
    .I1(__17__),
    .I0(__18__),
    .O(__29__)
  );
  LUT6 #(
    .INIT(64'h00000000bb04bf00)
  ) __84__ (
    .I5(CLR),
    .I4(__14__),
    .I3(__13__),
    .I2(__11__),
    .I1(__29__),
    .I0(__26__),
    .O(__30__)
  );
  LUT2 #(
    .INIT(4'h1)
  ) __85__ (
    .I1(__14__),
    .I0(__13__),
    .O(__31__)
  );
  LUT4 #(
    .INIT(16'h0100)
  ) __86__ (
    .I3(__14__),
    .I2(__13__),
    .I1(__11__),
    .I0(__4__),
    .O(__32__)
  );
  LUT6 #(
    .INIT(64'h000000008f88ff00)
  ) __87__ (
    .I5(CLR),
    .I4(__12__),
    .I3(__10__),
    .I2(__32__),
    .I1(__4__),
    .I0(__31__),
    .O(__33__)
  );
  LUT3 #(
    .INIT(8'h14)
  ) __88__ (
    .I2(__3__),
    .I1(TEST),
    .I0(CLR),
    .O(__34__)
  );
  LUT3 #(
    .INIT(8'h14)
  ) __89__ (
    .I2(__4__),
    .I1(FM),
    .I0(CLR),
    .O(__35__)
  );
  LUT6 #(
    .INIT(64'h0000aaab00004000)
  ) __90__ (
    .I5(__15__),
    .I4(CLR),
    .I3(__16__),
    .I2(__17__),
    .I1(__18__),
    .I0(__26__),
    .O(__36__)
  );
  LUT6 #(
    .INIT(64'h00000000a1a1a1a5)
  ) __91__ (
    .I5(CLR),
    .I4(__16__),
    .I3(__17__),
    .I2(__18__),
    .I1(__15__),
    .I0(__26__),
    .O(__37__)
  );
  LUT6 #(
    .INIT(64'hffffffff00000035)
  ) __92__ (
    .I5(CLR),
    .I4(__12__),
    .I3(__10__),
    .I2(__14__),
    .I1(__13__),
    .I0(__11__),
    .O(__38__)
  );
  LUT5 #(
    .INIT(32'h0000fe00)
  ) __93__ (
    .I4(__26__),
    .I3(__15__),
    .I2(__16__),
    .I1(__17__),
    .I0(__18__),
    .O(__39__)
  );
  LUT6 #(
    .INIT(64'h0000557f00000080)
  ) __94__ (
    .I5(__12__),
    .I4(CLR),
    .I3(__11__),
    .I2(__14__),
    .I1(__13__),
    .I0(__39__),
    .O(__40__)
  );
  LUT6 #(
    .INIT(64'hff00ff00ff00ff4f)
  ) __95__ (
    .I5(__12__),
    .I4(__10__),
    .I3(CLR),
    .I2(__11__),
    .I1(__14__),
    .I0(__13__),
    .O(__41__)
  );
  LUT5 #(
    .INIT(32'h00070008)
  ) __96__ (
    .I4(__20__),
    .I3(CLR),
    .I2(__19__),
    .I1(__22__),
    .I0(__21__),
    .O(__42__)
  );
  LUT6 #(
    .INIT(64'h0000001f00ff0000)
  ) __97__ (
    .I5(__39__),
    .I4(__14__),
    .I3(CLR),
    .I2(__11__),
    .I1(__12__),
    .I0(__13__),
    .O(__43__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __98__ (
    .I1(__12__),
    .I0(CLR),
    .O(__44__)
  );
  LUT6 #(
    .INIT(64'h005510fd00000000)
  ) __99__ (
    .I5(__44__),
    .I4(__11__),
    .I3(__10__),
    .I2(__14__),
    .I1(__13__),
    .I0(__4__),
    .O(__45__)
  );
  LUT6 #(
    .INIT(64'h0000555700008000)
  ) __100__ (
    .I5(__11__),
    .I4(CLR),
    .I3(__12__),
    .I2(__14__),
    .I1(__13__),
    .I0(__39__),
    .O(__46__)
  );
  LUT5 #(
    .INIT(32'h0000001f)
  ) __101__ (
    .I4(CLR),
    .I3(__22__),
    .I2(__19__),
    .I1(__21__),
    .I0(__20__),
    .O(__47__)
  );
  LUT4 #(
    .INIT(16'h0110)
  ) __102__ (
    .I3(__22__),
    .I2(__21__),
    .I1(CLR),
    .I0(__19__),
    .O(__48__)
  );
  LUT6 #(
    .INIT(64'h00000000ab10ab10)
  ) __103__ (
    .I5(CLR),
    .I4(__16__),
    .I3(__17__),
    .I2(__18__),
    .I1(__15__),
    .I0(__26__),
    .O(__49__)
  );
  LUT6 #(
    .INIT(64'h000000000002000c)
  ) __104__ (
    .I5(CLR),
    .I4(__12__),
    .I3(__14__),
    .I2(__13__),
    .I1(__11__),
    .I0(__4__),
    .O(__50__)
  );
  LUT5 #(
    .INIT(32'hd5d5cfd5)
  ) __105__ (
    .I4(CLR),
    .I3(__10__),
    .I2(__33__),
    .I1(__16__),
    .I0(__50__),
    .O(__51__)
  );
  LUT3 #(
    .INIT(8'h04)
  ) __106__ (
    .I2(CLR),
    .I1(__11__),
    .I0(__14__),
    .O(__52__)
  );
  LUT6 #(
    .INIT(64'hcfc5cfc5c0c0cfc5)
  ) __107__ (
    .I5(CLR),
    .I4(__12__),
    .I3(__13__),
    .I2(__33__),
    .I1(__16__),
    .I0(__52__),
    .O(__53__)
  );
  assign YLW2 = __2__;
  assign RED2 = __0__;
  assign GRN1 = __9__;
  assign RED1 = __7__;
  assign YLW1 = __1__;
  assign GRN2 = __8__;
endmodule
