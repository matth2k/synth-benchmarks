module s35932 (
  CK,
  DATA_0_0,
  DATA_0_1,
  DATA_0_10,
  DATA_0_11,
  DATA_0_12,
  DATA_0_13,
  DATA_0_14,
  DATA_0_15,
  DATA_0_16,
  DATA_0_17,
  DATA_0_18,
  DATA_0_19,
  DATA_0_2,
  DATA_0_20,
  DATA_0_21,
  DATA_0_22,
  DATA_0_23,
  DATA_0_24,
  DATA_0_25,
  DATA_0_26,
  DATA_0_27,
  DATA_0_28,
  DATA_0_29,
  DATA_0_3,
  DATA_0_30,
  DATA_0_31,
  DATA_0_4,
  DATA_0_5,
  DATA_0_6,
  DATA_0_7,
  DATA_0_8,
  DATA_0_9,
  RESET,
  TM0,
  TM1,
  CRC_OUT_9_24,
  CRC_OUT_5_23,
  CRC_OUT_2_14,
  CRC_OUT_7_5,
  CRC_OUT_4_23,
  CRC_OUT_1_28,
  CRC_OUT_6_13,
  CRC_OUT_1_19,
  CRC_OUT_9_31,
  CRC_OUT_4_14,
  CRC_OUT_5_3,
  CRC_OUT_2_15,
  CRC_OUT_7_15,
  CRC_OUT_2_3,
  CRC_OUT_3_12,
  CRC_OUT_1_6,
  CRC_OUT_6_21,
  CRC_OUT_9_25,
  CRC_OUT_2_25,
  DATA_9_15,
  CRC_OUT_6_26,
  DATA_9_4,
  CRC_OUT_6_3,
  CRC_OUT_2_29,
  CRC_OUT_3_10,
  CRC_OUT_5_6,
  CRC_OUT_2_20,
  CRC_OUT_3_27,
  CRC_OUT_6_30,
  CRC_OUT_2_5,
  CRC_OUT_1_20,
  CRC_OUT_6_11,
  CRC_OUT_7_29,
  CRC_OUT_9_19,
  CRC_OUT_1_16,
  CRC_OUT_5_1,
  CRC_OUT_3_8,
  CRC_OUT_7_3,
  CRC_OUT_2_8,
  DATA_9_20,
  CRC_OUT_9_11,
  CRC_OUT_7_26,
  CRC_OUT_1_7,
  CRC_OUT_2_17,
  CRC_OUT_2_6,
  CRC_OUT_4_11,
  CRC_OUT_9_4,
  CRC_OUT_9_6,
  CRC_OUT_8_3,
  DATA_9_21,
  CRC_OUT_7_19,
  CRC_OUT_7_22,
  DATA_9_17,
  CRC_OUT_9_22,
  CRC_OUT_4_31,
  CRC_OUT_2_12,
  CRC_OUT_9_21,
  CRC_OUT_8_29,
  CRC_OUT_9_7,
  CRC_OUT_9_5,
  CRC_OUT_6_7,
  DATA_9_11,
  CRC_OUT_3_9,
  CRC_OUT_4_18,
  CRC_OUT_7_20,
  CRC_OUT_1_11,
  CRC_OUT_3_15,
  CRC_OUT_8_31,
  CRC_OUT_5_13,
  CRC_OUT_1_31,
  CRC_OUT_6_28,
  CRC_OUT_5_19,
  CRC_OUT_3_3,
  CRC_OUT_6_0,
  DATA_9_8,
  CRC_OUT_9_29,
  CRC_OUT_8_21,
  DATA_9_0,
  CRC_OUT_9_26,
  CRC_OUT_1_4,
  CRC_OUT_1_22,
  CRC_OUT_4_24,
  CRC_OUT_6_6,
  CRC_OUT_4_13,
  CRC_OUT_3_16,
  CRC_OUT_4_10,
  CRC_OUT_5_25,
  CRC_OUT_7_2,
  CRC_OUT_5_12,
  CRC_OUT_8_10,
  CRC_OUT_4_0,
  CRC_OUT_6_16,
  CRC_OUT_7_4,
  CRC_OUT_5_14,
  CRC_OUT_3_24,
  CRC_OUT_6_18,
  CRC_OUT_9_14,
  CRC_OUT_3_7,
  CRC_OUT_6_24,
  CRC_OUT_5_5,
  CRC_OUT_6_19,
  CRC_OUT_3_11,
  CRC_OUT_8_11,
  CRC_OUT_6_20,
  CRC_OUT_5_24,
  CRC_OUT_4_2,
  CRC_OUT_3_6,
  CRC_OUT_4_27,
  CRC_OUT_6_9,
  CRC_OUT_2_2,
  CRC_OUT_5_4,
  CRC_OUT_7_27,
  CRC_OUT_2_26,
  CRC_OUT_5_7,
  CRC_OUT_2_27,
  CRC_OUT_5_20,
  CRC_OUT_4_17,
  CRC_OUT_8_6,
  CRC_OUT_2_11,
  CRC_OUT_4_3,
  CRC_OUT_8_26,
  CRC_OUT_1_5,
  CRC_OUT_4_4,
  CRC_OUT_5_0,
  CRC_OUT_4_22,
  CRC_OUT_9_27,
  CRC_OUT_9_8,
  DATA_9_13,
  DATA_9_7,
  CRC_OUT_3_14,
  CRC_OUT_3_2,
  CRC_OUT_3_5,
  CRC_OUT_3_20,
  CRC_OUT_8_2,
  CRC_OUT_7_17,
  CRC_OUT_2_24,
  CRC_OUT_8_25,
  DATA_9_1,
  CRC_OUT_2_16,
  CRC_OUT_5_29,
  DATA_9_29,
  CRC_OUT_2_22,
  CRC_OUT_4_19,
  DATA_9_27,
  CRC_OUT_1_15,
  CRC_OUT_2_4,
  CRC_OUT_9_28,
  CRC_OUT_4_5,
  CRC_OUT_2_7,
  DATA_9_30,
  CRC_OUT_5_30,
  CRC_OUT_2_23,
  CRC_OUT_6_31,
  CRC_OUT_1_17,
  CRC_OUT_4_7,
  CRC_OUT_4_25,
  CRC_OUT_6_14,
  CRC_OUT_3_18,
  CRC_OUT_5_26,
  CRC_OUT_5_28,
  CRC_OUT_1_27,
  CRC_OUT_7_12,
  CRC_OUT_3_28,
  CRC_OUT_9_16,
  CRC_OUT_4_12,
  CRC_OUT_7_7,
  CRC_OUT_4_15,
  CRC_OUT_6_10,
  DATA_9_25,
  CRC_OUT_7_8,
  CRC_OUT_9_30,
  CRC_OUT_8_1,
  CRC_OUT_8_16,
  CRC_OUT_3_31,
  CRC_OUT_1_3,
  CRC_OUT_2_30,
  CRC_OUT_4_8,
  CRC_OUT_1_23,
  CRC_OUT_8_30,
  CRC_OUT_6_1,
  CRC_OUT_8_7,
  CRC_OUT_8_8,
  CRC_OUT_9_13,
  CRC_OUT_5_11,
  CRC_OUT_1_0,
  CRC_OUT_3_29,
  CRC_OUT_7_9,
  CRC_OUT_5_8,
  CRC_OUT_5_21,
  CRC_OUT_9_2,
  CRC_OUT_2_0,
  DATA_9_26,
  CRC_OUT_3_17,
  CRC_OUT_8_15,
  DATA_9_2,
  CRC_OUT_2_28,
  DATA_9_14,
  CRC_OUT_9_17,
  CRC_OUT_9_3,
  DATA_9_9,
  CRC_OUT_8_17,
  DATA_9_19,
  DATA_9_10,
  CRC_OUT_7_13,
  CRC_OUT_7_23,
  CRC_OUT_2_1,
  CRC_OUT_1_26,
  CRC_OUT_9_9,
  CRC_OUT_8_14,
  CRC_OUT_1_14,
  CRC_OUT_7_16,
  CRC_OUT_3_23,
  CRC_OUT_8_13,
  CRC_OUT_9_23,
  CRC_OUT_8_19,
  DATA_9_23,
  CRC_OUT_8_28,
  CRC_OUT_9_18,
  CRC_OUT_1_21,
  CRC_OUT_4_1,
  CRC_OUT_1_24,
  CRC_OUT_2_21,
  CRC_OUT_4_26,
  CRC_OUT_6_2,
  CRC_OUT_7_25,
  CRC_OUT_3_25,
  CRC_OUT_9_12,
  CRC_OUT_9_15,
  DATA_9_22,
  CRC_OUT_1_1,
  DATA_9_5,
  CRC_OUT_8_0,
  DATA_9_31,
  CRC_OUT_7_21,
  DATA_9_16,
  CRC_OUT_2_13,
  CRC_OUT_9_10,
  DATA_9_28,
  CRC_OUT_8_4,
  CRC_OUT_4_29,
  CRC_OUT_6_8,
  CRC_OUT_3_13,
  CRC_OUT_3_30,
  CRC_OUT_1_30,
  CRC_OUT_8_5,
  CRC_OUT_6_15,
  CRC_OUT_6_5,
  CRC_OUT_1_10,
  CRC_OUT_7_18,
  CRC_OUT_4_9,
  CRC_OUT_1_13,
  CRC_OUT_8_27,
  CRC_OUT_5_2,
  CRC_OUT_8_12,
  CRC_OUT_8_22,
  CRC_OUT_7_11,
  CRC_OUT_7_10,
  CRC_OUT_6_25,
  CRC_OUT_6_23,
  CRC_OUT_1_9,
  CRC_OUT_7_0,
  CRC_OUT_7_1,
  CRC_OUT_4_21,
  CRC_OUT_9_0,
  CRC_OUT_1_2,
  CRC_OUT_6_17,
  CRC_OUT_5_10,
  CRC_OUT_8_9,
  CRC_OUT_7_24,
  CRC_OUT_5_22,
  CRC_OUT_7_14,
  DATA_9_18,
  CRC_OUT_7_28,
  CRC_OUT_3_22,
  CRC_OUT_6_29,
  CRC_OUT_8_20,
  CRC_OUT_6_22,
  CRC_OUT_5_17,
  CRC_OUT_3_1,
  CRC_OUT_3_19,
  CRC_OUT_5_9,
  CRC_OUT_3_4,
  CRC_OUT_1_18,
  CRC_OUT_5_16,
  CRC_OUT_6_4,
  CRC_OUT_8_24,
  CRC_OUT_2_10,
  DATA_9_24,
  CRC_OUT_8_23,
  CRC_OUT_8_18,
  CRC_OUT_1_8,
  CRC_OUT_2_31,
  CRC_OUT_2_19,
  CRC_OUT_4_16,
  CRC_OUT_7_31,
  CRC_OUT_2_18,
  CRC_OUT_4_6,
  CRC_OUT_2_9,
  CRC_OUT_5_31,
  CRC_OUT_5_18,
  CRC_OUT_6_27,
  CRC_OUT_3_21,
  CRC_OUT_1_25,
  CRC_OUT_4_30,
  DATA_9_3,
  CRC_OUT_1_12,
  CRC_OUT_7_6,
  CRC_OUT_9_1,
  CRC_OUT_5_15,
  CRC_OUT_5_27,
  CRC_OUT_7_30,
  CRC_OUT_3_26,
  CRC_OUT_3_0,
  CRC_OUT_1_29,
  CRC_OUT_9_20,
  DATA_9_12,
  CRC_OUT_6_12,
  DATA_9_6,
  CRC_OUT_4_20,
  CRC_OUT_4_28
);
  input CK;
  wire CK;
  input DATA_0_0;
  wire DATA_0_0;
  input DATA_0_1;
  wire DATA_0_1;
  input DATA_0_10;
  wire DATA_0_10;
  input DATA_0_11;
  wire DATA_0_11;
  input DATA_0_12;
  wire DATA_0_12;
  input DATA_0_13;
  wire DATA_0_13;
  input DATA_0_14;
  wire DATA_0_14;
  input DATA_0_15;
  wire DATA_0_15;
  input DATA_0_16;
  wire DATA_0_16;
  input DATA_0_17;
  wire DATA_0_17;
  input DATA_0_18;
  wire DATA_0_18;
  input DATA_0_19;
  wire DATA_0_19;
  input DATA_0_2;
  wire DATA_0_2;
  input DATA_0_20;
  wire DATA_0_20;
  input DATA_0_21;
  wire DATA_0_21;
  input DATA_0_22;
  wire DATA_0_22;
  input DATA_0_23;
  wire DATA_0_23;
  input DATA_0_24;
  wire DATA_0_24;
  input DATA_0_25;
  wire DATA_0_25;
  input DATA_0_26;
  wire DATA_0_26;
  input DATA_0_27;
  wire DATA_0_27;
  input DATA_0_28;
  wire DATA_0_28;
  input DATA_0_29;
  wire DATA_0_29;
  input DATA_0_3;
  wire DATA_0_3;
  input DATA_0_30;
  wire DATA_0_30;
  input DATA_0_31;
  wire DATA_0_31;
  input DATA_0_4;
  wire DATA_0_4;
  input DATA_0_5;
  wire DATA_0_5;
  input DATA_0_6;
  wire DATA_0_6;
  input DATA_0_7;
  wire DATA_0_7;
  input DATA_0_8;
  wire DATA_0_8;
  input DATA_0_9;
  wire DATA_0_9;
  input RESET;
  wire RESET;
  input TM0;
  wire TM0;
  input TM1;
  wire TM1;
  output CRC_OUT_9_24;
  wire CRC_OUT_9_24;
  output CRC_OUT_5_23;
  wire CRC_OUT_5_23;
  output CRC_OUT_2_14;
  wire CRC_OUT_2_14;
  output CRC_OUT_7_5;
  wire CRC_OUT_7_5;
  output CRC_OUT_4_23;
  wire CRC_OUT_4_23;
  output CRC_OUT_1_28;
  wire CRC_OUT_1_28;
  output CRC_OUT_6_13;
  wire CRC_OUT_6_13;
  output CRC_OUT_1_19;
  wire CRC_OUT_1_19;
  output CRC_OUT_9_31;
  wire CRC_OUT_9_31;
  output CRC_OUT_4_14;
  wire CRC_OUT_4_14;
  output CRC_OUT_5_3;
  wire CRC_OUT_5_3;
  output CRC_OUT_2_15;
  wire CRC_OUT_2_15;
  output CRC_OUT_7_15;
  wire CRC_OUT_7_15;
  output CRC_OUT_2_3;
  wire CRC_OUT_2_3;
  output CRC_OUT_3_12;
  wire CRC_OUT_3_12;
  output CRC_OUT_1_6;
  wire CRC_OUT_1_6;
  output CRC_OUT_6_21;
  wire CRC_OUT_6_21;
  output CRC_OUT_9_25;
  wire CRC_OUT_9_25;
  output CRC_OUT_2_25;
  wire CRC_OUT_2_25;
  output DATA_9_15;
  wire DATA_9_15;
  output CRC_OUT_6_26;
  wire CRC_OUT_6_26;
  output DATA_9_4;
  wire DATA_9_4;
  output CRC_OUT_6_3;
  wire CRC_OUT_6_3;
  output CRC_OUT_2_29;
  wire CRC_OUT_2_29;
  output CRC_OUT_3_10;
  wire CRC_OUT_3_10;
  output CRC_OUT_5_6;
  wire CRC_OUT_5_6;
  output CRC_OUT_2_20;
  wire CRC_OUT_2_20;
  output CRC_OUT_3_27;
  wire CRC_OUT_3_27;
  output CRC_OUT_6_30;
  wire CRC_OUT_6_30;
  output CRC_OUT_2_5;
  wire CRC_OUT_2_5;
  output CRC_OUT_1_20;
  wire CRC_OUT_1_20;
  output CRC_OUT_6_11;
  wire CRC_OUT_6_11;
  output CRC_OUT_7_29;
  wire CRC_OUT_7_29;
  output CRC_OUT_9_19;
  wire CRC_OUT_9_19;
  output CRC_OUT_1_16;
  wire CRC_OUT_1_16;
  output CRC_OUT_5_1;
  wire CRC_OUT_5_1;
  output CRC_OUT_3_8;
  wire CRC_OUT_3_8;
  output CRC_OUT_7_3;
  wire CRC_OUT_7_3;
  output CRC_OUT_2_8;
  wire CRC_OUT_2_8;
  output DATA_9_20;
  wire DATA_9_20;
  output CRC_OUT_9_11;
  wire CRC_OUT_9_11;
  output CRC_OUT_7_26;
  wire CRC_OUT_7_26;
  output CRC_OUT_1_7;
  wire CRC_OUT_1_7;
  output CRC_OUT_2_17;
  wire CRC_OUT_2_17;
  output CRC_OUT_2_6;
  wire CRC_OUT_2_6;
  output CRC_OUT_4_11;
  wire CRC_OUT_4_11;
  output CRC_OUT_9_4;
  wire CRC_OUT_9_4;
  output CRC_OUT_9_6;
  wire CRC_OUT_9_6;
  output CRC_OUT_8_3;
  wire CRC_OUT_8_3;
  output DATA_9_21;
  wire DATA_9_21;
  output CRC_OUT_7_19;
  wire CRC_OUT_7_19;
  output CRC_OUT_7_22;
  wire CRC_OUT_7_22;
  output DATA_9_17;
  wire DATA_9_17;
  output CRC_OUT_9_22;
  wire CRC_OUT_9_22;
  output CRC_OUT_4_31;
  wire CRC_OUT_4_31;
  output CRC_OUT_2_12;
  wire CRC_OUT_2_12;
  output CRC_OUT_9_21;
  wire CRC_OUT_9_21;
  output CRC_OUT_8_29;
  wire CRC_OUT_8_29;
  output CRC_OUT_9_7;
  wire CRC_OUT_9_7;
  output CRC_OUT_9_5;
  wire CRC_OUT_9_5;
  output CRC_OUT_6_7;
  wire CRC_OUT_6_7;
  output DATA_9_11;
  wire DATA_9_11;
  output CRC_OUT_3_9;
  wire CRC_OUT_3_9;
  output CRC_OUT_4_18;
  wire CRC_OUT_4_18;
  output CRC_OUT_7_20;
  wire CRC_OUT_7_20;
  output CRC_OUT_1_11;
  wire CRC_OUT_1_11;
  output CRC_OUT_3_15;
  wire CRC_OUT_3_15;
  output CRC_OUT_8_31;
  wire CRC_OUT_8_31;
  output CRC_OUT_5_13;
  wire CRC_OUT_5_13;
  output CRC_OUT_1_31;
  wire CRC_OUT_1_31;
  output CRC_OUT_6_28;
  wire CRC_OUT_6_28;
  output CRC_OUT_5_19;
  wire CRC_OUT_5_19;
  output CRC_OUT_3_3;
  wire CRC_OUT_3_3;
  output CRC_OUT_6_0;
  wire CRC_OUT_6_0;
  output DATA_9_8;
  wire DATA_9_8;
  output CRC_OUT_9_29;
  wire CRC_OUT_9_29;
  output CRC_OUT_8_21;
  wire CRC_OUT_8_21;
  output DATA_9_0;
  wire DATA_9_0;
  output CRC_OUT_9_26;
  wire CRC_OUT_9_26;
  output CRC_OUT_1_4;
  wire CRC_OUT_1_4;
  output CRC_OUT_1_22;
  wire CRC_OUT_1_22;
  output CRC_OUT_4_24;
  wire CRC_OUT_4_24;
  output CRC_OUT_6_6;
  wire CRC_OUT_6_6;
  output CRC_OUT_4_13;
  wire CRC_OUT_4_13;
  output CRC_OUT_3_16;
  wire CRC_OUT_3_16;
  output CRC_OUT_4_10;
  wire CRC_OUT_4_10;
  output CRC_OUT_5_25;
  wire CRC_OUT_5_25;
  output CRC_OUT_7_2;
  wire CRC_OUT_7_2;
  output CRC_OUT_5_12;
  wire CRC_OUT_5_12;
  output CRC_OUT_8_10;
  wire CRC_OUT_8_10;
  output CRC_OUT_4_0;
  wire CRC_OUT_4_0;
  output CRC_OUT_6_16;
  wire CRC_OUT_6_16;
  output CRC_OUT_7_4;
  wire CRC_OUT_7_4;
  output CRC_OUT_5_14;
  wire CRC_OUT_5_14;
  output CRC_OUT_3_24;
  wire CRC_OUT_3_24;
  output CRC_OUT_6_18;
  wire CRC_OUT_6_18;
  output CRC_OUT_9_14;
  wire CRC_OUT_9_14;
  output CRC_OUT_3_7;
  wire CRC_OUT_3_7;
  output CRC_OUT_6_24;
  wire CRC_OUT_6_24;
  output CRC_OUT_5_5;
  wire CRC_OUT_5_5;
  output CRC_OUT_6_19;
  wire CRC_OUT_6_19;
  output CRC_OUT_3_11;
  wire CRC_OUT_3_11;
  output CRC_OUT_8_11;
  wire CRC_OUT_8_11;
  output CRC_OUT_6_20;
  wire CRC_OUT_6_20;
  output CRC_OUT_5_24;
  wire CRC_OUT_5_24;
  output CRC_OUT_4_2;
  wire CRC_OUT_4_2;
  output CRC_OUT_3_6;
  wire CRC_OUT_3_6;
  output CRC_OUT_4_27;
  wire CRC_OUT_4_27;
  output CRC_OUT_6_9;
  wire CRC_OUT_6_9;
  output CRC_OUT_2_2;
  wire CRC_OUT_2_2;
  output CRC_OUT_5_4;
  wire CRC_OUT_5_4;
  output CRC_OUT_7_27;
  wire CRC_OUT_7_27;
  output CRC_OUT_2_26;
  wire CRC_OUT_2_26;
  output CRC_OUT_5_7;
  wire CRC_OUT_5_7;
  output CRC_OUT_2_27;
  wire CRC_OUT_2_27;
  output CRC_OUT_5_20;
  wire CRC_OUT_5_20;
  output CRC_OUT_4_17;
  wire CRC_OUT_4_17;
  output CRC_OUT_8_6;
  wire CRC_OUT_8_6;
  output CRC_OUT_2_11;
  wire CRC_OUT_2_11;
  output CRC_OUT_4_3;
  wire CRC_OUT_4_3;
  output CRC_OUT_8_26;
  wire CRC_OUT_8_26;
  output CRC_OUT_1_5;
  wire CRC_OUT_1_5;
  output CRC_OUT_4_4;
  wire CRC_OUT_4_4;
  output CRC_OUT_5_0;
  wire CRC_OUT_5_0;
  output CRC_OUT_4_22;
  wire CRC_OUT_4_22;
  output CRC_OUT_9_27;
  wire CRC_OUT_9_27;
  output CRC_OUT_9_8;
  wire CRC_OUT_9_8;
  output DATA_9_13;
  wire DATA_9_13;
  output DATA_9_7;
  wire DATA_9_7;
  output CRC_OUT_3_14;
  wire CRC_OUT_3_14;
  output CRC_OUT_3_2;
  wire CRC_OUT_3_2;
  output CRC_OUT_3_5;
  wire CRC_OUT_3_5;
  output CRC_OUT_3_20;
  wire CRC_OUT_3_20;
  output CRC_OUT_8_2;
  wire CRC_OUT_8_2;
  output CRC_OUT_7_17;
  wire CRC_OUT_7_17;
  output CRC_OUT_2_24;
  wire CRC_OUT_2_24;
  output CRC_OUT_8_25;
  wire CRC_OUT_8_25;
  output DATA_9_1;
  wire DATA_9_1;
  output CRC_OUT_2_16;
  wire CRC_OUT_2_16;
  output CRC_OUT_5_29;
  wire CRC_OUT_5_29;
  output DATA_9_29;
  wire DATA_9_29;
  output CRC_OUT_2_22;
  wire CRC_OUT_2_22;
  output CRC_OUT_4_19;
  wire CRC_OUT_4_19;
  output DATA_9_27;
  wire DATA_9_27;
  output CRC_OUT_1_15;
  wire CRC_OUT_1_15;
  output CRC_OUT_2_4;
  wire CRC_OUT_2_4;
  output CRC_OUT_9_28;
  wire CRC_OUT_9_28;
  output CRC_OUT_4_5;
  wire CRC_OUT_4_5;
  output CRC_OUT_2_7;
  wire CRC_OUT_2_7;
  output DATA_9_30;
  wire DATA_9_30;
  output CRC_OUT_5_30;
  wire CRC_OUT_5_30;
  output CRC_OUT_2_23;
  wire CRC_OUT_2_23;
  output CRC_OUT_6_31;
  wire CRC_OUT_6_31;
  output CRC_OUT_1_17;
  wire CRC_OUT_1_17;
  output CRC_OUT_4_7;
  wire CRC_OUT_4_7;
  output CRC_OUT_4_25;
  wire CRC_OUT_4_25;
  output CRC_OUT_6_14;
  wire CRC_OUT_6_14;
  output CRC_OUT_3_18;
  wire CRC_OUT_3_18;
  output CRC_OUT_5_26;
  wire CRC_OUT_5_26;
  output CRC_OUT_5_28;
  wire CRC_OUT_5_28;
  output CRC_OUT_1_27;
  wire CRC_OUT_1_27;
  output CRC_OUT_7_12;
  wire CRC_OUT_7_12;
  output CRC_OUT_3_28;
  wire CRC_OUT_3_28;
  output CRC_OUT_9_16;
  wire CRC_OUT_9_16;
  output CRC_OUT_4_12;
  wire CRC_OUT_4_12;
  output CRC_OUT_7_7;
  wire CRC_OUT_7_7;
  output CRC_OUT_4_15;
  wire CRC_OUT_4_15;
  output CRC_OUT_6_10;
  wire CRC_OUT_6_10;
  output DATA_9_25;
  wire DATA_9_25;
  output CRC_OUT_7_8;
  wire CRC_OUT_7_8;
  output CRC_OUT_9_30;
  wire CRC_OUT_9_30;
  output CRC_OUT_8_1;
  wire CRC_OUT_8_1;
  output CRC_OUT_8_16;
  wire CRC_OUT_8_16;
  output CRC_OUT_3_31;
  wire CRC_OUT_3_31;
  output CRC_OUT_1_3;
  wire CRC_OUT_1_3;
  output CRC_OUT_2_30;
  wire CRC_OUT_2_30;
  output CRC_OUT_4_8;
  wire CRC_OUT_4_8;
  output CRC_OUT_1_23;
  wire CRC_OUT_1_23;
  output CRC_OUT_8_30;
  wire CRC_OUT_8_30;
  output CRC_OUT_6_1;
  wire CRC_OUT_6_1;
  output CRC_OUT_8_7;
  wire CRC_OUT_8_7;
  output CRC_OUT_8_8;
  wire CRC_OUT_8_8;
  output CRC_OUT_9_13;
  wire CRC_OUT_9_13;
  output CRC_OUT_5_11;
  wire CRC_OUT_5_11;
  output CRC_OUT_1_0;
  wire CRC_OUT_1_0;
  output CRC_OUT_3_29;
  wire CRC_OUT_3_29;
  output CRC_OUT_7_9;
  wire CRC_OUT_7_9;
  output CRC_OUT_5_8;
  wire CRC_OUT_5_8;
  output CRC_OUT_5_21;
  wire CRC_OUT_5_21;
  output CRC_OUT_9_2;
  wire CRC_OUT_9_2;
  output CRC_OUT_2_0;
  wire CRC_OUT_2_0;
  output DATA_9_26;
  wire DATA_9_26;
  output CRC_OUT_3_17;
  wire CRC_OUT_3_17;
  output CRC_OUT_8_15;
  wire CRC_OUT_8_15;
  output DATA_9_2;
  wire DATA_9_2;
  output CRC_OUT_2_28;
  wire CRC_OUT_2_28;
  output DATA_9_14;
  wire DATA_9_14;
  output CRC_OUT_9_17;
  wire CRC_OUT_9_17;
  output CRC_OUT_9_3;
  wire CRC_OUT_9_3;
  output DATA_9_9;
  wire DATA_9_9;
  output CRC_OUT_8_17;
  wire CRC_OUT_8_17;
  output DATA_9_19;
  wire DATA_9_19;
  output DATA_9_10;
  wire DATA_9_10;
  output CRC_OUT_7_13;
  wire CRC_OUT_7_13;
  output CRC_OUT_7_23;
  wire CRC_OUT_7_23;
  output CRC_OUT_2_1;
  wire CRC_OUT_2_1;
  output CRC_OUT_1_26;
  wire CRC_OUT_1_26;
  output CRC_OUT_9_9;
  wire CRC_OUT_9_9;
  output CRC_OUT_8_14;
  wire CRC_OUT_8_14;
  output CRC_OUT_1_14;
  wire CRC_OUT_1_14;
  output CRC_OUT_7_16;
  wire CRC_OUT_7_16;
  output CRC_OUT_3_23;
  wire CRC_OUT_3_23;
  output CRC_OUT_8_13;
  wire CRC_OUT_8_13;
  output CRC_OUT_9_23;
  wire CRC_OUT_9_23;
  output CRC_OUT_8_19;
  wire CRC_OUT_8_19;
  output DATA_9_23;
  wire DATA_9_23;
  output CRC_OUT_8_28;
  wire CRC_OUT_8_28;
  output CRC_OUT_9_18;
  wire CRC_OUT_9_18;
  output CRC_OUT_1_21;
  wire CRC_OUT_1_21;
  output CRC_OUT_4_1;
  wire CRC_OUT_4_1;
  output CRC_OUT_1_24;
  wire CRC_OUT_1_24;
  output CRC_OUT_2_21;
  wire CRC_OUT_2_21;
  output CRC_OUT_4_26;
  wire CRC_OUT_4_26;
  output CRC_OUT_6_2;
  wire CRC_OUT_6_2;
  output CRC_OUT_7_25;
  wire CRC_OUT_7_25;
  output CRC_OUT_3_25;
  wire CRC_OUT_3_25;
  output CRC_OUT_9_12;
  wire CRC_OUT_9_12;
  output CRC_OUT_9_15;
  wire CRC_OUT_9_15;
  output DATA_9_22;
  wire DATA_9_22;
  output CRC_OUT_1_1;
  wire CRC_OUT_1_1;
  output DATA_9_5;
  wire DATA_9_5;
  output CRC_OUT_8_0;
  wire CRC_OUT_8_0;
  output DATA_9_31;
  wire DATA_9_31;
  output CRC_OUT_7_21;
  wire CRC_OUT_7_21;
  output DATA_9_16;
  wire DATA_9_16;
  output CRC_OUT_2_13;
  wire CRC_OUT_2_13;
  output CRC_OUT_9_10;
  wire CRC_OUT_9_10;
  output DATA_9_28;
  wire DATA_9_28;
  output CRC_OUT_8_4;
  wire CRC_OUT_8_4;
  output CRC_OUT_4_29;
  wire CRC_OUT_4_29;
  output CRC_OUT_6_8;
  wire CRC_OUT_6_8;
  output CRC_OUT_3_13;
  wire CRC_OUT_3_13;
  output CRC_OUT_3_30;
  wire CRC_OUT_3_30;
  output CRC_OUT_1_30;
  wire CRC_OUT_1_30;
  output CRC_OUT_8_5;
  wire CRC_OUT_8_5;
  output CRC_OUT_6_15;
  wire CRC_OUT_6_15;
  output CRC_OUT_6_5;
  wire CRC_OUT_6_5;
  output CRC_OUT_1_10;
  wire CRC_OUT_1_10;
  output CRC_OUT_7_18;
  wire CRC_OUT_7_18;
  output CRC_OUT_4_9;
  wire CRC_OUT_4_9;
  output CRC_OUT_1_13;
  wire CRC_OUT_1_13;
  output CRC_OUT_8_27;
  wire CRC_OUT_8_27;
  output CRC_OUT_5_2;
  wire CRC_OUT_5_2;
  output CRC_OUT_8_12;
  wire CRC_OUT_8_12;
  output CRC_OUT_8_22;
  wire CRC_OUT_8_22;
  output CRC_OUT_7_11;
  wire CRC_OUT_7_11;
  output CRC_OUT_7_10;
  wire CRC_OUT_7_10;
  output CRC_OUT_6_25;
  wire CRC_OUT_6_25;
  output CRC_OUT_6_23;
  wire CRC_OUT_6_23;
  output CRC_OUT_1_9;
  wire CRC_OUT_1_9;
  output CRC_OUT_7_0;
  wire CRC_OUT_7_0;
  output CRC_OUT_7_1;
  wire CRC_OUT_7_1;
  output CRC_OUT_4_21;
  wire CRC_OUT_4_21;
  output CRC_OUT_9_0;
  wire CRC_OUT_9_0;
  output CRC_OUT_1_2;
  wire CRC_OUT_1_2;
  output CRC_OUT_6_17;
  wire CRC_OUT_6_17;
  output CRC_OUT_5_10;
  wire CRC_OUT_5_10;
  output CRC_OUT_8_9;
  wire CRC_OUT_8_9;
  output CRC_OUT_7_24;
  wire CRC_OUT_7_24;
  output CRC_OUT_5_22;
  wire CRC_OUT_5_22;
  output CRC_OUT_7_14;
  wire CRC_OUT_7_14;
  output DATA_9_18;
  wire DATA_9_18;
  output CRC_OUT_7_28;
  wire CRC_OUT_7_28;
  output CRC_OUT_3_22;
  wire CRC_OUT_3_22;
  output CRC_OUT_6_29;
  wire CRC_OUT_6_29;
  output CRC_OUT_8_20;
  wire CRC_OUT_8_20;
  output CRC_OUT_6_22;
  wire CRC_OUT_6_22;
  output CRC_OUT_5_17;
  wire CRC_OUT_5_17;
  output CRC_OUT_3_1;
  wire CRC_OUT_3_1;
  output CRC_OUT_3_19;
  wire CRC_OUT_3_19;
  output CRC_OUT_5_9;
  wire CRC_OUT_5_9;
  output CRC_OUT_3_4;
  wire CRC_OUT_3_4;
  output CRC_OUT_1_18;
  wire CRC_OUT_1_18;
  output CRC_OUT_5_16;
  wire CRC_OUT_5_16;
  output CRC_OUT_6_4;
  wire CRC_OUT_6_4;
  output CRC_OUT_8_24;
  wire CRC_OUT_8_24;
  output CRC_OUT_2_10;
  wire CRC_OUT_2_10;
  output DATA_9_24;
  wire DATA_9_24;
  output CRC_OUT_8_23;
  wire CRC_OUT_8_23;
  output CRC_OUT_8_18;
  wire CRC_OUT_8_18;
  output CRC_OUT_1_8;
  wire CRC_OUT_1_8;
  output CRC_OUT_2_31;
  wire CRC_OUT_2_31;
  output CRC_OUT_2_19;
  wire CRC_OUT_2_19;
  output CRC_OUT_4_16;
  wire CRC_OUT_4_16;
  output CRC_OUT_7_31;
  wire CRC_OUT_7_31;
  output CRC_OUT_2_18;
  wire CRC_OUT_2_18;
  output CRC_OUT_4_6;
  wire CRC_OUT_4_6;
  output CRC_OUT_2_9;
  wire CRC_OUT_2_9;
  output CRC_OUT_5_31;
  wire CRC_OUT_5_31;
  output CRC_OUT_5_18;
  wire CRC_OUT_5_18;
  output CRC_OUT_6_27;
  wire CRC_OUT_6_27;
  output CRC_OUT_3_21;
  wire CRC_OUT_3_21;
  output CRC_OUT_1_25;
  wire CRC_OUT_1_25;
  output CRC_OUT_4_30;
  wire CRC_OUT_4_30;
  output DATA_9_3;
  wire DATA_9_3;
  output CRC_OUT_1_12;
  wire CRC_OUT_1_12;
  output CRC_OUT_7_6;
  wire CRC_OUT_7_6;
  output CRC_OUT_9_1;
  wire CRC_OUT_9_1;
  output CRC_OUT_5_15;
  wire CRC_OUT_5_15;
  output CRC_OUT_5_27;
  wire CRC_OUT_5_27;
  output CRC_OUT_7_30;
  wire CRC_OUT_7_30;
  output CRC_OUT_3_26;
  wire CRC_OUT_3_26;
  output CRC_OUT_3_0;
  wire CRC_OUT_3_0;
  output CRC_OUT_1_29;
  wire CRC_OUT_1_29;
  output CRC_OUT_9_20;
  wire CRC_OUT_9_20;
  output DATA_9_12;
  wire DATA_9_12;
  output CRC_OUT_6_12;
  wire CRC_OUT_6_12;
  output DATA_9_6;
  wire DATA_9_6;
  output CRC_OUT_4_20;
  wire CRC_OUT_4_20;
  output CRC_OUT_4_28;
  wire CRC_OUT_4_28;
  wire __0__;
  wire __1__;
  wire __2__;
  wire __3__;
  wire __4__;
  wire __5__;
  wire __6__;
  wire __7__;
  wire __8__;
  wire __9__;
  wire __10__;
  wire __11__;
  wire __12__;
  wire __13__;
  wire __14__;
  wire __15__;
  wire __16__;
  wire __17__;
  wire __18__;
  wire __19__;
  wire __20__;
  wire __21__;
  wire __22__;
  wire __23__;
  wire __24__;
  wire __25__;
  wire __26__;
  wire __27__;
  wire __28__;
  wire __29__;
  wire __30__;
  wire __31__;
  wire __32__;
  wire __33__;
  wire __34__;
  wire __35__;
  wire __36__;
  wire __37__;
  wire __38__;
  wire __39__;
  wire __40__;
  wire __41__;
  wire __42__;
  wire __43__;
  wire __44__;
  wire __45__;
  wire __46__;
  wire __47__;
  wire __48__;
  wire __49__;
  wire __50__;
  wire __51__;
  wire __52__;
  wire __53__;
  wire __54__;
  wire __55__;
  wire __56__;
  wire __57__;
  wire __58__;
  wire __59__;
  wire __60__;
  wire __61__;
  wire __62__;
  wire __63__;
  wire __64__;
  wire __65__;
  wire __66__;
  wire __67__;
  wire __68__;
  wire __69__;
  wire __70__;
  wire __71__;
  wire __72__;
  wire __73__;
  wire __74__;
  wire __75__;
  wire __76__;
  wire __77__;
  wire __78__;
  wire __79__;
  wire __80__;
  wire __81__;
  wire __82__;
  wire __83__;
  wire __84__;
  wire __85__;
  wire __86__;
  wire __87__;
  wire __88__;
  wire __89__;
  wire __90__;
  wire __91__;
  wire __92__;
  wire __93__;
  wire __94__;
  wire __95__;
  wire __96__;
  wire __97__;
  wire __98__;
  wire __99__;
  wire __100__;
  wire __101__;
  wire __102__;
  wire __103__;
  wire __104__;
  wire __105__;
  wire __106__;
  wire __107__;
  wire __108__;
  wire __109__;
  wire __110__;
  wire __111__;
  wire __112__;
  wire __113__;
  wire __114__;
  wire __115__;
  wire __116__;
  wire __117__;
  wire __118__;
  wire __119__;
  wire __120__;
  wire __121__;
  wire __122__;
  wire __123__;
  wire __124__;
  wire __125__;
  wire __126__;
  wire __127__;
  wire __128__;
  wire __129__;
  wire __130__;
  wire __131__;
  wire __132__;
  wire __133__;
  wire __134__;
  wire __135__;
  wire __136__;
  wire __137__;
  wire __138__;
  wire __139__;
  wire __140__;
  wire __141__;
  wire __142__;
  wire __143__;
  wire __144__;
  wire __145__;
  wire __146__;
  wire __147__;
  wire __148__;
  wire __149__;
  wire __150__;
  wire __151__;
  wire __152__;
  wire __153__;
  wire __154__;
  wire __155__;
  wire __156__;
  wire __157__;
  wire __158__;
  wire __159__;
  wire __160__;
  wire __161__;
  wire __162__;
  wire __163__;
  wire __164__;
  wire __165__;
  wire __166__;
  wire __167__;
  wire __168__;
  wire __169__;
  wire __170__;
  wire __171__;
  wire __172__;
  wire __173__;
  wire __174__;
  wire __175__;
  wire __176__;
  wire __177__;
  wire __178__;
  wire __179__;
  wire __180__;
  wire __181__;
  wire __182__;
  wire __183__;
  wire __184__;
  wire __185__;
  wire __186__;
  wire __187__;
  wire __188__;
  wire __189__;
  wire __190__;
  wire __191__;
  wire __192__;
  wire __193__;
  wire __194__;
  wire __195__;
  wire __196__;
  wire __197__;
  wire __198__;
  wire __199__;
  wire __200__;
  wire __201__;
  wire __202__;
  wire __203__;
  wire __204__;
  wire __205__;
  wire __206__;
  wire __207__;
  wire __208__;
  wire __209__;
  wire __210__;
  wire __211__;
  wire __212__;
  wire __213__;
  wire __214__;
  wire __215__;
  wire __216__;
  wire __217__;
  wire __218__;
  wire __219__;
  wire __220__;
  wire __221__;
  wire __222__;
  wire __223__;
  wire __224__;
  wire __225__;
  wire __226__;
  wire __227__;
  wire __228__;
  wire __229__;
  wire __230__;
  wire __231__;
  wire __232__;
  wire __233__;
  wire __234__;
  wire __235__;
  wire __236__;
  wire __237__;
  wire __238__;
  wire __239__;
  wire __240__;
  wire __241__;
  wire __242__;
  wire __243__;
  wire __244__;
  wire __245__;
  wire __246__;
  wire __247__;
  wire __248__;
  wire __249__;
  wire __250__;
  wire __251__;
  wire __252__;
  wire __253__;
  wire __254__;
  wire __255__;
  wire __256__;
  wire __257__;
  wire __258__;
  wire __259__;
  wire __260__;
  wire __261__;
  wire __262__;
  wire __263__;
  wire __264__;
  wire __265__;
  wire __266__;
  wire __267__;
  wire __268__;
  wire __269__;
  wire __270__;
  wire __271__;
  wire __272__;
  wire __273__;
  wire __274__;
  wire __275__;
  wire __276__;
  wire __277__;
  wire __278__;
  wire __279__;
  wire __280__;
  wire __281__;
  wire __282__;
  wire __283__;
  wire __284__;
  wire __285__;
  wire __286__;
  wire __287__;
  wire __288__;
  wire __289__;
  wire __290__;
  wire __291__;
  wire __292__;
  wire __293__;
  wire __294__;
  wire __295__;
  wire __296__;
  wire __297__;
  wire __298__;
  wire __299__;
  wire __300__;
  wire __301__;
  wire __302__;
  wire __303__;
  wire __304__;
  wire __305__;
  wire __306__;
  wire __307__;
  wire __308__;
  wire __309__;
  wire __310__;
  wire __311__;
  wire __312__;
  wire __313__;
  wire __314__;
  wire __315__;
  wire __316__;
  wire __317__;
  wire __318__;
  wire __319__;
  wire __320__;
  wire __321__;
  wire __322__;
  wire __323__;
  wire __324__;
  wire __325__;
  wire __326__;
  wire __327__;
  wire __328__;
  wire __329__;
  wire __330__;
  wire __331__;
  wire __332__;
  wire __333__;
  wire __334__;
  wire __335__;
  wire __336__;
  wire __337__;
  wire __338__;
  wire __339__;
  wire __340__;
  wire __341__;
  wire __342__;
  wire __343__;
  wire __344__;
  wire __345__;
  wire __346__;
  wire __347__;
  wire __348__;
  wire __349__;
  wire __350__;
  wire __351__;
  wire __352__;
  wire __353__;
  wire __354__;
  wire __355__;
  wire __356__;
  wire __357__;
  wire __358__;
  wire __359__;
  wire __360__;
  wire __361__;
  wire __362__;
  wire __363__;
  wire __364__;
  wire __365__;
  wire __366__;
  wire __367__;
  wire __368__;
  wire __369__;
  wire __370__;
  wire __371__;
  wire __372__;
  wire __373__;
  wire __374__;
  wire __375__;
  wire __376__;
  wire __377__;
  wire __378__;
  wire __379__;
  wire __380__;
  wire __381__;
  wire __382__;
  wire __383__;
  wire __384__;
  wire __385__;
  wire __386__;
  wire __387__;
  wire __388__;
  wire __389__;
  wire __390__;
  wire __391__;
  wire __392__;
  wire __393__;
  wire __394__;
  wire __395__;
  wire __396__;
  wire __397__;
  wire __398__;
  wire __399__;
  wire __400__;
  wire __401__;
  wire __402__;
  wire __403__;
  wire __404__;
  wire __405__;
  wire __406__;
  wire __407__;
  wire __408__;
  wire __409__;
  wire __410__;
  wire __411__;
  wire __412__;
  wire __413__;
  wire __414__;
  wire __415__;
  wire __416__;
  wire __417__;
  wire __418__;
  wire __419__;
  wire __420__;
  wire __421__;
  wire __422__;
  wire __423__;
  wire __424__;
  wire __425__;
  wire __426__;
  wire __427__;
  wire __428__;
  wire __429__;
  wire __430__;
  wire __431__;
  wire __432__;
  wire __433__;
  wire __434__;
  wire __435__;
  wire __436__;
  wire __437__;
  wire __438__;
  wire __439__;
  wire __440__;
  wire __441__;
  wire __442__;
  wire __443__;
  wire __444__;
  wire __445__;
  wire __446__;
  wire __447__;
  wire __448__;
  wire __449__;
  wire __450__;
  wire __451__;
  wire __452__;
  wire __453__;
  wire __454__;
  wire __455__;
  wire __456__;
  wire __457__;
  wire __458__;
  wire __459__;
  wire __460__;
  wire __461__;
  wire __462__;
  wire __463__;
  wire __464__;
  wire __465__;
  wire __466__;
  wire __467__;
  wire __468__;
  wire __469__;
  wire __470__;
  wire __471__;
  wire __472__;
  wire __473__;
  wire __474__;
  wire __475__;
  wire __476__;
  wire __477__;
  wire __478__;
  wire __479__;
  wire __480__;
  wire __481__;
  wire __482__;
  wire __483__;
  wire __484__;
  wire __485__;
  wire __486__;
  wire __487__;
  wire __488__;
  wire __489__;
  wire __490__;
  wire __491__;
  wire __492__;
  wire __493__;
  wire __494__;
  wire __495__;
  wire __496__;
  wire __497__;
  wire __498__;
  wire __499__;
  wire __500__;
  wire __501__;
  wire __502__;
  wire __503__;
  wire __504__;
  wire __505__;
  wire __506__;
  wire __507__;
  wire __508__;
  wire __509__;
  wire __510__;
  wire __511__;
  wire __512__;
  wire __513__;
  wire __514__;
  wire __515__;
  wire __516__;
  wire __517__;
  wire __518__;
  wire __519__;
  wire __520__;
  wire __521__;
  wire __522__;
  wire __523__;
  wire __524__;
  wire __525__;
  wire __526__;
  wire __527__;
  wire __528__;
  wire __529__;
  wire __530__;
  wire __531__;
  wire __532__;
  wire __533__;
  wire __534__;
  wire __535__;
  wire __536__;
  wire __537__;
  wire __538__;
  wire __539__;
  wire __540__;
  wire __541__;
  wire __542__;
  wire __543__;
  wire __544__;
  wire __545__;
  wire __546__;
  wire __547__;
  wire __548__;
  wire __549__;
  wire __550__;
  wire __551__;
  wire __552__;
  wire __553__;
  wire __554__;
  wire __555__;
  wire __556__;
  wire __557__;
  wire __558__;
  wire __559__;
  wire __560__;
  wire __561__;
  wire __562__;
  wire __563__;
  wire __564__;
  wire __565__;
  wire __566__;
  wire __567__;
  wire __568__;
  wire __569__;
  wire __570__;
  wire __571__;
  wire __572__;
  wire __573__;
  wire __574__;
  wire __575__;
  wire __576__;
  wire __577__;
  wire __578__;
  wire __579__;
  wire __580__;
  wire __581__;
  wire __582__;
  wire __583__;
  wire __584__;
  wire __585__;
  wire __586__;
  wire __587__;
  wire __588__;
  wire __589__;
  wire __590__;
  wire __591__;
  wire __592__;
  wire __593__;
  wire __594__;
  wire __595__;
  wire __596__;
  wire __597__;
  wire __598__;
  wire __599__;
  wire __600__;
  wire __601__;
  wire __602__;
  wire __603__;
  wire __604__;
  wire __605__;
  wire __606__;
  wire __607__;
  wire __608__;
  wire __609__;
  wire __610__;
  wire __611__;
  wire __612__;
  wire __613__;
  wire __614__;
  wire __615__;
  wire __616__;
  wire __617__;
  wire __618__;
  wire __619__;
  wire __620__;
  wire __621__;
  wire __622__;
  wire __623__;
  wire __624__;
  wire __625__;
  wire __626__;
  wire __627__;
  wire __628__;
  wire __629__;
  wire __630__;
  wire __631__;
  wire __632__;
  wire __633__;
  wire __634__;
  wire __635__;
  wire __636__;
  wire __637__;
  wire __638__;
  wire __639__;
  wire __640__;
  wire __641__;
  wire __642__;
  wire __643__;
  wire __644__;
  wire __645__;
  wire __646__;
  wire __647__;
  wire __648__;
  wire __649__;
  wire __650__;
  wire __651__;
  wire __652__;
  wire __653__;
  wire __654__;
  wire __655__;
  wire __656__;
  wire __657__;
  wire __658__;
  wire __659__;
  wire __660__;
  wire __661__;
  wire __662__;
  wire __663__;
  wire __664__;
  wire __665__;
  wire __666__;
  wire __667__;
  wire __668__;
  wire __669__;
  wire __670__;
  wire __671__;
  wire __672__;
  wire __673__;
  wire __674__;
  wire __675__;
  wire __676__;
  wire __677__;
  wire __678__;
  wire __679__;
  wire __680__;
  wire __681__;
  wire __682__;
  wire __683__;
  wire __684__;
  wire __685__;
  wire __686__;
  wire __687__;
  wire __688__;
  wire __689__;
  wire __690__;
  wire __691__;
  wire __692__;
  wire __693__;
  wire __694__;
  wire __695__;
  wire __696__;
  wire __697__;
  wire __698__;
  wire __699__;
  wire __700__;
  wire __701__;
  wire __702__;
  wire __703__;
  wire __704__;
  wire __705__;
  wire __706__;
  wire __707__;
  wire __708__;
  wire __709__;
  wire __710__;
  wire __711__;
  wire __712__;
  wire __713__;
  wire __714__;
  wire __715__;
  wire __716__;
  wire __717__;
  wire __718__;
  wire __719__;
  wire __720__;
  wire __721__;
  wire __722__;
  wire __723__;
  wire __724__;
  wire __725__;
  wire __726__;
  wire __727__;
  wire __728__;
  wire __729__;
  wire __730__;
  wire __731__;
  wire __732__;
  wire __733__;
  wire __734__;
  wire __735__;
  wire __736__;
  wire __737__;
  wire __738__;
  wire __739__;
  wire __740__;
  wire __741__;
  wire __742__;
  wire __743__;
  wire __744__;
  wire __745__;
  wire __746__;
  wire __747__;
  wire __748__;
  wire __749__;
  wire __750__;
  wire __751__;
  wire __752__;
  wire __753__;
  wire __754__;
  wire __755__;
  wire __756__;
  wire __757__;
  wire __758__;
  wire __759__;
  wire __760__;
  wire __761__;
  wire __762__;
  wire __763__;
  wire __764__;
  wire __765__;
  wire __766__;
  wire __767__;
  wire __768__;
  wire __769__;
  wire __770__;
  wire __771__;
  wire __772__;
  wire __773__;
  wire __774__;
  wire __775__;
  wire __776__;
  wire __777__;
  wire __778__;
  wire __779__;
  wire __780__;
  wire __781__;
  wire __782__;
  wire __783__;
  wire __784__;
  wire __785__;
  wire __786__;
  wire __787__;
  wire __788__;
  wire __789__;
  wire __790__;
  wire __791__;
  wire __792__;
  wire __793__;
  wire __794__;
  wire __795__;
  wire __796__;
  wire __797__;
  wire __798__;
  wire __799__;
  wire __800__;
  wire __801__;
  wire __802__;
  wire __803__;
  wire __804__;
  wire __805__;
  wire __806__;
  wire __807__;
  wire __808__;
  wire __809__;
  wire __810__;
  wire __811__;
  wire __812__;
  wire __813__;
  wire __814__;
  wire __815__;
  wire __816__;
  wire __817__;
  wire __818__;
  wire __819__;
  wire __820__;
  wire __821__;
  wire __822__;
  wire __823__;
  wire __824__;
  wire __825__;
  wire __826__;
  wire __827__;
  wire __828__;
  wire __829__;
  wire __830__;
  wire __831__;
  wire __832__;
  wire __833__;
  wire __834__;
  wire __835__;
  wire __836__;
  wire __837__;
  wire __838__;
  wire __839__;
  wire __840__;
  wire __841__;
  wire __842__;
  wire __843__;
  wire __844__;
  wire __845__;
  wire __846__;
  wire __847__;
  wire __848__;
  wire __849__;
  wire __850__;
  wire __851__;
  wire __852__;
  wire __853__;
  wire __854__;
  wire __855__;
  wire __856__;
  wire __857__;
  wire __858__;
  wire __859__;
  wire __860__;
  wire __861__;
  wire __862__;
  wire __863__;
  wire __864__;
  wire __865__;
  wire __866__;
  wire __867__;
  wire __868__;
  wire __869__;
  wire __870__;
  wire __871__;
  wire __872__;
  wire __873__;
  wire __874__;
  wire __875__;
  wire __876__;
  wire __877__;
  wire __878__;
  wire __879__;
  wire __880__;
  wire __881__;
  wire __882__;
  wire __883__;
  wire __884__;
  wire __885__;
  wire __886__;
  wire __887__;
  wire __888__;
  wire __889__;
  wire __890__;
  wire __891__;
  wire __892__;
  wire __893__;
  wire __894__;
  wire __895__;
  wire __896__;
  wire __897__;
  wire __898__;
  wire __899__;
  wire __900__;
  wire __901__;
  wire __902__;
  wire __903__;
  wire __904__;
  wire __905__;
  wire __906__;
  wire __907__;
  wire __908__;
  wire __909__;
  wire __910__;
  wire __911__;
  wire __912__;
  wire __913__;
  wire __914__;
  wire __915__;
  wire __916__;
  wire __917__;
  wire __918__;
  wire __919__;
  wire __920__;
  wire __921__;
  wire __922__;
  wire __923__;
  wire __924__;
  wire __925__;
  wire __926__;
  wire __927__;
  wire __928__;
  wire __929__;
  wire __930__;
  wire __931__;
  wire __932__;
  wire __933__;
  wire __934__;
  wire __935__;
  wire __936__;
  wire __937__;
  wire __938__;
  wire __939__;
  wire __940__;
  wire __941__;
  wire __942__;
  wire __943__;
  wire __944__;
  wire __945__;
  wire __946__;
  wire __947__;
  wire __948__;
  wire __949__;
  wire __950__;
  wire __951__;
  wire __952__;
  wire __953__;
  wire __954__;
  wire __955__;
  wire __956__;
  wire __957__;
  wire __958__;
  wire __959__;
  wire __960__;
  wire __961__;
  wire __962__;
  wire __963__;
  wire __964__;
  wire __965__;
  wire __966__;
  wire __967__;
  wire __968__;
  wire __969__;
  wire __970__;
  wire __971__;
  wire __972__;
  wire __973__;
  wire __974__;
  wire __975__;
  wire __976__;
  wire __977__;
  wire __978__;
  wire __979__;
  wire __980__;
  wire __981__;
  wire __982__;
  wire __983__;
  wire __984__;
  wire __985__;
  wire __986__;
  wire __987__;
  wire __988__;
  wire __989__;
  wire __990__;
  wire __991__;
  wire __992__;
  wire __993__;
  wire __994__;
  wire __995__;
  wire __996__;
  wire __997__;
  wire __998__;
  wire __999__;
  wire __1000__;
  wire __1001__;
  wire __1002__;
  wire __1003__;
  wire __1004__;
  wire __1005__;
  wire __1006__;
  wire __1007__;
  wire __1008__;
  wire __1009__;
  wire __1010__;
  wire __1011__;
  wire __1012__;
  wire __1013__;
  wire __1014__;
  wire __1015__;
  wire __1016__;
  wire __1017__;
  wire __1018__;
  wire __1019__;
  wire __1020__;
  wire __1021__;
  wire __1022__;
  wire __1023__;
  wire __1024__;
  wire __1025__;
  wire __1026__;
  wire __1027__;
  wire __1028__;
  wire __1029__;
  wire __1030__;
  wire __1031__;
  wire __1032__;
  wire __1033__;
  wire __1034__;
  wire __1035__;
  wire __1036__;
  wire __1037__;
  wire __1038__;
  wire __1039__;
  wire __1040__;
  wire __1041__;
  wire __1042__;
  wire __1043__;
  wire __1044__;
  wire __1045__;
  wire __1046__;
  wire __1047__;
  wire __1048__;
  wire __1049__;
  wire __1050__;
  wire __1051__;
  wire __1052__;
  wire __1053__;
  wire __1054__;
  wire __1055__;
  wire __1056__;
  wire __1057__;
  wire __1058__;
  wire __1059__;
  wire __1060__;
  wire __1061__;
  wire __1062__;
  wire __1063__;
  wire __1064__;
  wire __1065__;
  wire __1066__;
  wire __1067__;
  wire __1068__;
  wire __1069__;
  wire __1070__;
  wire __1071__;
  wire __1072__;
  wire __1073__;
  wire __1074__;
  wire __1075__;
  wire __1076__;
  wire __1077__;
  wire __1078__;
  wire __1079__;
  wire __1080__;
  wire __1081__;
  wire __1082__;
  wire __1083__;
  wire __1084__;
  wire __1085__;
  wire __1086__;
  wire __1087__;
  wire __1088__;
  wire __1089__;
  wire __1090__;
  wire __1091__;
  wire __1092__;
  wire __1093__;
  wire __1094__;
  wire __1095__;
  wire __1096__;
  wire __1097__;
  wire __1098__;
  wire __1099__;
  wire __1100__;
  wire __1101__;
  wire __1102__;
  wire __1103__;
  wire __1104__;
  wire __1105__;
  wire __1106__;
  wire __1107__;
  wire __1108__;
  wire __1109__;
  wire __1110__;
  wire __1111__;
  wire __1112__;
  wire __1113__;
  wire __1114__;
  wire __1115__;
  wire __1116__;
  wire __1117__;
  wire __1118__;
  wire __1119__;
  wire __1120__;
  wire __1121__;
  wire __1122__;
  wire __1123__;
  wire __1124__;
  wire __1125__;
  wire __1126__;
  wire __1127__;
  wire __1128__;
  wire __1129__;
  wire __1130__;
  wire __1131__;
  wire __1132__;
  wire __1133__;
  wire __1134__;
  wire __1135__;
  wire __1136__;
  wire __1137__;
  wire __1138__;
  wire __1139__;
  wire __1140__;
  wire __1141__;
  wire __1142__;
  wire __1143__;
  wire __1144__;
  wire __1145__;
  wire __1146__;
  wire __1147__;
  wire __1148__;
  wire __1149__;
  wire __1150__;
  wire __1151__;
  wire __1152__;
  wire __1153__;
  wire __1154__;
  wire __1155__;
  wire __1156__;
  wire __1157__;
  wire __1158__;
  wire __1159__;
  wire __1160__;
  wire __1161__;
  wire __1162__;
  wire __1163__;
  wire __1164__;
  wire __1165__;
  wire __1166__;
  wire __1167__;
  wire __1168__;
  wire __1169__;
  wire __1170__;
  wire __1171__;
  wire __1172__;
  wire __1173__;
  wire __1174__;
  wire __1175__;
  wire __1176__;
  wire __1177__;
  wire __1178__;
  wire __1179__;
  wire __1180__;
  wire __1181__;
  wire __1182__;
  wire __1183__;
  wire __1184__;
  wire __1185__;
  wire __1186__;
  wire __1187__;
  wire __1188__;
  wire __1189__;
  wire __1190__;
  wire __1191__;
  wire __1192__;
  wire __1193__;
  wire __1194__;
  wire __1195__;
  wire __1196__;
  wire __1197__;
  wire __1198__;
  wire __1199__;
  wire __1200__;
  wire __1201__;
  wire __1202__;
  wire __1203__;
  wire __1204__;
  wire __1205__;
  wire __1206__;
  wire __1207__;
  wire __1208__;
  wire __1209__;
  wire __1210__;
  wire __1211__;
  wire __1212__;
  wire __1213__;
  wire __1214__;
  wire __1215__;
  wire __1216__;
  wire __1217__;
  wire __1218__;
  wire __1219__;
  wire __1220__;
  wire __1221__;
  wire __1222__;
  wire __1223__;
  wire __1224__;
  wire __1225__;
  wire __1226__;
  wire __1227__;
  wire __1228__;
  wire __1229__;
  wire __1230__;
  wire __1231__;
  wire __1232__;
  wire __1233__;
  wire __1234__;
  wire __1235__;
  wire __1236__;
  wire __1237__;
  wire __1238__;
  wire __1239__;
  wire __1240__;
  wire __1241__;
  wire __1242__;
  wire __1243__;
  wire __1244__;
  wire __1245__;
  wire __1246__;
  wire __1247__;
  wire __1248__;
  wire __1249__;
  wire __1250__;
  wire __1251__;
  wire __1252__;
  wire __1253__;
  wire __1254__;
  wire __1255__;
  wire __1256__;
  wire __1257__;
  wire __1258__;
  wire __1259__;
  wire __1260__;
  wire __1261__;
  wire __1262__;
  wire __1263__;
  wire __1264__;
  wire __1265__;
  wire __1266__;
  wire __1267__;
  wire __1268__;
  wire __1269__;
  wire __1270__;
  wire __1271__;
  wire __1272__;
  wire __1273__;
  wire __1274__;
  wire __1275__;
  wire __1276__;
  wire __1277__;
  wire __1278__;
  wire __1279__;
  wire __1280__;
  wire __1281__;
  wire __1282__;
  wire __1283__;
  wire __1284__;
  wire __1285__;
  wire __1286__;
  wire __1287__;
  wire __1288__;
  wire __1289__;
  wire __1290__;
  wire __1291__;
  wire __1292__;
  wire __1293__;
  wire __1294__;
  wire __1295__;
  wire __1296__;
  wire __1297__;
  wire __1298__;
  wire __1299__;
  wire __1300__;
  wire __1301__;
  wire __1302__;
  wire __1303__;
  wire __1304__;
  wire __1305__;
  wire __1306__;
  wire __1307__;
  wire __1308__;
  wire __1309__;
  wire __1310__;
  wire __1311__;
  wire __1312__;
  wire __1313__;
  wire __1314__;
  wire __1315__;
  wire __1316__;
  wire __1317__;
  wire __1318__;
  wire __1319__;
  wire __1320__;
  wire __1321__;
  wire __1322__;
  wire __1323__;
  wire __1324__;
  wire __1325__;
  wire __1326__;
  wire __1327__;
  wire __1328__;
  wire __1329__;
  wire __1330__;
  wire __1331__;
  wire __1332__;
  wire __1333__;
  wire __1334__;
  wire __1335__;
  wire __1336__;
  wire __1337__;
  wire __1338__;
  wire __1339__;
  wire __1340__;
  wire __1341__;
  wire __1342__;
  wire __1343__;
  wire __1344__;
  wire __1345__;
  wire __1346__;
  wire __1347__;
  wire __1348__;
  wire __1349__;
  wire __1350__;
  wire __1351__;
  wire __1352__;
  wire __1353__;
  wire __1354__;
  wire __1355__;
  wire __1356__;
  wire __1357__;
  wire __1358__;
  wire __1359__;
  wire __1360__;
  wire __1361__;
  wire __1362__;
  wire __1363__;
  wire __1364__;
  wire __1365__;
  wire __1366__;
  wire __1367__;
  wire __1368__;
  wire __1369__;
  wire __1370__;
  wire __1371__;
  wire __1372__;
  wire __1373__;
  wire __1374__;
  wire __1375__;
  wire __1376__;
  wire __1377__;
  wire __1378__;
  wire __1379__;
  wire __1380__;
  wire __1381__;
  wire __1382__;
  wire __1383__;
  wire __1384__;
  wire __1385__;
  wire __1386__;
  wire __1387__;
  wire __1388__;
  wire __1389__;
  wire __1390__;
  wire __1391__;
  wire __1392__;
  wire __1393__;
  wire __1394__;
  wire __1395__;
  wire __1396__;
  wire __1397__;
  wire __1398__;
  wire __1399__;
  wire __1400__;
  wire __1401__;
  wire __1402__;
  wire __1403__;
  wire __1404__;
  wire __1405__;
  wire __1406__;
  wire __1407__;
  wire __1408__;
  wire __1409__;
  wire __1410__;
  wire __1411__;
  wire __1412__;
  wire __1413__;
  wire __1414__;
  wire __1415__;
  wire __1416__;
  wire __1417__;
  wire __1418__;
  wire __1419__;
  wire __1420__;
  wire __1421__;
  wire __1422__;
  wire __1423__;
  wire __1424__;
  wire __1425__;
  wire __1426__;
  wire __1427__;
  wire __1428__;
  wire __1429__;
  wire __1430__;
  wire __1431__;
  wire __1432__;
  wire __1433__;
  wire __1434__;
  wire __1435__;
  wire __1436__;
  wire __1437__;
  wire __1438__;
  wire __1439__;
  wire __1440__;
  wire __1441__;
  wire __1442__;
  wire __1443__;
  wire __1444__;
  wire __1445__;
  wire __1446__;
  wire __1447__;
  wire __1448__;
  wire __1449__;
  wire __1450__;
  wire __1451__;
  wire __1452__;
  wire __1453__;
  wire __1454__;
  wire __1455__;
  wire __1456__;
  wire __1457__;
  wire __1458__;
  wire __1459__;
  wire __1460__;
  wire __1461__;
  wire __1462__;
  wire __1463__;
  wire __1464__;
  wire __1465__;
  wire __1466__;
  wire __1467__;
  wire __1468__;
  wire __1469__;
  wire __1470__;
  wire __1471__;
  wire __1472__;
  wire __1473__;
  wire __1474__;
  wire __1475__;
  wire __1476__;
  wire __1477__;
  wire __1478__;
  wire __1479__;
  wire __1480__;
  wire __1481__;
  wire __1482__;
  wire __1483__;
  wire __1484__;
  wire __1485__;
  wire __1486__;
  wire __1487__;
  wire __1488__;
  wire __1489__;
  wire __1490__;
  wire __1491__;
  wire __1492__;
  wire __1493__;
  wire __1494__;
  wire __1495__;
  wire __1496__;
  wire __1497__;
  wire __1498__;
  wire __1499__;
  wire __1500__;
  wire __1501__;
  wire __1502__;
  wire __1503__;
  wire __1504__;
  wire __1505__;
  wire __1506__;
  wire __1507__;
  wire __1508__;
  wire __1509__;
  wire __1510__;
  wire __1511__;
  wire __1512__;
  wire __1513__;
  wire __1514__;
  wire __1515__;
  wire __1516__;
  wire __1517__;
  wire __1518__;
  wire __1519__;
  wire __1520__;
  wire __1521__;
  wire __1522__;
  wire __1523__;
  wire __1524__;
  wire __1525__;
  wire __1526__;
  wire __1527__;
  wire __1528__;
  wire __1529__;
  wire __1530__;
  wire __1531__;
  wire __1532__;
  wire __1533__;
  wire __1534__;
  wire __1535__;
  wire __1536__;
  wire __1537__;
  wire __1538__;
  wire __1539__;
  wire __1540__;
  wire __1541__;
  wire __1542__;
  wire __1543__;
  wire __1544__;
  wire __1545__;
  wire __1546__;
  wire __1547__;
  wire __1548__;
  wire __1549__;
  wire __1550__;
  wire __1551__;
  wire __1552__;
  wire __1553__;
  wire __1554__;
  wire __1555__;
  wire __1556__;
  wire __1557__;
  wire __1558__;
  wire __1559__;
  wire __1560__;
  wire __1561__;
  wire __1562__;
  wire __1563__;
  wire __1564__;
  wire __1565__;
  wire __1566__;
  wire __1567__;
  wire __1568__;
  wire __1569__;
  wire __1570__;
  wire __1571__;
  wire __1572__;
  wire __1573__;
  wire __1574__;
  wire __1575__;
  wire __1576__;
  wire __1577__;
  wire __1578__;
  wire __1579__;
  wire __1580__;
  wire __1581__;
  wire __1582__;
  wire __1583__;
  wire __1584__;
  wire __1585__;
  wire __1586__;
  wire __1587__;
  wire __1588__;
  wire __1589__;
  wire __1590__;
  wire __1591__;
  wire __1592__;
  wire __1593__;
  wire __1594__;
  wire __1595__;
  wire __1596__;
  wire __1597__;
  wire __1598__;
  wire __1599__;
  wire __1600__;
  wire __1601__;
  wire __1602__;
  wire __1603__;
  wire __1604__;
  wire __1605__;
  wire __1606__;
  wire __1607__;
  wire __1608__;
  wire __1609__;
  wire __1610__;
  wire __1611__;
  wire __1612__;
  wire __1613__;
  wire __1614__;
  wire __1615__;
  wire __1616__;
  wire __1617__;
  wire __1618__;
  wire __1619__;
  wire __1620__;
  wire __1621__;
  wire __1622__;
  wire __1623__;
  wire __1624__;
  wire __1625__;
  wire __1626__;
  wire __1627__;
  wire __1628__;
  wire __1629__;
  wire __1630__;
  wire __1631__;
  wire __1632__;
  wire __1633__;
  wire __1634__;
  wire __1635__;
  wire __1636__;
  wire __1637__;
  wire __1638__;
  wire __1639__;
  wire __1640__;
  wire __1641__;
  wire __1642__;
  wire __1643__;
  wire __1644__;
  wire __1645__;
  wire __1646__;
  wire __1647__;
  wire __1648__;
  wire __1649__;
  wire __1650__;
  wire __1651__;
  wire __1652__;
  wire __1653__;
  wire __1654__;
  wire __1655__;
  wire __1656__;
  wire __1657__;
  wire __1658__;
  wire __1659__;
  wire __1660__;
  wire __1661__;
  wire __1662__;
  wire __1663__;
  wire __1664__;
  wire __1665__;
  wire __1666__;
  wire __1667__;
  wire __1668__;
  wire __1669__;
  wire __1670__;
  wire __1671__;
  wire __1672__;
  wire __1673__;
  wire __1674__;
  wire __1675__;
  wire __1676__;
  wire __1677__;
  wire __1678__;
  wire __1679__;
  wire __1680__;
  wire __1681__;
  wire __1682__;
  wire __1683__;
  wire __1684__;
  wire __1685__;
  wire __1686__;
  wire __1687__;
  wire __1688__;
  wire __1689__;
  wire __1690__;
  wire __1691__;
  wire __1692__;
  wire __1693__;
  wire __1694__;
  wire __1695__;
  wire __1696__;
  wire __1697__;
  wire __1698__;
  wire __1699__;
  wire __1700__;
  wire __1701__;
  wire __1702__;
  wire __1703__;
  wire __1704__;
  wire __1705__;
  wire __1706__;
  wire __1707__;
  wire __1708__;
  wire __1709__;
  wire __1710__;
  wire __1711__;
  wire __1712__;
  wire __1713__;
  wire __1714__;
  wire __1715__;
  wire __1716__;
  wire __1717__;
  wire __1718__;
  wire __1719__;
  wire __1720__;
  wire __1721__;
  wire __1722__;
  wire __1723__;
  wire __1724__;
  wire __1725__;
  wire __1726__;
  wire __1727__;
  wire __1730__;
  wire __1731__;
  wire __1732__;
  wire __1733__;
  wire __1734__;
  wire __1735__;
  wire __1736__;
  wire __1737__;
  wire __1738__;
  wire __1739__;
  wire __1740__;
  wire __1741__;
  wire __1742__;
  wire __1743__;
  wire __1744__;
  wire __1745__;
  wire __1746__;
  wire __1747__;
  wire __1748__;
  wire __1749__;
  wire __1750__;
  wire __1751__;
  wire __1752__;
  wire __1753__;
  wire __1754__;
  wire __1755__;
  wire __1756__;
  wire __1757__;
  wire __1758__;
  wire __1759__;
  wire __1760__;
  wire __1761__;
  wire __1762__;
  wire __1763__;
  wire __1764__;
  wire __1765__;
  wire __1766__;
  wire __1767__;
  wire __1768__;
  wire __1769__;
  wire __1770__;
  wire __1771__;
  wire __1772__;
  wire __1773__;
  wire __1774__;
  wire __1775__;
  wire __1776__;
  wire __1777__;
  wire __1778__;
  wire __1779__;
  wire __1780__;
  wire __1781__;
  wire __1782__;
  wire __1783__;
  wire __1784__;
  wire __1785__;
  wire __1786__;
  wire __1787__;
  wire __1788__;
  wire __1789__;
  wire __1790__;
  wire __1791__;
  wire __1792__;
  wire __1793__;
  wire __1794__;
  wire __1795__;
  wire __1796__;
  wire __1797__;
  wire __1798__;
  wire __1799__;
  wire __1800__;
  wire __1801__;
  wire __1802__;
  wire __1803__;
  wire __1804__;
  wire __1805__;
  wire __1806__;
  wire __1807__;
  wire __1808__;
  wire __1809__;
  wire __1810__;
  wire __1811__;
  wire __1812__;
  wire __1813__;
  wire __1814__;
  wire __1815__;
  wire __1816__;
  wire __1817__;
  wire __1818__;
  wire __1819__;
  wire __1820__;
  wire __1821__;
  wire __1822__;
  wire __1823__;
  wire __1824__;
  wire __1825__;
  wire __1826__;
  wire __1827__;
  wire __1828__;
  wire __1829__;
  wire __1830__;
  wire __1831__;
  wire __1832__;
  wire __1833__;
  wire __1834__;
  wire __1835__;
  wire __1836__;
  wire __1837__;
  wire __1838__;
  wire __1839__;
  wire __1840__;
  wire __1841__;
  wire __1842__;
  wire __1843__;
  wire __1844__;
  wire __1845__;
  wire __1846__;
  wire __1847__;
  wire __1848__;
  wire __1849__;
  wire __1850__;
  wire __1851__;
  wire __1852__;
  wire __1853__;
  wire __1854__;
  wire __1855__;
  wire __1856__;
  wire __1857__;
  wire __1858__;
  wire __1859__;
  wire __1860__;
  wire __1861__;
  wire __1862__;
  wire __1863__;
  wire __1864__;
  wire __1865__;
  wire __1866__;
  wire __1867__;
  wire __1868__;
  wire __1869__;
  wire __1870__;
  wire __1871__;
  wire __1872__;
  wire __1873__;
  wire __1874__;
  wire __1875__;
  wire __1876__;
  wire __1877__;
  wire __1878__;
  wire __1879__;
  wire __1880__;
  wire __1881__;
  wire __1882__;
  wire __1883__;
  wire __1884__;
  wire __1885__;
  wire __1886__;
  wire __1887__;
  wire __1888__;
  wire __1889__;
  wire __1890__;
  wire __1891__;
  wire __1892__;
  wire __1893__;
  wire __1894__;
  wire __1895__;
  wire __1896__;
  wire __1897__;
  wire __1898__;
  wire __1899__;
  wire __1900__;
  wire __1901__;
  wire __1902__;
  wire __1903__;
  wire __1904__;
  wire __1905__;
  wire __1906__;
  wire __1907__;
  wire __1908__;
  wire __1909__;
  wire __1910__;
  wire __1911__;
  wire __1912__;
  wire __1913__;
  wire __1914__;
  wire __1915__;
  wire __1916__;
  wire __1917__;
  wire __1918__;
  wire __1919__;
  wire __1920__;
  wire __1921__;
  wire __1922__;
  wire __1923__;
  wire __1924__;
  wire __1925__;
  wire __1926__;
  wire __1927__;
  wire __1928__;
  wire __1929__;
  wire __1930__;
  wire __1931__;
  wire __1932__;
  wire __1933__;
  wire __1934__;
  wire __1935__;
  wire __1936__;
  wire __1937__;
  wire __1938__;
  wire __1939__;
  wire __1940__;
  wire __1941__;
  wire __1942__;
  wire __1943__;
  wire __1944__;
  wire __1945__;
  wire __1946__;
  wire __1947__;
  wire __1948__;
  wire __1949__;
  wire __1950__;
  wire __1951__;
  wire __1952__;
  wire __1953__;
  wire __1954__;
  wire __1955__;
  wire __1956__;
  wire __1957__;
  wire __1958__;
  wire __1959__;
  wire __1960__;
  wire __1961__;
  wire __1962__;
  wire __1963__;
  wire __1964__;
  wire __1965__;
  wire __1966__;
  wire __1967__;
  wire __1968__;
  wire __1969__;
  wire __1970__;
  wire __1971__;
  wire __1972__;
  wire __1973__;
  wire __1974__;
  wire __1975__;
  wire __1976__;
  wire __1977__;
  wire __1978__;
  wire __1979__;
  wire __1980__;
  wire __1981__;
  wire __1982__;
  wire __1983__;
  wire __1984__;
  wire __1985__;
  wire __1986__;
  wire __1987__;
  wire __1988__;
  wire __1989__;
  wire __1990__;
  wire __1991__;
  wire __1992__;
  wire __1993__;
  wire __1994__;
  wire __1995__;
  wire __1996__;
  wire __1997__;
  wire __1998__;
  wire __1999__;
  wire __2000__;
  wire __2001__;
  wire __2002__;
  wire __2003__;
  wire __2004__;
  wire __2005__;
  wire __2006__;
  wire __2007__;
  wire __2008__;
  wire __2009__;
  wire __2010__;
  wire __2011__;
  wire __2012__;
  wire __2013__;
  wire __2014__;
  wire __2015__;
  wire __2016__;
  wire __2017__;
  wire __2018__;
  wire __2019__;
  wire __2020__;
  wire __2021__;
  wire __2022__;
  wire __2023__;
  wire __2024__;
  wire __2025__;
  wire __2026__;
  wire __2027__;
  wire __2028__;
  wire __2029__;
  wire __2030__;
  wire __2031__;
  wire __2032__;
  wire __2033__;
  wire __2034__;
  wire __2035__;
  wire __2036__;
  wire __2037__;
  wire __2038__;
  wire __2039__;
  wire __2040__;
  wire __2041__;
  wire __2042__;
  wire __2043__;
  wire __2044__;
  wire __2045__;
  wire __2046__;
  wire __2047__;
  wire __2048__;
  wire __2049__;
  wire __2050__;
  wire __2051__;
  wire __2052__;
  wire __2053__;
  wire __2054__;
  wire __2055__;
  wire __2056__;
  wire __2057__;
  wire __2058__;
  wire __2059__;
  wire __2060__;
  wire __2061__;
  wire __2062__;
  wire __2063__;
  wire __2064__;
  wire __2065__;
  wire __2066__;
  wire __2067__;
  wire __2068__;
  wire __2069__;
  wire __2070__;
  wire __2071__;
  wire __2072__;
  wire __2073__;
  wire __2074__;
  wire __2075__;
  wire __2076__;
  wire __2077__;
  wire __2078__;
  wire __2079__;
  wire __2080__;
  wire __2081__;
  wire __2082__;
  wire __2083__;
  wire __2084__;
  wire __2085__;
  wire __2086__;
  wire __2087__;
  wire __2088__;
  wire __2089__;
  wire __2090__;
  wire __2091__;
  wire __2092__;
  wire __2093__;
  wire __2094__;
  wire __2095__;
  wire __2096__;
  wire __2097__;
  wire __2098__;
  wire __2099__;
  wire __2100__;
  wire __2101__;
  wire __2102__;
  wire __2103__;
  wire __2104__;
  wire __2105__;
  wire __2106__;
  wire __2107__;
  wire __2108__;
  wire __2109__;
  wire __2110__;
  wire __2111__;
  wire __2112__;
  wire __2113__;
  wire __2114__;
  wire __2115__;
  wire __2116__;
  wire __2117__;
  wire __2118__;
  wire __2119__;
  wire __2120__;
  wire __2121__;
  wire __2122__;
  wire __2123__;
  wire __2124__;
  wire __2125__;
  wire __2126__;
  wire __2127__;
  wire __2128__;
  wire __2129__;
  wire __2130__;
  wire __2131__;
  wire __2132__;
  wire __2133__;
  wire __2134__;
  wire __2135__;
  wire __2136__;
  wire __2137__;
  wire __2138__;
  wire __2139__;
  wire __2140__;
  wire __2141__;
  wire __2142__;
  wire __2143__;
  wire __2144__;
  wire __2145__;
  wire __2146__;
  wire __2147__;
  wire __2148__;
  wire __2149__;
  wire __2150__;
  wire __2151__;
  wire __2152__;
  wire __2153__;
  wire __2154__;
  wire __2155__;
  wire __2156__;
  wire __2157__;
  wire __2158__;
  wire __2159__;
  wire __2160__;
  wire __2161__;
  wire __2162__;
  wire __2163__;
  wire __2164__;
  wire __2165__;
  wire __2166__;
  wire __2167__;
  wire __2168__;
  wire __2169__;
  wire __2170__;
  wire __2171__;
  wire __2172__;
  wire __2173__;
  wire __2174__;
  wire __2175__;
  wire __2176__;
  wire __2177__;
  wire __2178__;
  wire __2179__;
  wire __2180__;
  wire __2181__;
  wire __2182__;
  wire __2183__;
  wire __2184__;
  wire __2185__;
  wire __2186__;
  wire __2187__;
  wire __2188__;
  wire __2189__;
  wire __2190__;
  wire __2191__;
  wire __2192__;
  wire __2193__;
  wire __2194__;
  wire __2195__;
  wire __2196__;
  wire __2197__;
  wire __2198__;
  wire __2199__;
  wire __2200__;
  wire __2201__;
  wire __2202__;
  wire __2203__;
  wire __2204__;
  wire __2205__;
  wire __2206__;
  wire __2207__;
  wire __2208__;
  wire __2209__;
  wire __2210__;
  wire __2211__;
  wire __2212__;
  wire __2213__;
  wire __2214__;
  wire __2215__;
  wire __2216__;
  wire __2217__;
  wire __2218__;
  wire __2219__;
  wire __2220__;
  wire __2221__;
  wire __2222__;
  wire __2223__;
  wire __2224__;
  wire __2225__;
  wire __2226__;
  wire __2227__;
  wire __2228__;
  wire __2229__;
  wire __2230__;
  wire __2231__;
  wire __2232__;
  wire __2233__;
  wire __2234__;
  wire __2235__;
  wire __2236__;
  wire __2237__;
  wire __2238__;
  wire __2239__;
  wire __2240__;
  wire __2241__;
  wire __2242__;
  wire __2243__;
  wire __2244__;
  wire __2245__;
  wire __2246__;
  wire __2247__;
  wire __2248__;
  wire __2249__;
  wire __2250__;
  wire __2251__;
  wire __2252__;
  wire __2253__;
  wire __2254__;
  wire __2255__;
  wire __2256__;
  wire __2257__;
  wire __2258__;
  wire __2259__;
  wire __2260__;
  wire __2261__;
  wire __2262__;
  wire __2263__;
  wire __2264__;
  wire __2265__;
  wire __2266__;
  wire __2267__;
  wire __2268__;
  wire __2269__;
  wire __2270__;
  wire __2271__;
  wire __2272__;
  wire __2273__;
  wire __2274__;
  wire __2275__;
  wire __2276__;
  wire __2277__;
  wire __2278__;
  wire __2279__;
  wire __2280__;
  wire __2281__;
  wire __2282__;
  wire __2283__;
  wire __2284__;
  wire __2285__;
  wire __2286__;
  wire __2287__;
  wire __2288__;
  wire __2289__;
  wire __2290__;
  wire __2291__;
  wire __2292__;
  wire __2293__;
  wire __2294__;
  wire __2295__;
  wire __2296__;
  wire __2297__;
  wire __2298__;
  wire __2299__;
  wire __2300__;
  wire __2301__;
  wire __2302__;
  wire __2303__;
  wire __2304__;
  wire __2305__;
  wire __2306__;
  wire __2307__;
  wire __2308__;
  wire __2309__;
  wire __2310__;
  wire __2311__;
  wire __2312__;
  wire __2313__;
  wire __2314__;
  wire __2315__;
  wire __2316__;
  wire __2317__;
  wire __2318__;
  wire __2319__;
  wire __2320__;
  wire __2321__;
  wire __2322__;
  wire __2323__;
  wire __2324__;
  wire __2325__;
  wire __2326__;
  wire __2327__;
  wire __2328__;
  wire __2329__;
  wire __2330__;
  wire __2331__;
  wire __2332__;
  wire __2333__;
  wire __2334__;
  wire __2335__;
  wire __2336__;
  wire __2337__;
  wire __2338__;
  wire __2339__;
  wire __2340__;
  wire __2341__;
  wire __2342__;
  wire __2343__;
  wire __2344__;
  wire __2345__;
  wire __2346__;
  wire __2347__;
  wire __2348__;
  wire __2349__;
  wire __2350__;
  wire __2351__;
  wire __2352__;
  wire __2353__;
  wire __2354__;
  wire __2355__;
  wire __2356__;
  wire __2357__;
  wire __2358__;
  wire __2359__;
  wire __2360__;
  wire __2361__;
  wire __2362__;
  wire __2363__;
  wire __2364__;
  wire __2365__;
  wire __2366__;
  wire __2367__;
  wire __2368__;
  wire __2369__;
  wire __2370__;
  wire __2371__;
  wire __2372__;
  wire __2373__;
  wire __2374__;
  wire __2375__;
  wire __2376__;
  wire __2377__;
  wire __2378__;
  wire __2379__;
  wire __2380__;
  wire __2381__;
  wire __2382__;
  wire __2383__;
  wire __2384__;
  wire __2385__;
  wire __2386__;
  wire __2387__;
  wire __2388__;
  wire __2389__;
  wire __2390__;
  wire __2391__;
  wire __2392__;
  wire __2393__;
  wire __2394__;
  wire __2395__;
  wire __2396__;
  wire __2397__;
  wire __2398__;
  wire __2399__;
  wire __2400__;
  wire __2401__;
  wire __2402__;
  wire __2403__;
  wire __2404__;
  wire __2405__;
  wire __2406__;
  wire __2407__;
  wire __2408__;
  wire __2409__;
  wire __2410__;
  wire __2411__;
  wire __2412__;
  wire __2413__;
  wire __2414__;
  wire __2415__;
  wire __2416__;
  wire __2417__;
  wire __2418__;
  wire __2419__;
  wire __2420__;
  wire __2421__;
  wire __2422__;
  wire __2423__;
  wire __2424__;
  wire __2425__;
  wire __2426__;
  wire __2427__;
  wire __2428__;
  wire __2429__;
  wire __2430__;
  wire __2431__;
  wire __2432__;
  wire __2433__;
  wire __2434__;
  wire __2435__;
  wire __2436__;
  wire __2437__;
  wire __2438__;
  wire __2439__;
  wire __2440__;
  wire __2441__;
  wire __2442__;
  wire __2443__;
  wire __2444__;
  wire __2445__;
  wire __2446__;
  wire __2447__;
  wire __2448__;
  wire __2449__;
  wire __2450__;
  wire __2451__;
  wire __2452__;
  wire __2453__;
  wire __2454__;
  wire __2455__;
  wire __2456__;
  wire __2457__;
  wire __2458__;
  wire __2459__;
  wire __2460__;
  wire __2461__;
  wire __2462__;
  wire __2463__;
  wire __2464__;
  wire __2465__;
  wire __2466__;
  wire __2467__;
  wire __2468__;
  wire __2469__;
  wire __2470__;
  wire __2471__;
  wire __2472__;
  wire __2473__;
  wire __2474__;
  wire __2475__;
  wire __2476__;
  wire __2477__;
  wire __2478__;
  wire __2479__;
  wire __2480__;
  wire __2481__;
  wire __2482__;
  wire __2483__;
  wire __2484__;
  wire __2485__;
  wire __2486__;
  wire __2487__;
  wire __2488__;
  wire __2489__;
  wire __2490__;
  wire __2491__;
  wire __2492__;
  wire __2493__;
  wire __2494__;
  wire __2495__;
  wire __2496__;
  wire __2497__;
  wire __2498__;
  wire __2499__;
  wire __2500__;
  wire __2501__;
  wire __2502__;
  wire __2503__;
  wire __2504__;
  wire __2505__;
  wire __2506__;
  wire __2507__;
  wire __2508__;
  wire __2509__;
  wire __2510__;
  wire __2511__;
  wire __2512__;
  wire __2513__;
  wire __2514__;
  wire __2515__;
  wire __2516__;
  wire __2517__;
  wire __2518__;
  wire __2519__;
  wire __2520__;
  wire __2521__;
  wire __2522__;
  wire __2523__;
  wire __2524__;
  wire __2525__;
  wire __2526__;
  wire __2527__;
  wire __2528__;
  wire __2529__;
  wire __2530__;
  wire __2531__;
  wire __2532__;
  wire __2533__;
  wire __2534__;
  wire __2535__;
  wire __2536__;
  wire __2537__;
  wire __2538__;
  wire __2539__;
  wire __2540__;
  wire __2541__;
  wire __2542__;
  wire __2543__;
  wire __2544__;
  wire __2545__;
  wire __2546__;
  wire __2547__;
  wire __2548__;
  wire __2549__;
  wire __2550__;
  wire __2551__;
  wire __2552__;
  wire __2553__;
  wire __2554__;
  wire __2555__;
  wire __2556__;
  wire __2557__;
  wire __2558__;
  wire __2559__;
  wire __2560__;
  wire __2561__;
  wire __2562__;
  wire __2563__;
  wire __2564__;
  wire __2565__;
  wire __2566__;
  wire __2567__;
  wire __2568__;
  wire __2569__;
  wire __2570__;
  wire __2571__;
  wire __2572__;
  wire __2573__;
  wire __2574__;
  wire __2575__;
  wire __2576__;
  wire __2577__;
  wire __2578__;
  wire __2579__;
  wire __2580__;
  wire __2581__;
  wire __2582__;
  wire __2583__;
  wire __2584__;
  wire __2585__;
  wire __2586__;
  wire __2587__;
  wire __2588__;
  wire __2589__;
  wire __2590__;
  wire __2591__;
  wire __2592__;
  wire __2593__;
  wire __2594__;
  wire __2595__;
  wire __2596__;
  wire __2597__;
  wire __2598__;
  wire __2599__;
  wire __2600__;
  wire __2601__;
  wire __2602__;
  wire __2603__;
  wire __2604__;
  wire __2605__;
  wire __2606__;
  wire __2607__;
  wire __2608__;
  wire __2609__;
  wire __2610__;
  wire __2611__;
  wire __2612__;
  wire __2613__;
  wire __2614__;
  wire __2615__;
  wire __2616__;
  wire __2617__;
  wire __2618__;
  wire __2619__;
  wire __2620__;
  wire __2621__;
  wire __2622__;
  wire __2623__;
  wire __2624__;
  wire __2625__;
  wire __2626__;
  wire __2627__;
  wire __2628__;
  wire __2629__;
  wire __2630__;
  wire __2631__;
  wire __2632__;
  wire __2633__;
  wire __2634__;
  wire __2635__;
  wire __2636__;
  wire __2637__;
  wire __2638__;
  wire __2639__;
  wire __2640__;
  wire __2641__;
  wire __2642__;
  wire __2643__;
  wire __2644__;
  wire __2645__;
  wire __2646__;
  wire __2647__;
  wire __2648__;
  wire __2649__;
  wire __2650__;
  wire __2651__;
  wire __2652__;
  wire __2653__;
  wire __2654__;
  wire __2655__;
  wire __2656__;
  wire __2657__;
  wire __2658__;
  wire __2659__;
  wire __2660__;
  wire __2661__;
  wire __2662__;
  wire __2663__;
  wire __2664__;
  wire __2665__;
  wire __2666__;
  wire __2667__;
  wire __2668__;
  wire __2669__;
  wire __2670__;
  wire __2671__;
  wire __2672__;
  wire __2673__;
  wire __2674__;
  wire __2675__;
  wire __2676__;
  wire __2677__;
  wire __2678__;
  wire __2679__;
  wire __2680__;
  wire __2681__;
  wire __2682__;
  wire __2683__;
  wire __2684__;
  wire __2685__;
  wire __2686__;
  wire __2687__;
  wire __2688__;
  wire __2689__;
  wire __2690__;
  wire __2691__;
  wire __2692__;
  wire __2693__;
  wire __2694__;
  wire __2695__;
  wire __2696__;
  wire __2697__;
  wire __2698__;
  wire __2699__;
  wire __2700__;
  wire __2701__;
  wire __2702__;
  wire __2703__;
  wire __2704__;
  wire __2705__;
  wire __2706__;
  wire __2707__;
  wire __2708__;
  wire __2709__;
  wire __2710__;
  wire __2711__;
  wire __2712__;
  wire __2713__;
  wire __2714__;
  wire __2715__;
  wire __2716__;
  wire __2717__;
  wire __2718__;
  wire __2719__;
  wire __2720__;
  wire __2721__;
  wire __2722__;
  wire __2723__;
  wire __2724__;
  wire __2725__;
  wire __2726__;
  wire __2727__;
  wire __2728__;
  wire __2729__;
  wire __2730__;
  wire __2731__;
  wire __2732__;
  wire __2733__;
  wire __2734__;
  wire __2735__;
  wire __2736__;
  wire __2737__;
  wire __2738__;
  wire __2739__;
  wire __2740__;
  wire __2741__;
  wire __2742__;
  wire __2743__;
  wire __2744__;
  wire __2745__;
  wire __2746__;
  wire __2747__;
  wire __2748__;
  wire __2749__;
  wire __2750__;
  wire __2751__;
  wire __2752__;
  wire __2753__;
  wire __2754__;
  wire __2755__;
  wire __2756__;
  wire __2757__;
  wire __2758__;
  wire __2759__;
  wire __2760__;
  wire __2761__;
  wire __2762__;
  wire __2763__;
  wire __2764__;
  wire __2765__;
  wire __2766__;
  wire __2767__;
  wire __2768__;
  wire __2769__;
  wire __2770__;
  wire __2771__;
  wire __2772__;
  wire __2773__;
  wire __2774__;
  wire __2775__;
  wire __2776__;
  wire __2777__;
  wire __2778__;
  wire __2779__;
  wire __2780__;
  wire __2781__;
  wire __2782__;
  wire __2783__;
  wire __2784__;
  wire __2785__;
  wire __2786__;
  wire __2787__;
  wire __2788__;
  wire __2789__;
  wire __2790__;
  wire __2791__;
  wire __2792__;
  wire __2793__;
  wire __2794__;
  wire __2795__;
  wire __2796__;
  wire __2797__;
  wire __2798__;
  wire __2799__;
  wire __2800__;
  wire __2801__;
  wire __2802__;
  wire __2803__;
  wire __2804__;
  wire __2805__;
  wire __2806__;
  wire __2807__;
  wire __2808__;
  wire __2809__;
  wire __2810__;
  wire __2811__;
  wire __2812__;
  wire __2813__;
  wire __2814__;
  wire __2815__;
  wire __2816__;
  wire __2817__;
  wire __2818__;
  wire __2819__;
  wire __2820__;
  wire __2821__;
  wire __2822__;
  wire __2823__;
  wire __2824__;
  wire __2825__;
  wire __2826__;
  wire __2827__;
  wire __2828__;
  wire __2829__;
  wire __2830__;
  wire __2831__;
  wire __2832__;
  wire __2833__;
  wire __2834__;
  wire __2835__;
  wire __2836__;
  wire __2837__;
  wire __2838__;
  wire __2839__;
  wire __2840__;
  wire __2841__;
  wire __2842__;
  wire __2843__;
  wire __2844__;
  wire __2845__;
  wire __2846__;
  wire __2847__;
  wire __2848__;
  wire __2849__;
  wire __2850__;
  wire __2851__;
  wire __2852__;
  wire __2853__;
  wire __2854__;
  wire __2855__;
  wire __2856__;
  wire __2857__;
  wire __2858__;
  wire __2859__;
  wire __2860__;
  wire __2861__;
  wire __2862__;
  wire __2863__;
  wire __2864__;
  wire __2865__;
  wire __2866__;
  wire __2867__;
  wire __2868__;
  wire __2869__;
  wire __2870__;
  wire __2871__;
  wire __2872__;
  wire __2873__;
  wire __2874__;
  wire __2875__;
  wire __2876__;
  wire __2877__;
  wire __2878__;
  wire __2879__;
  wire __2880__;
  wire __2881__;
  wire __2882__;
  wire __2883__;
  wire __2884__;
  wire __2885__;
  wire __2886__;
  wire __2887__;
  wire __2888__;
  wire __2889__;
  wire __2890__;
  wire __2891__;
  wire __2892__;
  wire __2893__;
  wire __2894__;
  wire __2895__;
  wire __2896__;
  wire __2897__;
  wire __2898__;
  wire __2899__;
  wire __2900__;
  wire __2901__;
  wire __2902__;
  wire __2903__;
  wire __2904__;
  wire __2905__;
  wire __2906__;
  wire __2907__;
  wire __2908__;
  wire __2909__;
  wire __2910__;
  wire __2911__;
  wire __2912__;
  wire __2913__;
  wire __2914__;
  wire __2915__;
  wire __2916__;
  wire __2917__;
  wire __2918__;
  wire __2919__;
  wire __2920__;
  wire __2921__;
  wire __2922__;
  wire __2923__;
  wire __2924__;
  wire __2925__;
  wire __2926__;
  wire __2927__;
  wire __2928__;
  wire __2929__;
  wire __2930__;
  wire __2931__;
  wire __2932__;
  wire __2933__;
  wire __2934__;
  wire __2935__;
  wire __2936__;
  wire __2937__;
  wire __2938__;
  wire __2939__;
  wire __2940__;
  wire __2941__;
  wire __2942__;
  wire __2943__;
  wire __2944__;
  wire __2945__;
  wire __2946__;
  wire __2947__;
  wire __2948__;
  wire __2949__;
  wire __2950__;
  wire __2951__;
  wire __2952__;
  wire __2953__;
  wire __2954__;
  wire __2955__;
  wire __2956__;
  wire __2957__;
  wire __2958__;
  wire __2959__;
  wire __2960__;
  wire __2961__;
  wire __2962__;
  wire __2963__;
  wire __2964__;
  wire __2965__;
  wire __2966__;
  wire __2967__;
  wire __2968__;
  wire __2969__;
  wire __2970__;
  wire __2971__;
  wire __2972__;
  wire __2973__;
  wire __2974__;
  wire __2975__;
  wire __2976__;
  wire __2977__;
  wire __2978__;
  wire __2979__;
  wire __2980__;
  wire __2981__;
  wire __2982__;
  wire __2983__;
  wire __2984__;
  wire __2985__;
  wire __2986__;
  wire __2987__;
  wire __2988__;
  wire __2989__;
  wire __2990__;
  wire __2991__;
  wire __2992__;
  wire __2993__;
  wire __2994__;
  wire __2995__;
  wire __2996__;
  wire __2997__;
  wire __2998__;
  wire __2999__;
  wire __3000__;
  wire __3001__;
  wire __3002__;
  wire __3003__;
  wire __3004__;
  wire __3005__;
  wire __3006__;
  wire __3007__;
  wire __3008__;
  wire __3009__;
  wire __3010__;
  wire __3011__;
  wire __3012__;
  wire __3013__;
  wire __3014__;
  wire __3015__;
  wire __3016__;
  wire __3017__;
  wire __3018__;
  wire __3019__;
  wire __3020__;
  wire __3021__;
  wire __3022__;
  wire __3023__;
  wire __3024__;
  wire __3025__;
  wire __3026__;
  wire __3027__;
  wire __3028__;
  wire __3029__;
  wire __3030__;
  wire __3031__;
  wire __3032__;
  wire __3033__;
  wire __3034__;
  wire __3035__;
  wire __3036__;
  wire __3037__;
  wire __3038__;
  wire __3039__;
  wire __3040__;
  wire __3041__;
  wire __3042__;
  wire __3043__;
  wire __3044__;
  wire __3045__;
  wire __3046__;
  wire __3047__;
  wire __3048__;
  wire __3049__;
  wire __3050__;
  wire __3051__;
  wire __3052__;
  wire __3053__;
  wire __3054__;
  wire __3055__;
  wire __3056__;
  wire __3057__;
  wire __3058__;
  wire __3059__;
  wire __3060__;
  wire __3061__;
  wire __3062__;
  wire __3063__;
  wire __3064__;
  wire __3065__;
  wire __3066__;
  wire __3067__;
  wire __3068__;
  wire __3069__;
  wire __3070__;
  wire __3071__;
  wire __3072__;
  wire __3073__;
  wire __3074__;
  wire __3075__;
  wire __3076__;
  wire __3077__;
  wire __3078__;
  wire __3079__;
  wire __3080__;
  wire __3081__;
  wire __3082__;
  wire __3083__;
  wire __3084__;
  wire __3085__;
  wire __3086__;
  wire __3087__;
  wire __3088__;
  wire __3089__;
  wire __3090__;
  wire __3091__;
  wire __3092__;
  wire __3093__;
  wire __3094__;
  wire __3095__;
  wire __3096__;
  wire __3097__;
  wire __3098__;
  wire __3099__;
  wire __3100__;
  wire __3101__;
  wire __3102__;
  wire __3103__;
  wire __3104__;
  wire __3105__;
  wire __3106__;
  wire __3107__;
  wire __3108__;
  wire __3109__;
  wire __3110__;
  wire __3111__;
  wire __3112__;
  wire __3113__;
  wire __3114__;
  wire __3115__;
  wire __3116__;
  wire __3117__;
  wire __3118__;
  wire __3119__;
  wire __3120__;
  wire __3121__;
  wire __3122__;
  wire __3123__;
  wire __3124__;
  wire __3125__;
  wire __3126__;
  wire __3127__;
  wire __3128__;
  wire __3129__;
  wire __3130__;
  wire __3131__;
  wire __3132__;
  wire __3133__;
  wire __3134__;
  wire __3135__;
  wire __3136__;
  wire __3137__;
  wire __3138__;
  wire __3139__;
  wire __3140__;
  wire __3141__;
  wire __3142__;
  wire __3143__;
  wire __3144__;
  wire __3145__;
  wire __3146__;
  wire __3147__;
  wire __3148__;
  wire __3149__;
  wire __3150__;
  wire __3151__;
  wire __3152__;
  wire __3153__;
  wire __3154__;
  wire __3155__;
  wire __3156__;
  wire __3157__;
  wire __3158__;
  wire __3159__;
  wire __3160__;
  wire __3161__;
  wire __3162__;
  wire __3163__;
  wire __3164__;
  wire __3165__;
  wire __3166__;
  wire __3167__;
  wire __3168__;
  wire __3169__;
  wire __3170__;
  wire __3171__;
  wire __3172__;
  wire __3173__;
  wire __3174__;
  wire __3175__;
  wire __3176__;
  wire __3177__;
  wire __3178__;
  wire __3179__;
  wire __3180__;
  wire __3181__;
  wire __3182__;
  wire __3183__;
  wire __3184__;
  wire __3185__;
  wire __3186__;
  wire __3187__;
  wire __3188__;
  wire __3189__;
  wire __3190__;
  wire __3191__;
  wire __3192__;
  wire __3193__;
  wire __3194__;
  wire __3195__;
  wire __3196__;
  wire __3197__;
  wire __3198__;
  wire __3199__;
  wire __3200__;
  wire __3201__;
  wire __3202__;
  wire __3203__;
  wire __3204__;
  wire __3205__;
  wire __3206__;
  wire __3207__;
  wire __3208__;
  wire __3209__;
  wire __3210__;
  wire __3211__;
  wire __3212__;
  wire __3213__;
  wire __3214__;
  wire __3215__;
  wire __3216__;
  wire __3217__;
  wire __3218__;
  wire __3219__;
  wire __3220__;
  wire __3221__;
  wire __3222__;
  wire __3223__;
  wire __3224__;
  wire __3225__;
  wire __3226__;
  wire __3227__;
  wire __3228__;
  wire __3229__;
  wire __3230__;
  wire __3231__;
  wire __3232__;
  wire __3233__;
  wire __3234__;
  wire __3235__;
  wire __3236__;
  wire __3237__;
  wire __3238__;
  wire __3239__;
  wire __3240__;
  wire __3241__;
  wire __3242__;
  wire __3243__;
  wire __3244__;
  wire __3245__;
  wire __3246__;
  wire __3247__;
  wire __3248__;
  wire __3249__;
  wire __3250__;
  wire __3251__;
  wire __3252__;
  wire __3253__;
  wire __3254__;
  wire __3255__;
  wire __3256__;
  wire __3257__;
  wire __3258__;
  wire __3259__;
  wire __3260__;
  wire __3261__;
  wire __3262__;
  wire __3263__;
  wire __3264__;
  wire __3265__;
  wire __3266__;
  wire __3267__;
  wire __3268__;
  wire __3269__;
  wire __3270__;
  wire __3271__;
  wire __3272__;
  wire __3273__;
  wire __3274__;
  wire __3275__;
  wire __3276__;
  wire __3277__;
  wire __3278__;
  wire __3279__;
  wire __3280__;
  wire __3281__;
  wire __3282__;
  wire __3283__;
  wire __3284__;
  wire __3285__;
  wire __3286__;
  wire __3287__;
  wire __3288__;
  wire __3289__;
  wire __3290__;
  wire __3291__;
  wire __3292__;
  wire __3293__;
  wire __3294__;
  wire __3295__;
  wire __3296__;
  wire __3297__;
  wire __3298__;
  wire __3299__;
  wire __3300__;
  wire __3301__;
  wire __3302__;
  wire __3303__;
  wire __3304__;
  wire __3305__;
  wire __3306__;
  wire __3307__;
  wire __3308__;
  wire __3309__;
  wire __3310__;
  wire __3311__;
  wire __3312__;
  wire __3313__;
  wire __3314__;
  wire __3315__;
  wire __3316__;
  wire __3317__;
  wire __3318__;
  wire __3319__;
  wire __3320__;
  wire __3321__;
  wire __3322__;
  wire __3323__;
  wire __3324__;
  wire __3325__;
  wire __3326__;
  wire __3327__;
  wire __3328__;
  wire __3329__;
  wire __3330__;
  wire __3331__;
  wire __3332__;
  wire __3333__;
  wire __3334__;
  wire __3335__;
  wire __3336__;
  wire __3337__;
  wire __3338__;
  wire __3339__;
  wire __3340__;
  wire __3341__;
  wire __3342__;
  wire __3343__;
  wire __3344__;
  wire __3345__;
  wire __3346__;
  wire __3347__;
  wire __3348__;
  wire __3349__;
  wire __3350__;
  wire __3351__;
  wire __3352__;
  wire __3353__;
  wire __3354__;
  wire __3355__;
  wire __3356__;
  wire __3357__;
  wire __3358__;
  wire __3359__;
  wire __3360__;
  wire __3361__;
  wire __3362__;
  wire __3363__;
  wire __3364__;
  wire __3365__;
  wire __3366__;
  wire __3367__;
  wire __3368__;
  wire __3369__;
  wire __3370__;
  wire __3371__;
  wire __3372__;
  wire __3373__;
  wire __3374__;
  wire __3375__;
  wire __3376__;
  wire __3377__;
  wire __3378__;
  wire __3379__;
  wire __3380__;
  wire __3381__;
  wire __3382__;
  wire __3383__;
  wire __3384__;
  wire __3385__;
  wire __3386__;
  wire __3387__;
  wire __3388__;
  wire __3389__;
  wire __3390__;
  wire __3391__;
  wire __3392__;
  wire __3393__;
  wire __3394__;
  wire __3395__;
  wire __3396__;
  wire __3397__;
  wire __3398__;
  wire __3399__;
  wire __3400__;
  wire __3401__;
  wire __3402__;
  wire __3403__;
  wire __3404__;
  wire __3405__;
  wire __3406__;
  wire __3407__;
  wire __3408__;
  wire __3409__;
  wire __3410__;
  wire __3411__;
  wire __3412__;
  wire __3413__;
  wire __3414__;
  wire __3415__;
  wire __3416__;
  wire __3417__;
  wire __3418__;
  wire __3419__;
  wire __3420__;
  wire __3421__;
  wire __3422__;
  wire __3423__;
  wire __3424__;
  wire __3425__;
  wire __3426__;
  wire __3427__;
  wire __3428__;
  wire __3429__;
  wire __3430__;
  wire __3431__;
  wire __3432__;
  wire __3433__;
  wire __3434__;
  wire __3435__;
  wire __3436__;
  wire __3437__;
  wire __3438__;
  wire __3439__;
  wire __3440__;
  wire __3441__;
  wire __3442__;
  wire __3443__;
  wire __3444__;
  wire __3445__;
  wire __3446__;
  wire __3447__;
  wire __3448__;
  wire __3449__;
  wire __3450__;
  wire __3451__;
  wire __3452__;
  wire __3453__;
  wire __3454__;
  wire __3455__;
  wire __3456__;
  wire __3457__;
  wire __3458__;
  wire __3459__;
  wire __3460__;
  wire __3461__;
  wire __3462__;
  wire __3463__;
  wire __3464__;
  wire __3465__;
  wire __3466__;
  wire __3467__;
  wire __3468__;
  wire __3469__;
  wire __3470__;
  wire __3471__;
  wire __3472__;
  wire __3473__;
  wire __3474__;
  wire __3475__;
  wire __3476__;
  wire __3477__;
  wire __3478__;
  wire __3479__;
  wire __3480__;
  wire __3481__;
  wire __3482__;
  wire __3483__;
  wire __3484__;
  wire __3485__;
  wire __3486__;
  wire __3487__;
  wire __3488__;
  wire __3489__;
  wire __3490__;
  wire __3491__;
  wire __3492__;
  wire __3493__;
  wire __3494__;
  wire __3495__;
  wire __3496__;
  wire __3497__;
  wire __3498__;
  wire __3499__;
  wire __3500__;
  wire __3501__;
  wire __3502__;
  wire __3503__;
  wire __3504__;
  wire __3505__;
  wire __3506__;
  wire __3507__;
  wire __3508__;
  wire __3509__;
  wire __3510__;
  wire __3511__;
  wire __3512__;
  wire __3513__;
  wire __3514__;
  wire __3515__;
  wire __3516__;
  wire __3517__;
  wire __3518__;
  wire __3519__;
  wire __3520__;
  wire __3521__;
  wire __3522__;
  wire __3523__;
  wire __3524__;
  wire __3525__;
  wire __3526__;
  wire __3527__;
  wire __3528__;
  wire __3529__;
  wire __3530__;
  wire __3531__;
  wire __3532__;
  wire __3533__;
  wire __3534__;
  wire __3535__;
  wire __3536__;
  wire __3537__;
  wire __3538__;
  wire __3539__;
  wire __3540__;
  wire __3541__;
  wire __3542__;
  wire __3543__;
  wire __3544__;
  wire __3545__;
  wire __3546__;
  wire __3547__;
  wire __3548__;
  wire __3549__;
  wire __3550__;
  wire __3551__;
  wire __3552__;
  wire __3553__;
  wire __3554__;
  wire __3555__;
  wire __3556__;
  wire __3557__;
  wire __3558__;
  wire __3559__;
  wire __3560__;
  wire __3561__;
  wire __3562__;
  wire __3563__;
  wire __3564__;
  wire __3565__;
  wire __3566__;
  wire __3567__;
  wire __3568__;
  wire __3569__;
  wire __3570__;
  wire __3571__;
  wire __3572__;
  wire __3573__;
  wire __3574__;
  wire __3575__;
  wire __3576__;
  wire __3577__;
  wire __3578__;
  wire __3579__;
  wire __3580__;
  wire __3581__;
  wire __3582__;
  wire __3583__;
  wire __3584__;
  wire __3585__;
  wire __3586__;
  wire __3587__;
  wire __3588__;
  wire __3589__;
  wire __3590__;
  wire __3591__;
  wire __3592__;
  wire __3593__;
  wire __3594__;
  wire __3595__;
  wire __3596__;
  wire __3597__;
  wire __3598__;
  wire __3599__;
  wire __3600__;
  wire __3601__;
  wire __3602__;
  wire __3603__;
  wire __3604__;
  wire __3605__;
  wire __3606__;
  wire __3607__;
  wire __3608__;
  wire __3609__;
  wire __3610__;
  wire __3611__;
  wire __3612__;
  wire __3613__;
  wire __3614__;
  wire __3615__;
  wire __3616__;
  wire __3617__;
  wire __3618__;
  wire __3619__;
  wire __3620__;
  wire __3621__;
  wire __3622__;
  wire __3623__;
  wire __3624__;
  wire __3625__;
  wire __3626__;
  wire __3627__;
  wire __3628__;
  wire __3629__;
  wire __3630__;
  wire __3631__;
  wire __3632__;
  wire __3633__;
  wire __3634__;
  wire __3635__;
  wire __3636__;
  wire __3637__;
  wire __3638__;
  wire __3639__;
  wire __3640__;
  wire __3641__;
  wire __3642__;
  wire __3643__;
  wire __3644__;
  wire __3645__;
  wire __3646__;
  wire __3647__;
  wire __3648__;
  wire __3649__;
  wire __3650__;
  wire __3651__;
  wire __3652__;
  wire __3653__;
  wire __3654__;
  wire __3655__;
  wire __3656__;
  wire __3657__;
  wire __3658__;
  wire __3659__;
  wire __3660__;
  wire __3661__;
  wire __3662__;
  wire __3663__;
  wire __3664__;
  wire __3665__;
  wire __3666__;
  wire __3667__;
  wire __3668__;
  wire __3669__;
  wire __3670__;
  wire __3671__;
  wire __3672__;
  wire __3673__;
  wire __3674__;
  wire __3675__;
  wire __3676__;
  wire __3677__;
  wire __3678__;
  wire __3679__;
  wire __3680__;
  wire __3681__;
  wire __3682__;
  wire __3683__;
  wire __3684__;
  wire __3685__;
  wire __3686__;
  wire __3687__;
  wire __3688__;
  wire __3689__;
  wire __3690__;
  wire __3691__;
  wire __3692__;
  wire __3693__;
  wire __3694__;
  wire __3695__;
  wire __3696__;
  wire __3697__;
  wire __3698__;
  wire __3699__;
  wire __3700__;
  wire __3701__;
  wire __3702__;
  wire __3703__;
  wire __3704__;
  wire __3705__;
  wire __3706__;
  wire __3707__;
  wire __3708__;
  wire __3709__;
  wire __3710__;
  wire __3711__;
  wire __3712__;
  wire __3713__;
  wire __3714__;
  wire __3715__;
  wire __3716__;
  wire __3717__;
  wire __3718__;
  wire __3719__;
  wire __3720__;
  wire __3721__;
  wire __3722__;
  wire __3723__;
  wire __3724__;
  wire __3725__;
  wire __3726__;
  wire __3727__;
  wire __3728__;
  wire __3729__;
  wire __3730__;
  wire __3731__;
  wire __3732__;
  wire __3733__;
  wire __3734__;
  wire __3735__;
  wire __3736__;
  wire __3737__;
  wire __3738__;
  wire __3739__;
  wire __3740__;
  wire __3741__;
  wire __3742__;
  wire __3743__;
  wire __3744__;
  wire __3745__;
  wire __3746__;
  wire __3747__;
  wire __3748__;
  wire __3749__;
  wire __3750__;
  wire __3751__;
  wire __3752__;
  wire __3753__;
  wire __3754__;
  wire __3755__;
  wire __3756__;
  wire __3757__;
  wire __3758__;
  wire __3759__;
  wire __3760__;
  wire __3761__;
  wire __3762__;
  wire __3763__;
  wire __3764__;
  wire __3765__;
  wire __3766__;
  wire __3767__;
  wire __3768__;
  wire __3769__;
  wire __3770__;
  wire __3771__;
  wire __3772__;
  wire __3773__;
  wire __3774__;
  wire __3775__;
  wire __3776__;
  wire __3777__;
  wire __3778__;
  wire __3779__;
  wire __3780__;
  wire __3781__;
  wire __3782__;
  wire __3783__;
  wire __3784__;
  wire __3785__;
  wire __3786__;
  wire __3787__;
  wire __3788__;
  wire __3789__;
  wire __3790__;
  wire __3791__;
  wire __3792__;
  wire __3793__;
  wire __3794__;
  wire __3795__;
  wire __3796__;
  wire __3797__;
  wire __3798__;
  wire __3799__;
  wire __3800__;
  wire __3801__;
  wire __3802__;
  wire __3803__;
  wire __3804__;
  wire __3805__;
  wire __3806__;
  wire __3807__;
  wire __3808__;
  wire __3809__;
  wire __3810__;
  wire __3811__;
  wire __3812__;
  wire __3813__;
  wire __3814__;
  wire __3815__;
  wire __3816__;
  wire __3817__;
  wire __3818__;
  wire __3819__;
  wire __3820__;
  wire __3821__;
  wire __3822__;
  wire __3823__;
  wire __3824__;
  wire __3825__;
  wire __3826__;
  wire __3827__;
  wire __3828__;
  wire __3829__;
  wire __3830__;
  wire __3831__;
  wire __3832__;
  wire __3833__;
  wire __3834__;
  wire __3835__;
  wire __3836__;
  wire __3837__;
  wire __3838__;
  wire __3839__;
  wire __3840__;
  wire __3841__;
  wire __3842__;
  wire __3843__;
  wire __3844__;
  wire __3845__;
  wire __3846__;
  wire __3847__;
  wire __3848__;
  wire __3849__;
  wire __3850__;
  wire __3851__;
  wire __3852__;
  wire __3853__;
  wire __3854__;
  wire __3855__;
  wire __3856__;
  wire __3857__;
  wire __3858__;
  wire __3859__;
  wire __3860__;
  wire __3861__;
  wire __3862__;
  wire __3863__;
  wire __3864__;
  wire __3865__;
  wire __3866__;
  wire __3867__;
  wire __3868__;
  wire __3869__;
  wire __3870__;
  wire __3871__;
  wire __3872__;
  wire __3873__;
  wire __3874__;
  wire __3875__;
  wire __3876__;
  wire __3877__;
  wire __3878__;
  wire __3879__;
  wire __3880__;
  wire __3881__;
  wire __3882__;
  wire __3883__;
  wire __3884__;
  wire __3885__;
  wire __3886__;
  wire __3887__;
  wire __3888__;
  wire __3889__;
  wire __3890__;
  wire __3891__;
  wire __3892__;
  wire __3893__;
  wire __3894__;
  wire __3895__;
  wire __3896__;
  wire __3897__;
  wire __3898__;
  wire __3899__;
  wire __3900__;
  wire __3901__;
  wire __3902__;
  wire __3903__;
  wire __3904__;
  wire __3905__;
  wire __3906__;
  wire __3907__;
  wire __3908__;
  wire __3909__;
  wire __3910__;
  wire __3911__;
  wire __3912__;
  wire __3913__;
  wire __3914__;
  wire __3915__;
  wire __3916__;
  wire __3917__;
  wire __3918__;
  wire __3919__;
  wire __3920__;
  wire __3921__;
  wire __3922__;
  wire __3923__;
  wire __3924__;
  wire __3925__;
  wire __3926__;
  wire __3927__;
  wire __3928__;
  wire __3929__;
  wire __3930__;
  wire __3931__;
  wire __3932__;
  wire __3933__;
  wire __3934__;
  wire __3935__;
  wire __3936__;
  wire __3937__;
  wire __3938__;
  wire __3939__;
  wire __3940__;
  wire __3941__;
  wire __3942__;
  wire __3943__;
  wire __3944__;
  wire __3945__;
  wire __3946__;
  wire __3947__;
  wire __3948__;
  wire __3949__;
  wire __3950__;
  wire __3951__;
  wire __3952__;
  wire __3953__;
  wire __3954__;
  wire __3955__;
  wire __3956__;
  wire __3957__;
  wire __3958__;
  wire __3959__;
  wire __3960__;
  wire __3961__;
  wire __3962__;
  wire __3963__;
  wire __3964__;
  wire __3965__;
  wire __3966__;
  wire __3967__;
  wire __3968__;
  wire __3969__;
  wire __3970__;
  wire __3971__;
  wire __3972__;
  wire __3973__;
  wire __3974__;
  wire __3975__;
  wire __3976__;
  wire __3977__;
  wire __3978__;
  wire __3979__;
  wire __3980__;
  wire __3981__;
  wire __3982__;
  wire __3983__;
  wire __3984__;
  wire __3985__;
  wire __3986__;
  wire __3987__;
  wire __3988__;
  wire __3989__;
  wire __3990__;
  wire __3991__;
  wire __3992__;
  wire __3993__;
  wire __3994__;
  wire __3995__;
  wire __3996__;
  wire __3997__;
  wire __3998__;
  wire __3999__;
  wire __4000__;
  wire __4001__;
  wire __4002__;
  wire __4003__;
  wire __4004__;
  wire __4005__;
  wire __4006__;
  wire __4007__;
  wire __4008__;
  wire __4009__;
  wire __4010__;
  wire __4011__;
  wire __4012__;
  wire __4013__;
  wire __4014__;
  wire __4015__;
  wire __4016__;
  wire __4017__;
  wire __4018__;
  wire __4019__;
  wire __4020__;
  wire __4021__;
  wire __4022__;
  wire __4023__;
  wire __4024__;
  wire __4025__;
  wire __4026__;
  wire __4027__;
  wire __4028__;
  wire __4029__;
  wire __4030__;
  wire __4031__;
  wire __4032__;
  wire __4033__;
  wire __4034__;
  wire __4035__;
  wire __4036__;
  wire __4037__;
  wire __4038__;
  wire __4039__;
  wire __4040__;
  wire __4041__;
  wire __4042__;
  wire __4043__;
  wire __4044__;
  wire __4045__;
  wire __4046__;
  wire __4047__;
  wire __4048__;
  wire __4049__;
  wire __4050__;
  wire __4051__;
  wire __4052__;
  wire __4053__;
  wire __4054__;
  wire __4055__;
  wire __4056__;
  wire __4057__;
  wire __4058__;
  wire __4059__;
  wire __4060__;
  wire __4061__;
  wire __4062__;
  wire __4063__;
  wire __4064__;
  wire __4065__;
  wire __4066__;
  wire __4067__;
  wire __4068__;
  wire __4069__;
  wire __4070__;
  wire __4071__;
  wire __4072__;
  wire __4073__;
  wire __4074__;
  wire __4075__;
  wire __4076__;
  wire __4077__;
  wire __4078__;
  wire __4079__;
  wire __4080__;
  wire __4081__;
  wire __4082__;
  wire __4083__;
  wire __4084__;
  wire __4085__;
  wire __4086__;
  wire __4087__;
  wire __4088__;
  wire __4089__;
  wire __4090__;
  wire __4091__;
  wire __4092__;
  wire __4093__;
  wire __4094__;
  wire __4095__;
  wire __4096__;
  wire __4097__;
  wire __4098__;
  wire __4099__;
  wire __4100__;
  wire __4101__;
  wire __4102__;
  wire __4103__;
  wire __4104__;
  wire __4105__;
  wire __4106__;
  wire __4107__;
  wire __4108__;
  wire __4109__;
  wire __4110__;
  wire __4111__;
  wire __4112__;
  wire __4113__;
  wire __4114__;
  wire __4115__;
  wire __4116__;
  wire __4117__;
  wire __4118__;
  wire __4119__;
  wire __4120__;
  wire __4121__;
  wire __4122__;
  wire __4123__;
  wire __4124__;
  wire __4125__;
  wire __4126__;
  wire __4127__;
  wire __4128__;
  wire __4129__;
  wire __4130__;
  wire __4131__;
  wire __4132__;
  wire __4133__;
  wire __4134__;
  wire __4135__;
  wire __4136__;
  wire __4137__;
  wire __4138__;
  wire __4139__;
  wire __4140__;
  wire __4141__;
  wire __4142__;
  wire __4143__;
  wire __4144__;
  wire __4145__;
  wire __4146__;
  wire __4147__;
  wire __4148__;
  wire __4149__;
  wire __4150__;
  wire __4151__;
  wire __4152__;
  wire __4153__;
  wire __4154__;
  wire __4155__;
  wire __4156__;
  wire __4157__;
  wire __4158__;
  wire __4159__;
  wire __4160__;
  wire __4161__;
  FDRE #(
    .INIT(1'bx)
  ) __4162__ (
    .D(__3195__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__0__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4163__ (
    .D(__3403__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4164__ (
    .D(__2290__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__2__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4165__ (
    .D(__2161__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__3__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4166__ (
    .D(__3623__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__4__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4167__ (
    .D(__2393__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__5__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4168__ (
    .D(__3755__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__6__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4169__ (
    .D(__2301__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__7__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4170__ (
    .D(__3020__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__8__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4171__ (
    .D(__3445__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__9__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4172__ (
    .D(__1854__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__10__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4173__ (
    .D(__3212__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__11__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4174__ (
    .D(__3649__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__12__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4175__ (
    .D(__3972__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__13__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4176__ (
    .D(__3749__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__14__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4177__ (
    .D(__3917__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__15__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4178__ (
    .D(__2653__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__16__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4179__ (
    .D(__3828__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__17__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4180__ (
    .D(__2438__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__18__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4181__ (
    .D(__2797__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__19__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4182__ (
    .D(__1781__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__20__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4183__ (
    .D(__2629__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__21__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4184__ (
    .D(__3933__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__22__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4185__ (
    .D(__2926__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__23__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4186__ (
    .D(__3388__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__24__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4187__ (
    .D(__2019__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__25__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4188__ (
    .D(__3053__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__26__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4189__ (
    .D(__3779__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__27__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4190__ (
    .D(__3251__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__28__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4191__ (
    .D(__3678__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__29__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4192__ (
    .D(__2789__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__30__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4193__ (
    .D(__2961__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__31__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4194__ (
    .D(__3333__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__32__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4195__ (
    .D(__3732__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__33__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4196__ (
    .D(__2820__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__34__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4197__ (
    .D(__2956__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__35__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4198__ (
    .D(__2921__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__36__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4199__ (
    .D(__2620__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__37__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4200__ (
    .D(__2062__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__38__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4201__ (
    .D(__3497__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__39__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4202__ (
    .D(__1925__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__40__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4203__ (
    .D(__2662__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__41__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4204__ (
    .D(__2348__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__42__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4205__ (
    .D(__1835__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__43__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4206__ (
    .D(__3647__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__44__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4207__ (
    .D(__2090__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__45__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4208__ (
    .D(__3542__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__46__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4209__ (
    .D(__3826__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__47__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4210__ (
    .D(__2354__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__48__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4211__ (
    .D(__3559__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__49__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4212__ (
    .D(__3356__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__50__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4213__ (
    .D(__2726__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__51__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4214__ (
    .D(__2560__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__52__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4215__ (
    .D(__1957__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__53__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4216__ (
    .D(__3200__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__54__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4217__ (
    .D(__1940__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__55__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4218__ (
    .D(__3980__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__56__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4219__ (
    .D(__2248__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__57__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4220__ (
    .D(__3841__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__58__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4221__ (
    .D(__4088__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__59__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4222__ (
    .D(__3947__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__60__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4223__ (
    .D(__2268__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__61__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4224__ (
    .D(__3130__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__62__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4225__ (
    .D(__4132__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__63__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4226__ (
    .D(__3485__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__64__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4227__ (
    .D(__3017__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__65__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4228__ (
    .D(__2588__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__66__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4229__ (
    .D(__2755__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__67__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4230__ (
    .D(__3340__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__68__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4231__ (
    .D(__3913__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__69__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4232__ (
    .D(__2279__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__70__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4233__ (
    .D(__4087__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__71__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4234__ (
    .D(__3704__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__72__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4235__ (
    .D(__3687__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__73__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4236__ (
    .D(__3465__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__74__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4237__ (
    .D(__3379__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__75__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4238__ (
    .D(__2278__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__76__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4239__ (
    .D(__2167__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__77__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4240__ (
    .D(__4124__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__78__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4241__ (
    .D(__2246__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__79__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4242__ (
    .D(__3083__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__80__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4243__ (
    .D(__3328__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__81__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4244__ (
    .D(__3285__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__82__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4245__ (
    .D(__3278__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__83__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4246__ (
    .D(__2449__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__84__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4247__ (
    .D(__3548__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__85__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4248__ (
    .D(__1754__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__86__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4249__ (
    .D(__4054__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__87__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4250__ (
    .D(__4099__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__88__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4251__ (
    .D(__1751__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__89__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4252__ (
    .D(__4114__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__90__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4253__ (
    .D(__2963__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__91__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4254__ (
    .D(__3105__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__92__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4255__ (
    .D(__2192__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__93__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4256__ (
    .D(__3392__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__94__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4257__ (
    .D(__3508__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__95__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4258__ (
    .D(__4021__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__96__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4259__ (
    .D(__3601__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__97__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4260__ (
    .D(__1788__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__98__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4261__ (
    .D(__1973__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__99__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4262__ (
    .D(__3555__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__100__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4263__ (
    .D(__2381__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__101__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4264__ (
    .D(__3394__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__102__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4265__ (
    .D(__4152__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__103__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4266__ (
    .D(__1756__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__104__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4267__ (
    .D(__3574__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__105__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4268__ (
    .D(__2537__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__106__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4269__ (
    .D(__3939__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__107__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4270__ (
    .D(__3132__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__108__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4271__ (
    .D(__2888__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__109__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4272__ (
    .D(__2306__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__110__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4273__ (
    .D(__2384__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__111__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4274__ (
    .D(__1975__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__112__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4275__ (
    .D(__3436__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__113__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4276__ (
    .D(__2158__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__114__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4277__ (
    .D(__3502__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__115__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4278__ (
    .D(__3573__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__116__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4279__ (
    .D(__3744__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__117__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4280__ (
    .D(__2086__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__118__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4281__ (
    .D(__2948__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__119__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4282__ (
    .D(__3946__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__120__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4283__ (
    .D(__2115__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__121__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4284__ (
    .D(__2491__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__122__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4285__ (
    .D(__3725__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__123__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4286__ (
    .D(__3271__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__124__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4287__ (
    .D(__2220__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__125__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4288__ (
    .D(__3534__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__126__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4289__ (
    .D(__2859__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__127__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4290__ (
    .D(__3851__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__128__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4291__ (
    .D(__2110__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__129__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4292__ (
    .D(__1812__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__130__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4293__ (
    .D(__1796__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__131__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4294__ (
    .D(__1926__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__132__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4295__ (
    .D(__3214__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__133__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4296__ (
    .D(__1997__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__134__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4297__ (
    .D(__3170__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__135__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4298__ (
    .D(__2845__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__136__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4299__ (
    .D(__4066__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__137__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4300__ (
    .D(__3644__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__138__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4301__ (
    .D(__3452__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__139__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4302__ (
    .D(__3422__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__140__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4303__ (
    .D(__4029__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__141__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4304__ (
    .D(__2933__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__142__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4305__ (
    .D(__3843__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__143__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4306__ (
    .D(__3126__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__144__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4307__ (
    .D(__2974__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__145__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4308__ (
    .D(__3408__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__146__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4309__ (
    .D(__4059__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__147__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4310__ (
    .D(__3654__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__148__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4311__ (
    .D(__3054__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__149__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4312__ (
    .D(__1733__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__150__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4313__ (
    .D(__1996__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__151__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4314__ (
    .D(__2793__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__152__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4315__ (
    .D(__2863__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__153__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4316__ (
    .D(__2964__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__154__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4317__ (
    .D(__4004__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__155__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4318__ (
    .D(__2266__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__156__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4319__ (
    .D(__3169__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__157__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4320__ (
    .D(__3712__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__158__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4321__ (
    .D(__1795__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__159__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4322__ (
    .D(__3538__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__160__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4323__ (
    .D(__2494__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__161__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4324__ (
    .D(__2803__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__162__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4325__ (
    .D(__3078__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__163__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4326__ (
    .D(__3979__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__164__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4327__ (
    .D(__3364__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__165__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4328__ (
    .D(__2250__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__166__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4329__ (
    .D(__3243__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__167__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4330__ (
    .D(__3575__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__168__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4331__ (
    .D(__4103__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__169__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4332__ (
    .D(__2265__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__170__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4333__ (
    .D(__3808__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__171__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4334__ (
    .D(__3467__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__172__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4335__ (
    .D(__2850__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__173__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4336__ (
    .D(__3585__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__174__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4337__ (
    .D(__3656__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__175__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4338__ (
    .D(__3815__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__176__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4339__ (
    .D(__3997__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__177__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4340__ (
    .D(__3685__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__178__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4341__ (
    .D(__2556__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__179__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4342__ (
    .D(__2874__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__180__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4343__ (
    .D(__4012__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__181__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4344__ (
    .D(__1811__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__182__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4345__ (
    .D(__2612__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__183__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4346__ (
    .D(__4045__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__184__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4347__ (
    .D(__3145__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__185__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4348__ (
    .D(__3213__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__186__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4349__ (
    .D(__4089__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__187__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4350__ (
    .D(__2065__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__188__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4351__ (
    .D(__2935__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__189__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4352__ (
    .D(__3553__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__190__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4353__ (
    .D(__3657__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__191__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4354__ (
    .D(__2994__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__192__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4355__ (
    .D(__2819__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__193__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4356__ (
    .D(__2498__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__194__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4357__ (
    .D(__1734__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__195__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4358__ (
    .D(__1904__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__196__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4359__ (
    .D(__3123__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__197__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4360__ (
    .D(__2120__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__198__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4361__ (
    .D(__3719__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__199__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4362__ (
    .D(__2940__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__200__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4363__ (
    .D(__4007__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__201__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4364__ (
    .D(__1792__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__202__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4365__ (
    .D(__3205__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__203__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4366__ (
    .D(__1864__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__204__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4367__ (
    .D(__2397__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__205__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4368__ (
    .D(__3895__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__206__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4369__ (
    .D(__2918__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__207__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4370__ (
    .D(__3790__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__208__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4371__ (
    .D(__2518__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__209__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4372__ (
    .D(__3859__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__210__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4373__ (
    .D(__1881__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__211__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4374__ (
    .D(__1949__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__212__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4375__ (
    .D(__1814__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__213__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4376__ (
    .D(__2298__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__214__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4377__ (
    .D(__2545__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__215__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4378__ (
    .D(__3560__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__216__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4379__ (
    .D(__3745__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__217__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4380__ (
    .D(__3273__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__218__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4381__ (
    .D(__2608__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__219__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4382__ (
    .D(__3840__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__220__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4383__ (
    .D(__3387__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__221__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4384__ (
    .D(__3839__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__222__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4385__ (
    .D(__2541__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__223__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4386__ (
    .D(__3873__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__224__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4387__ (
    .D(__2055__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__225__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4388__ (
    .D(__3516__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__226__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4389__ (
    .D(__3910__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__227__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4390__ (
    .D(__3478__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__228__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4391__ (
    .D(__2795__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__229__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4392__ (
    .D(__2338__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__230__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4393__ (
    .D(__2224__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__231__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4394__ (
    .D(__2232__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__232__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4395__ (
    .D(__2909__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__233__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4396__ (
    .D(__2533__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__234__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4397__ (
    .D(__3218__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__235__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4398__ (
    .D(__4108__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__236__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4399__ (
    .D(__1916__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__237__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4400__ (
    .D(__2827__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__238__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4401__ (
    .D(__3197__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__239__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4402__ (
    .D(__2913__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__240__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4403__ (
    .D(__3876__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__241__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4404__ (
    .D(__3891__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__242__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4405__ (
    .D(__3651__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__243__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4406__ (
    .D(__4028__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__244__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4407__ (
    .D(__2580__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__245__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4408__ (
    .D(__2891__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__246__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4409__ (
    .D(__4001__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__247__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4410__ (
    .D(__2005__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__248__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4411__ (
    .D(__3450__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__249__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4412__ (
    .D(__1743__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__250__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4413__ (
    .D(__2322__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__251__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4414__ (
    .D(__1890__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__252__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4415__ (
    .D(__3302__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__253__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4416__ (
    .D(__2683__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__254__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4417__ (
    .D(__2034__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__255__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4418__ (
    .D(__2057__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__256__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4419__ (
    .D(__3076__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__257__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4420__ (
    .D(__3541__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__258__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4421__ (
    .D(__2693__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__259__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4422__ (
    .D(__3688__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__260__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4423__ (
    .D(__3770__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__261__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4424__ (
    .D(__3330__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__262__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4425__ (
    .D(__2075__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__263__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4426__ (
    .D(__3985__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__264__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4427__ (
    .D(__3359__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__265__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4428__ (
    .D(__3262__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__266__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4429__ (
    .D(__2808__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__267__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4430__ (
    .D(__2263__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__268__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4431__ (
    .D(__3354__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__269__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4432__ (
    .D(__2902__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__270__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4433__ (
    .D(__3860__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__271__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4434__ (
    .D(__3537__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__272__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4435__ (
    .D(__3008__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__273__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4436__ (
    .D(__2117__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__274__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4437__ (
    .D(__2884__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__275__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4438__ (
    .D(__2641__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__276__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4439__ (
    .D(__2425__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__277__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4440__ (
    .D(__3874__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__278__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4441__ (
    .D(__3501__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__279__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4442__ (
    .D(__3655__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__280__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4443__ (
    .D(__2339__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__281__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4444__ (
    .D(__4074__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__282__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4445__ (
    .D(__2864__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__283__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4446__ (
    .D(__2743__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__284__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4447__ (
    .D(__2331__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__285__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4448__ (
    .D(__2297__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__286__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4449__ (
    .D(__3270__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__287__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4450__ (
    .D(__2261__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__288__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4451__ (
    .D(__3035__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__289__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4452__ (
    .D(__4115__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__290__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4453__ (
    .D(__2765__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__291__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4454__ (
    .D(__2513__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__292__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4455__ (
    .D(__2187__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__293__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4456__ (
    .D(__3799__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__294__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4457__ (
    .D(__3703__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__295__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4458__ (
    .D(__3412__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__296__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4459__ (
    .D(__2242__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__297__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4460__ (
    .D(__3432__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__298__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4461__ (
    .D(__4051__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__299__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4462__ (
    .D(__3357__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__300__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4463__ (
    .D(__2231__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__301__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4464__ (
    .D(__3362__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__302__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4465__ (
    .D(__3858__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__303__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4466__ (
    .D(__3982__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__304__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4467__ (
    .D(__3802__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__305__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4468__ (
    .D(__4010__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__306__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4469__ (
    .D(__3100__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__307__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4470__ (
    .D(__2087__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__308__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4471__ (
    .D(__2344__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__309__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4472__ (
    .D(__3492__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__310__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4473__ (
    .D(__3025__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__311__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4474__ (
    .D(__3376__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__312__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4475__ (
    .D(__4086__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__313__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4476__ (
    .D(__4050__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__314__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4477__ (
    .D(__3971__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__315__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4478__ (
    .D(__3973__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__316__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4479__ (
    .D(__3691__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__317__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4480__ (
    .D(__2071__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__318__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4481__ (
    .D(__4049__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__319__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4482__ (
    .D(__3215__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__320__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4483__ (
    .D(__2267__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__321__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4484__ (
    .D(__1831__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__322__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4485__ (
    .D(__2223__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__323__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4486__ (
    .D(__3063__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__324__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4487__ (
    .D(__4067__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__325__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4488__ (
    .D(__2636__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__326__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4489__ (
    .D(__3586__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__327__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4490__ (
    .D(__1966__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__328__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4491__ (
    .D(__2353__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__329__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4492__ (
    .D(__1932__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__330__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4493__ (
    .D(__3684__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__331__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4494__ (
    .D(__1730__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__332__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4495__ (
    .D(__4151__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__333__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4496__ (
    .D(__3294__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__334__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4497__ (
    .D(__1938__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__335__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4498__ (
    .D(__3201__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__336__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4499__ (
    .D(__3098__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__337__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4500__ (
    .D(__2419__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__338__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4501__ (
    .D(__1982__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__339__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4502__ (
    .D(__2098__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__340__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4503__ (
    .D(__4069__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__341__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4504__ (
    .D(__1992__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__342__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4505__ (
    .D(__4048__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__343__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4506__ (
    .D(__3632__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__344__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4507__ (
    .D(__3730__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__345__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4508__ (
    .D(__2626__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__346__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4509__ (
    .D(__2140__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__347__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4510__ (
    .D(__2881__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__348__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4511__ (
    .D(__1840__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__349__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4512__ (
    .D(__1755__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__350__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4513__ (
    .D(__3967__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__351__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4514__ (
    .D(__2546__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__352__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4515__ (
    .D(__1769__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__353__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4516__ (
    .D(__3321__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__354__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4517__ (
    .D(__2054__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__355__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4518__ (
    .D(__2345__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__356__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4519__ (
    .D(__3666__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__357__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4520__ (
    .D(__4060__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__358__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4521__ (
    .D(__4138__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__359__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4522__ (
    .D(__2524__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__360__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4523__ (
    .D(__3571__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__361__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4524__ (
    .D(__2391__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__362__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4525__ (
    .D(__1737__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__363__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4526__ (
    .D(__3423__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__364__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4527__ (
    .D(__2817__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__365__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4528__ (
    .D(__2666__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__366__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4529__ (
    .D(__3561__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__367__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4530__ (
    .D(__3713__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__368__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4531__ (
    .D(__3958__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__369__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4532__ (
    .D(__1971__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__370__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4533__ (
    .D(__3295__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__371__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4534__ (
    .D(__3286__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__372__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4535__ (
    .D(__2327__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__373__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4536__ (
    .D(__2138__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__374__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4537__ (
    .D(__3924__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__375__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4538__ (
    .D(__3493__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__376__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4539__ (
    .D(__3028__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__377__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4540__ (
    .D(__3753__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__378__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4541__ (
    .D(__3238__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__379__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4542__ (
    .D(__3477__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__380__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4543__ (
    .D(__2531__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__381__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4544__ (
    .D(__2953__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__382__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4545__ (
    .D(__2794__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__383__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4546__ (
    .D(__2151__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__384__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4547__ (
    .D(__3429__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__385__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4548__ (
    .D(__3070__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__386__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4549__ (
    .D(__3077__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__387__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4550__ (
    .D(__2333__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__388__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4551__ (
    .D(__3399__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__389__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4552__ (
    .D(__1878__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__390__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4553__ (
    .D(__4003__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__391__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4554__ (
    .D(__3265__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__392__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4555__ (
    .D(__2495__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__393__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4556__ (
    .D(__3852__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__394__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4557__ (
    .D(__2284__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__395__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4558__ (
    .D(__3384__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__396__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4559__ (
    .D(__2766__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__397__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4560__ (
    .D(__2993__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__398__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4561__ (
    .D(__4081__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__399__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4562__ (
    .D(__4057__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__400__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4563__ (
    .D(__2230__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__401__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4564__ (
    .D(__3996__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__402__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4565__ (
    .D(__4121__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__403__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4566__ (
    .D(__1870__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__404__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4567__ (
    .D(__2941__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__405__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4568__ (
    .D(__2768__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__406__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4569__ (
    .D(__4161__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__407__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4570__ (
    .D(__3183__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__408__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4571__ (
    .D(__2867__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__409__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4572__ (
    .D(__2479__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__410__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4573__ (
    .D(__2426__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__411__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4574__ (
    .D(__3618__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__412__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4575__ (
    .D(__2406__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__413__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4576__ (
    .D(__3948__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__414__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4577__ (
    .D(__2462__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__415__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4578__ (
    .D(__2900__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__416__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4579__ (
    .D(__2952__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__417__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4580__ (
    .D(__2930__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__418__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4581__ (
    .D(__2924__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__419__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4582__ (
    .D(__2488__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__420__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4583__ (
    .D(__3904__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__421__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4584__ (
    .D(__2219__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__422__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4585__ (
    .D(__2617__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__423__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4586__ (
    .D(__1914__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__424__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4587__ (
    .D(__3616__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__425__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4588__ (
    .D(__3192__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__426__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4589__ (
    .D(__2717__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__427__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4590__ (
    .D(__2442__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__428__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4591__ (
    .D(__4093__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__429__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4592__ (
    .D(__3661__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__430__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4593__ (
    .D(__3608__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__431__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4594__ (
    .D(__2772__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__432__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4595__ (
    .D(__2987__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__433__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4596__ (
    .D(__2701__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__434__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4597__ (
    .D(__2132__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__435__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4598__ (
    .D(__1990__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__436__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4599__ (
    .D(__3162__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__437__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4600__ (
    .D(__2571__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__438__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4601__ (
    .D(__4149__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__439__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4602__ (
    .D(__3676__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__440__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4603__ (
    .D(__2414__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__441__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4604__ (
    .D(__2461__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__442__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4605__ (
    .D(__3977__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__443__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4606__ (
    .D(__3210__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__444__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4607__ (
    .D(__2907__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__445__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4608__ (
    .D(__4080__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__446__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4609__ (
    .D(__2357__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__447__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4610__ (
    .D(__2824__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__448__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4611__ (
    .D(__3291__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__449__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4612__ (
    .D(__3466__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__450__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4613__ (
    .D(__3099__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__451__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4614__ (
    .D(__3609__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__452__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4615__ (
    .D(__3934__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__453__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4616__ (
    .D(__3011__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__454__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4617__ (
    .D(__2939__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__455__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4618__ (
    .D(__3045__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__456__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4619__ (
    .D(__2547__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__457__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4620__ (
    .D(__4016__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__458__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4621__ (
    .D(__2002__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__459__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4622__ (
    .D(__2866__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__460__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4623__ (
    .D(__1740__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__461__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4624__ (
    .D(__2865__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__462__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4625__ (
    .D(__2194__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__463__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4626__ (
    .D(__3296__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__464__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4627__ (
    .D(__3260__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__465__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4628__ (
    .D(__2959__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__466__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4629__ (
    .D(__2212__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__467__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4630__ (
    .D(__3353__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__468__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4631__ (
    .D(__1746__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__469__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4632__ (
    .D(__1768__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__470__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4633__ (
    .D(__3455__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__471__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4634__ (
    .D(__3697__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__472__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4635__ (
    .D(__2779__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__473__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4636__ (
    .D(__2112__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__474__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4637__ (
    .D(__3919__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__475__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4638__ (
    .D(__2730__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__476__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4639__ (
    .D(__2172__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__477__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4640__ (
    .D(__4073__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__478__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4641__ (
    .D(__3796__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__479__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4642__ (
    .D(__4129__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__480__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4643__ (
    .D(__1838__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__481__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4644__ (
    .D(__3926__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__482__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4645__ (
    .D(__3325__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__483__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4646__ (
    .D(__1806__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__484__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4647__ (
    .D(__2473__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__485__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4648__ (
    .D(__3253__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__486__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4649__ (
    .D(__1823__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__487__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4650__ (
    .D(__2359__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__488__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4651__ (
    .D(__3978__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__489__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4652__ (
    .D(__2227__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__490__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4653__ (
    .D(__1945__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__491__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4654__ (
    .D(__2741__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__492__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4655__ (
    .D(__3500__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__493__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4656__ (
    .D(__3342__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__494__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4657__ (
    .D(__3889__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__495__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4658__ (
    .D(__3848__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__496__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4659__ (
    .D(__2934__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__497__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4660__ (
    .D(__1965__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__498__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4661__ (
    .D(__2162__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__499__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4662__ (
    .D(__3872__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__500__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4663__ (
    .D(__3803__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__501__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4664__ (
    .D(__4062__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__502__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4665__ (
    .D(__3363__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__503__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4666__ (
    .D(__2635__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__504__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4667__ (
    .D(__3293__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__505__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4668__ (
    .D(__2880__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__506__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4669__ (
    .D(__1797__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__507__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4670__ (
    .D(__3591__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__508__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4671__ (
    .D(__2654__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__509__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4672__ (
    .D(__2991__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__510__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4673__ (
    .D(__4076__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__511__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4674__ (
    .D(__3141__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__512__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4675__ (
    .D(__3989__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__513__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4676__ (
    .D(__2781__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__514__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4677__ (
    .D(__1827__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__515__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4678__ (
    .D(__2746__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__516__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4679__ (
    .D(__1839__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__517__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4680__ (
    .D(__1855__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__518__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4681__ (
    .D(__1837__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__519__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4682__ (
    .D(__2367__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__520__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4683__ (
    .D(__4068__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__521__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4684__ (
    .D(__2336__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__522__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4685__ (
    .D(__3963__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__523__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4686__ (
    .D(__1738__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__524__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4687__ (
    .D(__2759__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__525__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4688__ (
    .D(__3761__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__526__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4689__ (
    .D(__2868__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__527__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4690__ (
    .D(__2582__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__528__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4691__ (
    .D(__3758__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__529__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4692__ (
    .D(__3386__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__530__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4693__ (
    .D(__2033__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__531__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4694__ (
    .D(__3992__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__532__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4695__ (
    .D(__3778__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__533__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4696__ (
    .D(__1941__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__534__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4697__ (
    .D(__2295__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__535__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4698__ (
    .D(__3468__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__536__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4699__ (
    .D(__3337__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__537__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4700__ (
    .D(__1822__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__538__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4701__ (
    .D(__3857__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__539__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4702__ (
    .D(__3075__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__540__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4703__ (
    .D(__3303__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__541__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4704__ (
    .D(__2605__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__542__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4705__ (
    .D(__2445__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__543__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4706__ (
    .D(__3300__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__544__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4707__ (
    .D(__2651__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__545__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4708__ (
    .D(__2887__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__546__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4709__ (
    .D(__1829__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__547__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4710__ (
    .D(__3760__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__548__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4711__ (
    .D(__2281__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__549__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4712__ (
    .D(__2482__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__550__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4713__ (
    .D(__2032__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__551__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4714__ (
    .D(__1821__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__552__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4715__ (
    .D(__3185__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__553__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4716__ (
    .D(__4110__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__554__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4717__ (
    .D(__2228__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__555__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4718__ (
    .D(__2247__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__556__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4719__ (
    .D(__3398__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__557__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4720__ (
    .D(__2725__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__558__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4721__ (
    .D(__1922__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__559__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4722__ (
    .D(__3625__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__560__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4723__ (
    .D(__3856__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__561__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4724__ (
    .D(__3729__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__562__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4725__ (
    .D(__2296__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__563__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4726__ (
    .D(__1759__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__564__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4727__ (
    .D(__3523__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__565__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4728__ (
    .D(__2585__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__566__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4729__ (
    .D(__3288__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__567__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4730__ (
    .D(__3938__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__568__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4731__ (
    .D(__1793__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__569__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4732__ (
    .D(__3367__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__570__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4733__ (
    .D(__3121__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__571__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4734__ (
    .D(__2490__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__572__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4735__ (
    .D(__1885__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__573__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4736__ (
    .D(__2767__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__574__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4737__ (
    .D(__3550__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__575__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4738__ (
    .D(__2051__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__576__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4739__ (
    .D(__3572__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__577__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4740__ (
    .D(__3375__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__578__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4741__ (
    .D(__2038__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__579__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4742__ (
    .D(__3805__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__580__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4743__ (
    .D(__2037__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__581__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4744__ (
    .D(__2707__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__582__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4745__ (
    .D(__2758__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__583__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4746__ (
    .D(__2474__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__584__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4747__ (
    .D(__2225__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__585__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4748__ (
    .D(__3401__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__586__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4749__ (
    .D(__2573__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__587__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4750__ (
    .D(__2792__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__588__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4751__ (
    .D(__1842__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__589__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4752__ (
    .D(__3471__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__590__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4753__ (
    .D(__3718__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__591__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4754__ (
    .D(__4011__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__592__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4755__ (
    .D(__3003__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__593__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4756__ (
    .D(__2785__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__594__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4757__ (
    .D(__3414__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__595__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4758__ (
    .D(__1955__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__596__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4759__ (
    .D(__3235__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__597__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4760__ (
    .D(__1813__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__598__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4761__ (
    .D(__2222__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__599__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4762__ (
    .D(__4005__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__600__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4763__ (
    .D(__2704__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__601__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4764__ (
    .D(__1815__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__602__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4765__ (
    .D(__3767__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__603__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4766__ (
    .D(__2405__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__604__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4767__ (
    .D(__3629__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__605__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4768__ (
    .D(__2687__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__606__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4769__ (
    .D(__1798__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__607__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4770__ (
    .D(__2070__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__608__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4771__ (
    .D(__3476__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__609__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4772__ (
    .D(__2857__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__610__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4773__ (
    .D(__2403__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__611__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4774__ (
    .D(__4157__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__612__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4775__ (
    .D(__2179__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__613__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4776__ (
    .D(__3604__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__614__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4777__ (
    .D(__3774__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__615__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4778__ (
    .D(__2137__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__616__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4779__ (
    .D(__2754__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__617__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4780__ (
    .D(__1869__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__618__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4781__ (
    .D(__3096__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__619__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4782__ (
    .D(__2568__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__620__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4783__ (
    .D(__2649__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__621__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4784__ (
    .D(__2241__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__622__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4785__ (
    .D(__2508__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__623__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4786__ (
    .D(__3007__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__624__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4787__ (
    .D(__3930__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__625__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4788__ (
    .D(__3937__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__626__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4789__ (
    .D(__2127__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__627__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4790__ (
    .D(__3846__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__628__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4791__ (
    .D(__2634__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__629__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4792__ (
    .D(__3374__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__630__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4793__ (
    .D(__3777__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__631__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4794__ (
    .D(__3407__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__632__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4795__ (
    .D(__3417__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__633__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4796__ (
    .D(__2363__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__634__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4797__ (
    .D(__3093__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__635__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4798__ (
    .D(__1884__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__636__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4799__ (
    .D(__3526__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__637__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4800__ (
    .D(__1784__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__638__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4801__ (
    .D(__2737__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__639__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4802__ (
    .D(__3915__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__640__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4803__ (
    .D(__1745__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__641__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4804__ (
    .D(__3494__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__642__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4805__ (
    .D(__2080__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__643__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4806__ (
    .D(__1804__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__644__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4807__ (
    .D(__1880__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__645__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4808__ (
    .D(__3323__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__646__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4809__ (
    .D(__3371__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__647__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4810__ (
    .D(__2031__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__648__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4811__ (
    .D(__3628__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__649__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4812__ (
    .D(__1731__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__650__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4813__ (
    .D(__3642__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__651__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4814__ (
    .D(__3522__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__652__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4815__ (
    .D(__2018__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__653__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4816__ (
    .D(__3757__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__654__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4817__ (
    .D(__2310__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__655__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4818__ (
    .D(__4036__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__656__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4819__ (
    .D(__4130__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__657__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4820__ (
    .D(__2378__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__658__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4821__ (
    .D(__3366__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__659__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4822__ (
    .D(__2332__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__660__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4823__ (
    .D(__3172__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__661__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4824__ (
    .D(__3570__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__662__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4825__ (
    .D(__2463__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__663__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4826__ (
    .D(__3329__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__664__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4827__ (
    .D(__2206__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__665__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4828__ (
    .D(__2910__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__666__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4829__ (
    .D(__4071__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__667__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4830__ (
    .D(__2584__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__668__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4831__ (
    .D(__3955__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__669__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4832__ (
    .D(__1937__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__670__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4833__ (
    .D(__4106__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__671__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4834__ (
    .D(__2351__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__672__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4835__ (
    .D(__2697__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__673__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4836__ (
    .D(__4075__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__674__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4837__ (
    .D(__2497__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__675__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4838__ (
    .D(__3067__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__676__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4839__ (
    .D(__4102__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__677__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4840__ (
    .D(__2198__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__678__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4841__ (
    .D(__3319__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__679__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4842__ (
    .D(__3842__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__680__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4843__ (
    .D(__2229__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__681__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4844__ (
    .D(__3717__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__682__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4845__ (
    .D(__3365__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__683__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4846__ (
    .D(__1803__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__684__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4847__ (
    .D(__2828__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__685__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4848__ (
    .D(__3515__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__686__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4849__ (
    .D(__2139__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__687__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4850__ (
    .D(__2540__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__688__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4851__ (
    .D(__2152__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__689__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4852__ (
    .D(__2052__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__690__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4853__ (
    .D(__4070__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__691__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4854__ (
    .D(__3108__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__692__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4855__ (
    .D(__2661__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__693__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4856__ (
    .D(__3807__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__694__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4857__ (
    .D(__3279__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__695__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4858__ (
    .D(__1830__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__696__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4859__ (
    .D(__2042__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__697__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4860__ (
    .D(__1826__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__698__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4861__ (
    .D(__3284__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__699__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4862__ (
    .D(__3639__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__700__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4863__ (
    .D(__3166__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__701__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4864__ (
    .D(__2089__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__702__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4865__ (
    .D(__3327__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__703__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4866__ (
    .D(__1799__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__704__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4867__ (
    .D(__3690__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__705__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4868__ (
    .D(__2979__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__706__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4869__ (
    .D(__3009__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__707__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4870__ (
    .D(__3768__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__708__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4871__ (
    .D(__2492__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__709__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4872__ (
    .D(__3942__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__710__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4873__ (
    .D(__4104__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__711__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4874__ (
    .D(__3047__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__712__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4875__ (
    .D(__2702__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__713__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4876__ (
    .D(__3871__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__714__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4877__ (
    .D(__2925__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__715__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4878__ (
    .D(__3619__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__716__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4879__ (
    .D(__2349__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__717__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4880__ (
    .D(__1780__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__718__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4881__ (
    .D(__2030__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__719__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4882__ (
    .D(__2337__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__720__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4883__ (
    .D(__3174__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__721__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4884__ (
    .D(__2294__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__722__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4885__ (
    .D(__3816__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__723__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4886__ (
    .D(__3986__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__724__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4887__ (
    .D(__3954__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__725__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4888__ (
    .D(__3906__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__726__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4889__ (
    .D(__2015__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__727__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4890__ (
    .D(__3668__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__728__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4891__ (
    .D(__2623__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__729__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4892__ (
    .D(__1771__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__730__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4893__ (
    .D(__3498__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__731__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4894__ (
    .D(__2883__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__732__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4895__ (
    .D(__2823__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__733__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4896__ (
    .D(__3539__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__734__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4897__ (
    .D(__3763__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__735__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4898__ (
    .D(__1841__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__736__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4899__ (
    .D(__2740__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__737__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4900__ (
    .D(__3765__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__738__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4901__ (
    .D(__3613__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__739__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4902__ (
    .D(__3084__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__740__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4903__ (
    .D(__2998__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__741__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4904__ (
    .D(__3019__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__742__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4905__ (
    .D(__2101__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__743__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4906__ (
    .D(__2978__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__744__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4907__ (
    .D(__3669__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__745__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4908__ (
    .D(__3171__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__746__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4909__ (
    .D(__3189__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__747__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4910__ (
    .D(__2521__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__748__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4911__ (
    .D(__2133__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__749__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4912__ (
    .D(__2450__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__750__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4913__ (
    .D(__2885__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__751__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4914__ (
    .D(__3026__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__752__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4915__ (
    .D(__2643__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__753__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4916__ (
    .D(__3641__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__754__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4917__ (
    .D(__4009__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__755__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4918__ (
    .D(__3510__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__756__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4919__ (
    .D(__3069__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__757__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4920__ (
    .D(__2039__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__758__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4921__ (
    .D(__2606__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__759__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4922__ (
    .D(__2703__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__760__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4923__ (
    .D(__3287__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__761__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4924__ (
    .D(__2698__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__762__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4925__ (
    .D(__2437__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__763__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4926__ (
    .D(__2561__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__764__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4927__ (
    .D(__1786__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__765__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4928__ (
    .D(__3689__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__766__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4929__ (
    .D(__3334__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__767__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4930__ (
    .D(__2596__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__768__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4931__ (
    .D(__2782__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__769__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4932__ (
    .D(__2398__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__770__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4933__ (
    .D(__3909__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__771__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4934__ (
    .D(__1977__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__772__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4935__ (
    .D(__3727__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__773__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4936__ (
    .D(__1858__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__774__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4937__ (
    .D(__3734__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__775__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4938__ (
    .D(__3079__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__776__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4939__ (
    .D(__2631__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__777__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4940__ (
    .D(__2088__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__778__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4941__ (
    .D(__1995__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__779__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4942__ (
    .D(__3787__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__780__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4943__ (
    .D(__4043__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__781__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4944__ (
    .D(__1794__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__782__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4945__ (
    .D(__3533__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__783__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4946__ (
    .D(__1732__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__784__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4947__ (
    .D(__2457__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__785__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4948__ (
    .D(__4096__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__786__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4949__ (
    .D(__2059__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__787__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4950__ (
    .D(__3918__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__788__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4951__ (
    .D(__2967__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__789__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4952__ (
    .D(__3711__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__790__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4953__ (
    .D(__2957__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__791__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4954__ (
    .D(__2379__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__792__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4955__ (
    .D(__3336__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__793__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4956__ (
    .D(__1879__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__794__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4957__ (
    .D(__3038__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__795__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4958__ (
    .D(__3503__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__796__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4959__ (
    .D(__2694__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__797__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4960__ (
    .D(__3404__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__798__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4961__ (
    .D(__3469__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__799__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4962__ (
    .D(__3043__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__800__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4963__ (
    .D(__3257__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__801__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4964__ (
    .D(__3970__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__802__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4965__ (
    .D(__3945__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__803__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4966__ (
    .D(__4119__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__804__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4967__ (
    .D(__3673__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__805__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4968__ (
    .D(__2411__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__806__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4969__ (
    .D(__3638__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__807__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4970__ (
    .D(__1910__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__808__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4971__ (
    .D(__2319__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__809__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4972__ (
    .D(__4128__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__810__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4973__ (
    .D(__2682__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__811__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4974__ (
    .D(__2502__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__812__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4975__ (
    .D(__3600__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__813__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4976__ (
    .D(__2433__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__814__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4977__ (
    .D(__2945__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__815__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4978__ (
    .D(__1897__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__816__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4979__ (
    .D(__2734__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__817__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4980__ (
    .D(__3881__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__818__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4981__ (
    .D(__3443__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__819__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4982__ (
    .D(__3177__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__820__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4983__ (
    .D(__2536__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__821__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4984__ (
    .D(__2325__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__822__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4985__ (
    .D(__2970__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__823__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4986__ (
    .D(__3435__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__824__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4987__ (
    .D(__2559__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__825__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4988__ (
    .D(__1779__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__826__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4989__ (
    .D(__2997__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__827__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4990__ (
    .D(__2564__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__828__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4991__ (
    .D(__2721__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__829__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4992__ (
    .D(__2366__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__830__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4993__ (
    .D(__3484__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__831__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4994__ (
    .D(__1947__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__832__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4995__ (
    .D(__3764__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__833__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4996__ (
    .D(__2072__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__834__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4997__ (
    .D(__2932__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__835__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4998__ (
    .D(__4144__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__836__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __4999__ (
    .D(__3272__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__837__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5000__ (
    .D(__1899__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__838__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5001__ (
    .D(__2021__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__839__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5002__ (
    .D(__3061__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__840__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5003__ (
    .D(__3380__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__841__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5004__ (
    .D(__2347__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__842__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5005__ (
    .D(__3966__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__843__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5006__ (
    .D(__2064__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__844__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5007__ (
    .D(__2690__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__845__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5008__ (
    .D(__4027__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__846__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5009__ (
    .D(__3470__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__847__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5010__ (
    .D(__3073__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__848__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5011__ (
    .D(__2102__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__849__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5012__ (
    .D(__2544__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__850__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5013__ (
    .D(__3165__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__851__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5014__ (
    .D(__2429__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__852__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5015__ (
    .D(__2043__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__853__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5016__ (
    .D(__1994__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__854__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5017__ (
    .D(__3884__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__855__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5018__ (
    .D(__4044__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__856__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5019__ (
    .D(__3692__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__857__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5020__ (
    .D(__2209__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__858__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5021__ (
    .D(__2489__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__859__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5022__ (
    .D(__3850__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__860__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5023__ (
    .D(__4018__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__861__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5024__ (
    .D(__3031__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__862__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5025__ (
    .D(__3097__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__863__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5026__ (
    .D(__3046__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__864__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5027__ (
    .D(__3530__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__865__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5028__ (
    .D(__3702__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__866__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5029__ (
    .D(__3965__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__867__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5030__ (
    .D(__1886__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__868__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5031__ (
    .D(__3292__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__869__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5032__ (
    .D(__3239__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__870__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5033__ (
    .D(__3819__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__871__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5034__ (
    .D(__3499__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__872__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5035__ (
    .D(__3430__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__873__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5036__ (
    .D(__2599__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__874__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5037__ (
    .D(__3120__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__875__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5038__ (
    .D(__2017__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__876__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5039__ (
    .D(__2404__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__877__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5040__ (
    .D(__3062__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__878__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5041__ (
    .D(__2664__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__879__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5042__ (
    .D(__3223__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__880__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5043__ (
    .D(__2116__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__881__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5044__ (
    .D(__3624__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__882__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5045__ (
    .D(__3217__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__883__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5046__ (
    .D(__2630__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__884__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5047__ (
    .D(__3617__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__885__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5048__ (
    .D(__3818__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__886__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5049__ (
    .D(__2947__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__887__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5050__ (
    .D(__2153__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__888__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5051__ (
    .D(__4063__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__889__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5052__ (
    .D(__2879__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__890__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5053__ (
    .D(__3128__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__891__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5054__ (
    .D(__2205__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__892__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5055__ (
    .D(__3962__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__893__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5056__ (
    .D(__3428__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__894__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5057__ (
    .D(__2302__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__895__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5058__ (
    .D(__3395__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__896__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5059__ (
    .D(__3941__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__897__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5060__ (
    .D(__3227__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__898__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5061__ (
    .D(__2602__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__899__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5062__ (
    .D(__1809__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__900__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5063__ (
    .D(__3242__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__901__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5064__ (
    .D(__2352__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__902__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5065__ (
    .D(__3029__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__903__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5066__ (
    .D(__3875__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__904__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5067__ (
    .D(__3868__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__905__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5068__ (
    .D(__3320__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__906__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5069__ (
    .D(__3897__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__907__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5070__ (
    .D(__1789__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__908__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5071__ (
    .D(__3297__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__909__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5072__ (
    .D(__3479__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__910__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5073__ (
    .D(__2938__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__911__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5074__ (
    .D(__2519__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__912__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5075__ (
    .D(__3142__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__913__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5076__ (
    .D(__2014__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__914__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5077__ (
    .D(__3866__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__915__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5078__ (
    .D(__2142__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__916__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5079__ (
    .D(__3592__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__917__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5080__ (
    .D(__3596__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__918__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5081__ (
    .D(__2652__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__919__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5082__ (
    .D(__3317__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__920__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5083__ (
    .D(__1970__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__921__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5084__ (
    .D(__3987__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__922__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5085__ (
    .D(__2251__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__923__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5086__ (
    .D(__3480__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__924__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5087__ (
    .D(__2522__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__925__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5088__ (
    .D(__4105__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__926__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5089__ (
    .D(__1857__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__927__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5090__ (
    .D(__2802__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__928__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5091__ (
    .D(__2427__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__929__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5092__ (
    .D(__4111__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__930__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5093__ (
    .D(__1894__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__931__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5094__ (
    .D(__2154__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__932__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5095__ (
    .D(__3487__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__933__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5096__ (
    .D(__3361__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__934__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5097__ (
    .D(__3411__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__935__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5098__ (
    .D(__2723__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__936__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5099__ (
    .D(__2718__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__937__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5100__ (
    .D(__4065__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__938__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5101__ (
    .D(__3274__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__939__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5102__ (
    .D(__3427__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__940__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5103__ (
    .D(__3892__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__941__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5104__ (
    .D(__3558__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__942__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5105__ (
    .D(__2202__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__943__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5106__ (
    .D(__1825__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__944__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5107__ (
    .D(__2016__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__945__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5108__ (
    .D(__3186__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__946__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5109__ (
    .D(__2283__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__947__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5110__ (
    .D(__2539__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__948__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5111__ (
    .D(__3052__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__949__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5112__ (
    .D(__2805__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__950__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5113__ (
    .D(__3578__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__951__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5114__ (
    .D(__2852__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__952__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5115__ (
    .D(__3577__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__953__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5116__ (
    .D(__2157__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__954__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5117__ (
    .D(__2529__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__955__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5118__ (
    .D(__4056__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__956__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5119__ (
    .D(__3999__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__957__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5120__ (
    .D(__3959__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__958__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5121__ (
    .D(__3544__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__959__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5122__ (
    .D(__2965__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__960__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5123__ (
    .D(__3528__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__961__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5124__ (
    .D(__2786__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__962__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5125__ (
    .D(__2665__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__963__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5126__ (
    .D(__2826__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__964__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5127__ (
    .D(__3813__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__965__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5128__ (
    .D(__1958__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__966__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5129__ (
    .D(__3686__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__967__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5130__ (
    .D(__2705__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__968__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5131__ (
    .D(__1872__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__969__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5132__ (
    .D(__3631__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__970__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5133__ (
    .D(__3991__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__971__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5134__ (
    .D(__2644__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__972__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5135__ (
    .D(__2886__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__973__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5136__ (
    .D(__2234__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__974__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5137__ (
    .D(__3650__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__975__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5138__ (
    .D(__4037__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__976__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5139__ (
    .D(__1946__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__977__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5140__ (
    .D(__2390__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__978__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5141__ (
    .D(__2788__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__979__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5142__ (
    .D(__3806__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__980__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5143__ (
    .D(__2056__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__981__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5144__ (
    .D(__4109__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__982__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5145__ (
    .D(__3829__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__983__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5146__ (
    .D(__3801__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__984__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5147__ (
    .D(__2211__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__985__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5148__ (
    .D(__2493__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__986__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5149__ (
    .D(__3282__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__987__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5150__ (
    .D(__3232__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__988__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5151__ (
    .D(__2036__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__989__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5152__ (
    .D(__3746__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__990__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5153__ (
    .D(__3136__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__991__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5154__ (
    .D(__4137__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__992__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5155__ (
    .D(__2273__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__993__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5156__ (
    .D(__3795__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__994__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5157__ (
    .D(__2029__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__995__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5158__ (
    .D(__3834__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__996__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5159__ (
    .D(__3701__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__997__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5160__ (
    .D(__2710__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__998__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5161__ (
    .D(__1981__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__999__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5162__ (
    .D(__2373__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1000__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5163__ (
    .D(__3135__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1001__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5164__ (
    .D(__1820__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1002__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5165__ (
    .D(__1776__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1003__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5166__ (
    .D(__2472__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1004__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5167__ (
    .D(__4160__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1005__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5168__ (
    .D(__2671__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1006__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5169__ (
    .D(__3034__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1007__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5170__ (
    .D(__3683__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1008__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5171__ (
    .D(__3420__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1009__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5172__ (
    .D(__3521__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1010__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5173__ (
    .D(__3665__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1011__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5174__ (
    .D(__3737__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1012__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5175__ (
    .D(__2309__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1013__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5176__ (
    .D(__3014__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1014__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5177__ (
    .D(__3953__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1015__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5178__ (
    .D(__3250__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1016__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5179__ (
    .D(__2593__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1017__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5180__ (
    .D(__3348__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1018__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5181__ (
    .D(__3783__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1019__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5182__ (
    .D(__2552__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1020__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5183__ (
    .D(__3383__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1021__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5184__ (
    .D(__1964__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1022__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5185__ (
    .D(__3118__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1023__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5186__ (
    .D(__3648__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1024__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5187__ (
    .D(__2858__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1025__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5188__ (
    .D(__2509__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1026__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5189__ (
    .D(__2822__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1027__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5190__ (
    .D(__2621__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1028__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5191__ (
    .D(__3590__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1029__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5192__ (
    .D(__3545__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1030__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5193__ (
    .D(__2624__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1031__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5194__ (
    .D(__3037__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1032__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5195__ (
    .D(__1967__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1033__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5196__ (
    .D(__3817__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1034__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5197__ (
    .D(__2169__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1035__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5198__ (
    .D(__2722__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1036__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5199__ (
    .D(__2590__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1037__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5200__ (
    .D(__3605__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1038__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5201__ (
    .D(__3762__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1039__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5202__ (
    .D(__4139__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1040__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5203__ (
    .D(__1810__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1041__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5204__ (
    .D(__2063__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1042__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5205__ (
    .D(__3653__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1043__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5206__ (
    .D(__2256__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1044__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5207__ (
    .D(__3739__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1045__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5208__ (
    .D(__2382__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1046__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5209__ (
    .D(__2061__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1047__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5210__ (
    .D(__2619__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1048__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5211__ (
    .D(__2761__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1049__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5212__ (
    .D(__3804__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1050__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5213__ (
    .D(__3355__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1051__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5214__ (
    .D(__2920__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1052__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5215__ (
    .D(__3131__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1053__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5216__ (
    .D(__3049__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1054__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5217__ (
    .D(__3726__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1055__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5218__ (
    .D(__2171__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1056__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5219__ (
    .D(__3646__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1057__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5220__ (
    .D(__3912__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1058__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5221__ (
    .D(__1770__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1059__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5222__ (
    .D(__2081__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1060__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5223__ (
    .D(__3021__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1061__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5224__ (
    .D(__3144__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1062__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5225__ (
    .D(__2148__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1063__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5226__ (
    .D(__3740__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1064__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5227__ (
    .D(__2369__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1065__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5228__ (
    .D(__3206__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1066__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5229__ (
    .D(__3090__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1067__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5230__ (
    .D(__3643__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1068__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5231__ (
    .D(__2249__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1069__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5232__ (
    .D(__3464__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1070__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5233__ (
    .D(__4008__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1071__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5234__ (
    .D(__3950__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1072__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5235__ (
    .D(__3486__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1073__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5236__ (
    .D(__2581__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1074__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5237__ (
    .D(__4101__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1075__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5238__ (
    .D(__3667__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1076__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5239__ (
    .D(__3835__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1077__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5240__ (
    .D(__2443__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1078__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5241__ (
    .D(__2326__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1079__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5242__ (
    .D(__3332__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1080__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5243__ (
    .D(__3002__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1081__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5244__ (
    .D(__3584__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1082__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5245__ (
    .D(__3231__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1083__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5246__ (
    .D(__1758__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1084__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5247__ (
    .D(__3222__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1085__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5248__ (
    .D(__2642__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1086__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5249__ (
    .D(__3771__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1087__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5250__ (
    .D(__3089__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1088__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5251__ (
    .D(__2973__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1089__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5252__ (
    .D(__2554__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1090__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5253__ (
    .D(__2966__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1091__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5254__ (
    .D(__2618__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1092__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5255__ (
    .D(__2233__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1093__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5256__ (
    .D(__3877__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1094__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5257__ (
    .D(__3645__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1095__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5258__ (
    .D(__2530__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1096__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5259__ (
    .D(__1800__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1097__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5260__ (
    .D(__2870__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1098__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5261__ (
    .D(__2660__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1099__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5262__ (
    .D(__2214__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1100__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5263__ (
    .D(__3595__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1101__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5264__ (
    .D(__1808__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1102__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5265__ (
    .D(__3431__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1103__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5266__ (
    .D(__2769__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1104__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5267__ (
    .D(__3865__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1105__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5268__ (
    .D(__2103__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1106__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5269__ (
    .D(__1956__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1107__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5270__ (
    .D(__3378__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1108__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5271__ (
    .D(__3241__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1109__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5272__ (
    .D(__3335__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1110__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5273__ (
    .D(__3447__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1111__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5274__ (
    .D(__3220__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1112__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5275__ (
    .D(__2483__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1113__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5276__ (
    .D(__4077__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1114__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5277__ (
    .D(__2420__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1115__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5278__ (
    .D(__3759__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1116__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5279__ (
    .D(__3385__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1117__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5280__ (
    .D(__3168__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1118__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5281__ (
    .D(__3275__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1119__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5282__ (
    .D(__3298__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1120__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5283__ (
    .D(__4140__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1121__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5284__ (
    .D(__2607__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1122__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5285__ (
    .D(__2745__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1123__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5286__ (
    .D(__2603__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1124__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5287__ (
    .D(__1846__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1125__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5288__ (
    .D(__2000__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1126__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5289__ (
    .D(__3225__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1127__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5290__ (
    .D(__2204__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1128__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5291__ (
    .D(__3981__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1129__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5292__ (
    .D(__3731__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1130__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5293__ (
    .D(__3281__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1131__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5294__ (
    .D(__2255__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1132__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5295__ (
    .D(__2712__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1133__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5296__ (
    .D(__3072__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1134__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5297__ (
    .D(__2114__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1135__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5298__ (
    .D(__1871__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1136__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5299__ (
    .D(__2134__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1137__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5300__ (
    .D(__3396__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1138__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5301__ (
    .D(__2684__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1139__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5302__ (
    .D(__3532__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1140__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5303__ (
    .D(__3351__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1141__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5304__ (
    .D(__2097__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1142__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5305__ (
    .D(__2895__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1143__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5306__ (
    .D(__2481__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1144__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5307__ (
    .D(__3837__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1145__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5308__ (
    .D(__2919__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1146__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5309__ (
    .D(__2869__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1147__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5310__ (
    .D(__3581__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1148__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5311__ (
    .D(__3557__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1149__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5312__ (
    .D(__3377__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1150__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5313__ (
    .D(__3490__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1151__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5314__ (
    .D(__3143__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1152__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5315__ (
    .D(__2377__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1153__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5316__ (
    .D(__2960__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1154__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5317__ (
    .D(__2598__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1155__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5318__ (
    .D(__2790__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1156__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5319__ (
    .D(__1852__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1157__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5320__ (
    .D(__3211__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1158__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5321__ (
    .D(__2977__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1159__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5322__ (
    .D(__2833__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1160__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5323__ (
    .D(__2168__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1161__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5324__ (
    .D(__3995__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1162__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5325__ (
    .D(__3974__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1163__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5326__ (
    .D(__4085__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1164__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5327__ (
    .D(__2456__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1165__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5328__ (
    .D(__2053__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1166__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5329__ (
    .D(__2173__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1167__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5330__ (
    .D(__1752__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1168__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5331__ (
    .D(__3156__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1169__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5332__ (
    .D(__3463__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1170__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5333__ (
    .D(__2226__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1171__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5334__ (
    .D(__3048__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1172__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5335__ (
    .D(__3184__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1173__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5336__ (
    .D(__3036__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1174__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5337__ (
    .D(__1993__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1175__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5338__ (
    .D(__1834__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1176__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5339__ (
    .D(__2195__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1177__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5340__ (
    .D(__3583__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1178__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5341__ (
    .D(__2350__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1179__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5342__ (
    .D(__4025__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1180__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5343__ (
    .D(__3696__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1181__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5344__ (
    .D(__2818__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1182__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5345__ (
    .D(__3004__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1183__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5346__ (
    .D(__2839__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1184__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5347__ (
    .D(__3569__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1185__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5348__ (
    .D(__2844__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1186__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5349__ (
    .D(__2674__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1187__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5350__ (
    .D(__1954__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1188__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5351__ (
    .D(__3440__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1189__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5352__ (
    .D(__2389__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1190__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5353__ (
    .D(__1877__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1191__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5354__ (
    .D(__3182__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1192__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5355__ (
    .D(__2124__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1193__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5356__ (
    .D(__2454__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1194__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5357__ (
    .D(__2314__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1195__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5358__ (
    .D(__1851__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1196__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5359__ (
    .D(__2984__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1197__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5360__ (
    .D(__2878__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1198__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5361__ (
    .D(__2147__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1199__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5362__ (
    .D(__1935__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1200__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5363__ (
    .D(__3345__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1201__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5364__ (
    .D(__2468__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1202__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5365__ (
    .D(__2024__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1203__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5366__ (
    .D(__3148__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1204__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5367__ (
    .D(__2816__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1205__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5368__ (
    .D(__2013__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1206__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5369__ (
    .D(__2678__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1207__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5370__ (
    .D(__1931__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1208__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5371__ (
    .D(__1902__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1209__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5372__ (
    .D(__2085__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1210__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5373__ (
    .D(__4024__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1211__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5374__ (
    .D(__3001__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1212__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5375__ (
    .D(__3115__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1213__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5376__ (
    .D(__3316__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1214__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5377__ (
    .D(__2990__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1215__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5378__ (
    .D(__3280__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1216__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5379__ (
    .D(__2821__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1217__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5380__ (
    .D(__2128__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1218__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5381__ (
    .D(__2170__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1219__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5382__ (
    .D(__2583__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1220__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5383__ (
    .D(__3324__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1221__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5384__ (
    .D(__1903__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1222__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5385__ (
    .D(__2428__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1223__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5386__ (
    .D(__3318__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1224__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5387__ (
    .D(__3627__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1225__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5388__ (
    .D(__2675__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1226__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5389__ (
    .D(__2035__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1227__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5390__ (
    .D(__3173__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1228__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5391__ (
    .D(__3733__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1229__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5392__ (
    .D(__3956__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1230__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5393__ (
    .D(__2009__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1231__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5394__ (
    .D(__2092__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1232__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5395__ (
    .D(__4134__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1233__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5396__ (
    .D(__2040__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1234__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5397__ (
    .D(__4125__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1235__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5398__ (
    .D(__3491__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1236__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5399__ (
    .D(__3724__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1237__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5400__ (
    .D(__2368__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1238__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5401__ (
    .D(__2058__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1239__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5402__ (
    .D(__3562__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1240__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5403__ (
    .D(__4061__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1241__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5404__ (
    .D(__3066__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1242__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5405__ (
    .D(__2896__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1243__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5406__ (
    .D(__3698__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1244__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5407__ (
    .D(__2689__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1245__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5408__ (
    .D(__1760__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1246__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5409__ (
    .D(__3138__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1247__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5410__ (
    .D(__4042__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1248__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5411__ (
    .D(__2436__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1249__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5412__ (
    .D(__2663__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1250__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5413__ (
    .D(__2050__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1251__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5414__ (
    .D(__1836__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1252__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5415__ (
    .D(__2200__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1253__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5416__ (
    .D(__2542__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1254__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5417__ (
    .D(__2798__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1255__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5418__ (
    .D(__2475__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1256__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5419__ (
    .D(__3551__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1257__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5420__ (
    .D(__1969__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1258__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5421__ (
    .D(__3626__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1259__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5422__ (
    .D(__2458__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1260__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5423__ (
    .D(__3313__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1261__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5424__ (
    .D(__4047__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1262__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5425__ (
    .D(__2201__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1263__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5426__ (
    .D(__3446__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1264__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5427__ (
    .D(__2213__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1265__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5428__ (
    .D(__1976__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1266__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5429__ (
    .D(__1928__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1267__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5430__ (
    .D(__3814__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1268__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5431__ (
    .D(__4120__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1269__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5432__ (
    .D(__3556__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1270__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5433__ (
    .D(__2627__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1271__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5434__ (
    .D(__3994__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1272__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5435__ (
    .D(__3547__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1273__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5436__ (
    .D(__2958__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1274__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5437__ (
    .D(__4006__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1275__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5438__ (
    .D(__3451__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1276__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5439__ (
    .D(__3885__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1277__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5440__ (
    .D(__3051__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1278__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5441__ (
    .D(__3226__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1279__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5442__ (
    .D(__3549__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1280__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5443__ (
    .D(__3957__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1281__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5444__ (
    .D(__3680__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1282__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5445__ (
    .D(__3766__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1283__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5446__ (
    .D(__1921__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1284__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5447__ (
    .D(__2946__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1285__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5448__ (
    .D(__4064__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1286__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5449__ (
    .D(__3612__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1287__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5450__ (
    .D(__3421__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1288__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5451__ (
    .D(__3531__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1289__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5452__ (
    .D(__2150__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1290__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5453__ (
    .D(__3630__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1291__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5454__ (
    .D(__2834__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1292__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5455__ (
    .D(__2851__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1293__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5456__ (
    .D(__3721__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1294__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5457__ (
    .D(__3326__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1295__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5458__ (
    .D(__2597__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1296__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5459__ (
    .D(__3125__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1297__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5460__ (
    .D(__2955__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1298__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5461__ (
    .D(__2049__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1299__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5462__ (
    .D(__1845__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1300__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5463__ (
    .D(__3931__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1301__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5464__ (
    .D(__3914__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1302__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5465__ (
    .D(__2832__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1303__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5466__ (
    .D(__1856__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1304__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5467__ (
    .D(__2575__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1305__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5468__ (
    .D(__2901__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1306__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5469__ (
    .D(__4154__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1307__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5470__ (
    .D(__4141__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1308__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5471__ (
    .D(__1843__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1309__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5472__ (
    .D(__3747__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1310__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5473__ (
    .D(__2480__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1311__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5474__ (
    .D(__1757__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1312__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5475__ (
    .D(__2156__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1313__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5476__ (
    .D(__3139__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1314__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5477__ (
    .D(__4055__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1315__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5478__ (
    .D(__3723__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1316__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5479__ (
    .D(__3137__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1317__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5480__ (
    .D(__2113__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1318__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5481__ (
    .D(__3258__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1319__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5482__ (
    .D(__2904__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1320__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5483__ (
    .D(__3060__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1321__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5484__ (
    .D(__4015__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1322__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5485__ (
    .D(__2041__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1323__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5486__ (
    .D(__2208__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1324__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5487__ (
    .D(__3786__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1325__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5488__ (
    .D(__3163__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1326__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5489__ (
    .D(__3122__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1327__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5490__ (
    .D(__2335__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1328__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5491__ (
    .D(__1991__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1329__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5492__ (
    .D(__1939__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1330__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5493__ (
    .D(__4072__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1331__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5494__ (
    .D(__3576__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1332__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5495__ (
    .D(__2252__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1333__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5496__ (
    .D(__3756__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1334__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5497__ (
    .D(__1736__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1335__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5498__ (
    .D(__3505__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1336__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5499__ (
    .D(__2280__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1337__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5500__ (
    .D(__3074__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1338__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5501__ (
    .D(__1972__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1339__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5502__ (
    .D(__2264__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1340__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5503__ (
    .D(__3869__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1341__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5504__ (
    .D(__3579__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1342__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5505__ (
    .D(__3925__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1343__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5506__ (
    .D(__3923__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1344__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5507__ (
    .D(__3527__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1345__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5508__ (
    .D(__3228__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1346__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5509__ (
    .D(__3855__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1347__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5510__ (
    .D(__3198__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1348__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5511__ (
    .D(__3107__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1349__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5512__ (
    .D(__3864__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1350__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5513__ (
    .D(__2465__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1351__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5514__ (
    .D(__2221__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1352__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5515__ (
    .D(__4014__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1353__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5516__ (
    .D(__1787__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1354__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5517__ (
    .D(__3064__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1355__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5518__ (
    .D(__3722__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1356__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5519__ (
    .D(__2282__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1357__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5520__ (
    .D(__2182__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1358__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5521__ (
    .D(__4035__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1359__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5522__ (
    .D(__3811__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1360__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5523__ (
    .D(__3349__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1361__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5524__ (
    .D(__2174__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1362__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5525__ (
    .D(__3127__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1363__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5526__ (
    .D(__3338__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1364__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5527__ (
    .D(__1785__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1365__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5528__ (
    .D(__3196__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1366__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5529__ (
    .D(__2383__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1367__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5530__ (
    .D(__2873__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1368__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5531__ (
    .D(__2149__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1369__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5532__ (
    .D(__2236__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1370__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5533__ (
    .D(__1766__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1371__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5534__ (
    .D(__2555__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1372__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5535__ (
    .D(__1802__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1373__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5536__ (
    .D(__4100__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1374__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5537__ (
    .D(__3827__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1375__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5538__ (
    .D(__3307__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1376__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5539__ (
    .D(__3695__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1377__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5540__ (
    .D(__2778__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1378__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5541__ (
    .D(__2659__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1379__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5542__ (
    .D(__3922__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1380__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5543__ (
    .D(__2812__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1381__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5544__ (
    .D(__2096__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1382__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5545__ (
    .D(__3426__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1383__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5546__ (
    .D(__3246__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1384__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5547__ (
    .D(__1987__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1385__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5548__ (
    .D(__4040__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1386__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5549__ (
    .D(__3159__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1387__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5550__ (
    .D(__3709__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1388__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5551__ (
    .D(__4084__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1389__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5552__ (
    .D(__2048__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1390__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5553__ (
    .D(__3565__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1391__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5554__ (
    .D(__4034__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1392__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5555__ (
    .D(__2784__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1393__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5556__ (
    .D(__2528__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1394__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5557__ (
    .D(__3154__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1395__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5558__ (
    .D(__3825__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1396__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5559__ (
    .D(__3264__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1397__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5560__ (
    .D(__3112__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1398__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5561__ (
    .D(__4143__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1399__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5562__ (
    .D(__3785__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1400__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5563__ (
    .D(__2937__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1401__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5564__ (
    .D(__2343__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1402__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5565__ (
    .D(__2831__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1403__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5566__ (
    .D(__3961__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1404__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5567__ (
    .D(__2749__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1405__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5568__ (
    .D(__3743__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1406__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5569__ (
    .D(__3087__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1407__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5570__ (
    .D(__4013__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1408__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5571__ (
    .D(__3714__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1409__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5572__ (
    .D(__3993__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1410__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5573__ (
    .D(__2813__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1411__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5574__ (
    .D(__2082__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1412__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5575__ (
    .D(__3728__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1413__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5576__ (
    .D(__4090__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1414__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5577__ (
    .D(__3489__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1415__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5578__ (
    .D(__3350__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1416__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5579__ (
    .D(__2543__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1417__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5580__ (
    .D(__2840__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1418__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5581__ (
    .D(__3620__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1419__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5582__ (
    .D(__2464__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1420__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5583__ (
    .D(__2756__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1421__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5584__ (
    .D(__3454__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1422__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5585__ (
    .D(__3331__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1423__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5586__ (
    .D(__2548__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1424__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5587__ (
    .D(__3820__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1425__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5588__ (
    .D(__3720__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1426__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5589__ (
    .D(__4095__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1427__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5590__ (
    .D(__1828__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1428__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5591__ (
    .D(__1853__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1429__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5592__ (
    .D(__3890__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1430__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5593__ (
    .D(__3151__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1431__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5594__ (
    .D(__1807__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1432__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5595__ (
    .D(__3593__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1433__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5596__ (
    .D(__3899__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1434__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5597__ (
    .D(__2882__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1435__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5598__ (
    .D(__3509__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1436__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5599__ (
    .D(__2155__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1437__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5600__ (
    .D(__3410__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1438__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5601__ (
    .D(__4094__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1439__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5602__ (
    .D(__2574__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1440__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5603__ (
    .D(__2875__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1441__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5604__ (
    .D(__2744__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1442__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5605__ (
    .D(__1735__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1443__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5606__ (
    .D(__3290__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1444__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5607__ (
    .D(__3988__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1445__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5608__ (
    .D(__4041__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1446__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5609__ (
    .D(__4107__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1447__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5610__ (
    .D(__1767__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1448__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5611__ (
    .D(__2572__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1449__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5612__ (
    .D(__1753__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1450__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5613__ (
    .D(__2503__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1451__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5614__ (
    .D(__3457__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1452__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5615__ (
    .D(__2532__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1453__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5616__ (
    .D(__2525__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1454__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5617__ (
    .D(__3514__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1455__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5618__ (
    .D(__2773__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1456__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5619__ (
    .D(__2711__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1457__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5620__ (
    .D(__2334__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1458__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5621__ (
    .D(__2010__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1459__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5622__ (
    .D(__2109__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1460__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5623__ (
    .D(__3998__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1461__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5624__ (
    .D(__2079__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1462__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5625__ (
    .D(__2688__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1463__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5626__ (
    .D(__3911__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1464__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5627__ (
    .D(__3900__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1465__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5628__ (
    .D(__2553__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1466__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5629__ (
    .D(__3552__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1467__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5630__ (
    .D(__3109__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1468__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5631__ (
    .D(__1936__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1469__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5632__ (
    .D(__3027__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1470__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5633__ (
    .D(__2235__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1471__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5634__ (
    .D(__2787__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1472__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5635__ (
    .D(__3582__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1473__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5636__ (
    .D(__3119__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1474__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5637__ (
    .D(__3339__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1475__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5638__ (
    .D(__3752__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1476__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5639__ (
    .D(__2595__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1477__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5640__ (
    .D(__3738__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1478__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5641__ (
    .D(__4150__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1479__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5642__ (
    .D(__2589__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1480__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5643__ (
    .D(__2549__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1481__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5644__ (
    .D(__3059__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1482__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5645__ (
    .D(__3543__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1483__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5646__ (
    .D(__2496__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1484__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5647__ (
    .D(__1891__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1485__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5648__ (
    .D(__2141__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1486__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5649__ (
    .D(__2954__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1487__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5650__ (
    .D(__2254__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1488__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5651__ (
    .D(__3124__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1489__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5652__ (
    .D(__3888__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1490__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5653__ (
    .D(__3024__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1491__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5654__ (
    .D(__3662__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1492__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5655__ (
    .D(__3940__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1493__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5656__ (
    .D(__2077__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1494__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5657__ (
    .D(__2435__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1495__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5658__ (
    .D(__3299__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1496__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5659__ (
    .D(__3990__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1497__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5660__ (
    .D(__3106__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1498__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5661__ (
    .D(__3706__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1499__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5662__ (
    .D(__3233__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1500__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5663__ (
    .D(__3854__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1501__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5664__ (
    .D(__3360__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1502__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5665__ (
    .D(__2686__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1503__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5666__ (
    .D(__3473__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1504__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5667__ (
    .D(__2076__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1505__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5668__ (
    .D(__2739__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1506__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5669__ (
    .D(__2199__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1507__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5670__ (
    .D(__3010__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1508__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5671__ (
    .D(__2020__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1509__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5672__ (
    .D(__2622__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1510__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5673__ (
    .D(__3705__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1511__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5674__ (
    .D(__2706__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1512__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5675__ (
    .D(__3448__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1513__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5676__ (
    .D(__3838__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1514__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5677__ (
    .D(__1764__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1515__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5678__ (
    .D(__2601__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1516__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5679__ (
    .D(__1898__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1517__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5680__ (
    .D(__2181__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1518__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5681__ (
    .D(__1765__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1519__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5682__ (
    .D(__2444__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1520__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5683__ (
    .D(__3927__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1521__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5684__ (
    .D(__2418__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1522__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5685__ (
    .D(__3677__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1523__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5686__ (
    .D(__1968__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1524__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5687__ (
    .D(__2650__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1525__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5688__ (
    .D(__2849__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1526__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5689__ (
    .D(__3472__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1527__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5690__ (
    .D(__3240__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1528__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5691__ (
    .D(__2801__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1529__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5692__ (
    .D(__1948__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1530__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5693__ (
    .D(__1915__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1531__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5694__ (
    .D(__3898__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1532__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5695__ (
    .D(__3908__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1533__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5696__ (
    .D(__3504__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1534__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5697__ (
    .D(__1824__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1535__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5698__ (
    .D(__2100__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1536__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5699__ (
    .D(__3878__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1537__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5700__ (
    .D(__2415__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1538__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5701__ (
    .D(__2800__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1539__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5702__ (
    .D(__2197__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1540__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5703__ (
    .D(__3150__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1541__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5704__ (
    .D(__2060__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1542__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5705__ (
    .D(__1998__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1543__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5706__ (
    .D(__2303__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1544__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5707__ (
    .D(__2538__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1545__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5708__ (
    .D(__2434__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1546__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5709__ (
    .D(__3983__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1547__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5710__ (
    .D(__3058__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1548__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5711__ (
    .D(__2992__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1549__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5712__ (
    .D(__3546__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1550__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5713__ (
    .D(__3580__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1551__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5714__ (
    .D(__3633__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1552__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5715__ (
    .D(__3400__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1553__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5716__ (
    .D(__2825__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1554__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5717__ (
    .D(__3140__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1555__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5718__ (
    .D(__3155__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1556__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5719__ (
    .D(__2912__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1557__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5720__ (
    .D(__3715__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1558__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5721__ (
    .D(__3044__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1559__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5722__ (
    .D(__2872__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1560__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5723__ (
    .D(__3594__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1561__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5724__ (
    .D(__3836__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1562__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5725__ (
    .D(__2696__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1563__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5726__ (
    .D(__3769__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1564__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5727__ (
    .D(__2972__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1565__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5728__ (
    .D(__3462__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1566__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5729__ (
    .D(__3536__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1567__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5730__ (
    .D(__4146__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1568__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5731__ (
    .D(__3461__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1569__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5732__ (
    .D(__2894__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1570__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5733__ (
    .D(__2976__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1571__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5734__ (
    .D(__2108__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1572__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5735__ (
    .D(__2330__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1573__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5736__ (
    .D(__2008__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1574__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5737__ (
    .D(__1763__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1575__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5738__ (
    .D(__2287__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1576__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5739__ (
    .D(__3188__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1577__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5740__ (
    .D(__2729__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1578__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5741__ (
    .D(__1961__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1579__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5742__ (
    .D(__1944__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1580__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5743__ (
    .D(__3312__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1581__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5744__ (
    .D(__3023__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1582__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5745__ (
    .D(__1920__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1583__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5746__ (
    .D(__2376__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1584__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5747__ (
    .D(__2478__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1585__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5748__ (
    .D(__2293__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1586__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5749__ (
    .D(__3513__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1587__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5750__ (
    .D(__3863__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1588__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5751__ (
    .D(__2862__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1589__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5752__ (
    .D(__3057__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1590__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5753__ (
    .D(__3370__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1591__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5754__ (
    .D(__2848__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1592__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5755__ (
    .D(__2611__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1593__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5756__ (
    .D(__2417__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1594__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5757__ (
    .D(__4031__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1595__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5758__ (
    .D(__3589__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1596__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5759__ (
    .D(__3309__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1597__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5760__ (
    .D(__3887__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1598__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5761__ (
    .D(__3230__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1599__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5762__ (
    .D(__2742__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1600__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5763__ (
    .D(__2971__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1601__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5764__ (
    .D(__3853__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1602__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5765__ (
    .D(__1974__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1603__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5766__ (
    .D(__2931__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1604__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5767__ (
    .D(__3216__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1605__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5768__ (
    .D(__3444__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1606__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5769__ (
    .D(__1905__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1607__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5770__ (
    .D(__2908__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1608__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5771__ (
    .D(__2791__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1609__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5772__ (
    .D(__2203__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1610__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5773__ (
    .D(__3164__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1611__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5774__ (
    .D(__2911__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1612__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5775__ (
    .D(__3456__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1613__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5776__ (
    .D(__3219__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1614__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5777__ (
    .D(__4058__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1615__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5778__ (
    .D(__3283__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1616__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5779__ (
    .D(__3247__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1617__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5780__ (
    .D(__3964__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1618__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5781__ (
    .D(__4032__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1619__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5782__ (
    .D(__3341__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1620__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5783__ (
    .D(__2380__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1621__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5784__ (
    .D(__3149__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1622__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5785__ (
    .D(__2594__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1623__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5786__ (
    .D(__2757__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1624__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5787__ (
    .D(__2780__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1625__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5788__ (
    .D(__3352__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1626__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5789__ (
    .D(__3481__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1627__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5790__ (
    .D(__2262__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1628__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5791__ (
    .D(__3751__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1629__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5792__ (
    .D(__4133__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1630__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5793__ (
    .D(__3413__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1631__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5794__ (
    .D(__3050__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1632__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5795__ (
    .D(__2871__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1633__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5796__ (
    .D(__3511__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1634__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5797__ (
    .D(__1859__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1635__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5798__ (
    .D(__4002__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1636__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5799__ (
    .D(__3167__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1637__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5800__ (
    .D(__2455__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1638__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5801__ (
    .D(__3800__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1639__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5802__ (
    .D(__3867__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1640__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5803__ (
    .D(__4026__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1641__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5804__ (
    .D(__1739__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1642__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5805__ (
    .D(__2193__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1643__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5806__ (
    .D(__2514__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1644__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5807__ (
    .D(__2196__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1645__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5808__ (
    .D(__3822__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1646__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5809__ (
    .D(__2210__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1647__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5810__ (
    .D(__2903__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1648__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5811__ (
    .D(__2738__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1649__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5812__ (
    .D(__3397__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1650__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5813__ (
    .D(__1999__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1651__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5814__ (
    .D(__3488__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1652__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5815__ (
    .D(__2091__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1653__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5816__ (
    .D(__1917__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1654__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5817__ (
    .D(__3393__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1655__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5818__ (
    .D(__2600__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1656__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5819__ (
    .D(__2724__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1657__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5820__ (
    .D(__3039__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1658__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5821__ (
    .D(__1833__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1659__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5822__ (
    .D(__3710__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1660__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5823__ (
    .D(__3554__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1661__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5824__ (
    .D(__3611__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1662__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5825__ (
    .D(__1801__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1663__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5826__ (
    .D(__2796__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1664__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5827__ (
    .D(__2667__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1665__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5828__ (
    .D(__2523__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1666__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5829__ (
    .D(__3810__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1667__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5830__ (
    .D(__3849__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1668__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5831__ (
    .D(__2340__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1669__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5832__ (
    .D(__3679__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1670__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5833__ (
    .D(__3750__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1671__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5834__ (
    .D(__3289__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1672__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5835__ (
    .D(__2804__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1673__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5836__ (
    .D(__3830__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1674__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5837__ (
    .D(__3535__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1675__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5838__ (
    .D(__2760__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1676__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5839__ (
    .D(__2892__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1677__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5840__ (
    .D(__2695__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1678__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5841__ (
    .D(__2358__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1679__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5842__ (
    .D(__2207__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1680__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5843__ (
    .D(__2685__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1681__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5844__ (
    .D(__3178__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1682__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5845__ (
    .D(__2565__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1683__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5846__ (
    .D(__2625__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1684__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5847__ (
    .D(__3870__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1685__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5848__ (
    .D(__3640__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1686__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5849__ (
    .D(__1744__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1687__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5850__ (
    .D(__3234__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1688__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5851__ (
    .D(__3071__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1689__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5852__ (
    .D(__2628__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1690__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5853__ (
    .D(__3949__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1691__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5854__ (
    .D(__3259__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1692__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5855__ (
    .D(__2180__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1693__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5856__ (
    .D(__3207__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1694__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5857__ (
    .D(__2253__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1695__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5858__ (
    .D(__3529__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1696__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5859__ (
    .D(__3812__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1697__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5860__ (
    .D(__3621__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1698__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5861__ (
    .D(__2099__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1699__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5862__ (
    .D(__3652__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1700__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5863__ (
    .D(__3030__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1701__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5864__ (
    .D(__2587__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1702__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5865__ (
    .D(__3065__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1703__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5866__ (
    .D(__3821__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1704__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5867__ (
    .D(__3199__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1705__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5868__ (
    .D(__3110__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1706__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5869__ (
    .D(__2799__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1707__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5870__ (
    .D(__3409__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1708__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5871__ (
    .D(__2586__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1709__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5872__ (
    .D(__3453__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1710__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5873__ (
    .D(__3791__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1711__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5874__ (
    .D(__3458__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1712__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5875__ (
    .D(__3780__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1713__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5876__ (
    .D(__1844__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1714__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5877__ (
    .D(__3861__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1715__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5878__ (
    .D(__3517__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1716__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5879__ (
    .D(__2360__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1717__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5880__ (
    .D(__3252__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1718__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5881__ (
    .D(__2001__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1719__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5882__ (
    .D(__3018__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1720__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5883__ (
    .D(__1832__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1721__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5884__ (
    .D(__3896__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1722__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5885__ (
    .D(__3907__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1723__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5886__ (
    .D(__1927__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1724__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5887__ (
    .D(__3088__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1725__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5888__ (
    .D(__1887__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1726__)
  );
  FDRE #(
    .INIT(1'bx)
  ) __5889__ (
    .D(__2078__),
    .C(CK),
    .CE(1'b1),
    .R(1'b0),
    .Q(__1727__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5892__ (
    .I1(RESET),
    .I0(__300__),
    .O(__1730__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5893__ (
    .I1(RESET),
    .I0(__618__),
    .O(__1731__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5894__ (
    .I1(RESET),
    .I0(__785__),
    .O(__1732__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __5895__ (
    .I2(RESET),
    .I1(__146__),
    .I0(__151__),
    .O(__1733__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5896__ (
    .I1(RESET),
    .I0(__228__),
    .O(__1734__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5897__ (
    .I1(RESET),
    .I0(__1411__),
    .O(__1735__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __5898__ (
    .I2(RESET),
    .I1(__1334__),
    .I0(__1288__),
    .O(__1736__)
  );
  LUT4 #(
    .INIT(16'h6900)
  ) __5899__ (
    .I3(RESET),
    .I2(__383__),
    .I1(__362__),
    .I0(__340__),
    .O(__1737__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5900__ (
    .I1(RESET),
    .I0(__492__),
    .O(__1738__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5901__ (
    .I1(RESET),
    .I0(__1610__),
    .O(__1739__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5902__ (
    .I1(RESET),
    .I0(__429__),
    .O(__1740__)
  );
  LUT5 #(
    .INIT(32'h14414114)
  ) __5903__ (
    .I4(__21__),
    .I3(__315__),
    .I2(__15__),
    .I1(__347__),
    .I0(TM0),
    .O(__1741__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __5904__ (
    .I5(TM0),
    .I4(__218__),
    .I3(__250__),
    .I2(__152__),
    .I1(__184__),
    .I0(__283__),
    .O(__1742__)
  );
  LUT6 #(
    .INIT(64'h00fff8f800000000)
  ) __5905__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__1742__),
    .I2(__1741__),
    .I1(TM0),
    .I0(__145__),
    .O(__1743__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5906__ (
    .I1(RESET),
    .I0(__1655__),
    .O(__1744__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5907__ (
    .I1(RESET),
    .I0(__609__),
    .O(__1745__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5908__ (
    .I1(RESET),
    .I0(__437__),
    .O(__1746__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5909__ (
    .I1(TM0),
    .I0(__375__),
    .O(__1747__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __5910__ (
    .I5(TM1),
    .I4(__520__),
    .I3(__424__),
    .I2(__488__),
    .I1(__456__),
    .I0(TM0),
    .O(__1748__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5911__ (
    .I1(TM0),
    .I0(__123__),
    .O(__1749__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __5912__ (
    .I5(TM1),
    .I4(__328__),
    .I3(__36__),
    .I2(__89__),
    .I1(__26__),
    .I0(TM0),
    .O(__1750__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __5913__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__1750__),
    .I2(__1749__),
    .I1(__1748__),
    .I0(__1747__),
    .O(__1751__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5914__ (
    .I1(RESET),
    .I0(__1169__),
    .O(__1752__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5915__ (
    .I1(RESET),
    .I0(__1418__),
    .O(__1753__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5916__ (
    .I1(RESET),
    .I0(__98__),
    .O(__1754__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5917__ (
    .I1(RESET),
    .I0(__318__),
    .O(__1755__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5918__ (
    .I1(RESET),
    .I0(__137__),
    .O(__1756__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __5919__ (
    .I2(RESET),
    .I1(__1343__),
    .I0(__1311__),
    .O(__1757__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5920__ (
    .I1(RESET),
    .I0(__1052__),
    .O(__1758__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __5921__ (
    .I2(RESET),
    .I1(__523__),
    .I0(__563__),
    .O(__1759__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5922__ (
    .I1(RESET),
    .I0(__1214__),
    .O(__1760__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __5923__ (
    .I2(TM0),
    .I1(__1720__),
    .I0(DATA_0_24),
    .O(__1761__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __5924__ (
    .I5(TM1),
    .I4(__1607__),
    .I3(__1639__),
    .I2(__1575__),
    .I1(__1671__),
    .I0(TM0),
    .O(__1762__)
  );
  LUT6 #(
    .INIT(64'hff88f0f000000000)
  ) __5925__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__1762__),
    .I2(__1761__),
    .I1(TM0),
    .I0(__1543__),
    .O(__1763__)
  );
  LUT4 #(
    .INIT(16'h6900)
  ) __5926__ (
    .I3(RESET),
    .I2(__1492__),
    .I1(__1535__),
    .I0(__1514__),
    .O(__1764__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __5927__ (
    .I2(RESET),
    .I1(__1488__),
    .I0(__1518__),
    .O(__1765__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5928__ (
    .I1(RESET),
    .I0(__1372__),
    .O(__1766__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5929__ (
    .I1(RESET),
    .I0(__1416__),
    .O(__1767__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5930__ (
    .I1(RESET),
    .I0(__438__),
    .O(__1768__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __5931__ (
    .I2(RESET),
    .I1(__350__),
    .I0(__352__),
    .O(__1769__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5932__ (
    .I1(RESET),
    .I0(__1027__),
    .O(__1770__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5933__ (
    .I1(RESET),
    .I0(__698__),
    .O(__1771__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5934__ (
    .I1(TM0),
    .I0(__1140__),
    .O(__1772__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __5935__ (
    .I5(TM1),
    .I4(__1259__),
    .I3(__1227__),
    .I2(__1291__),
    .I1(__1195__),
    .I0(TM0),
    .O(__1773__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5936__ (
    .I1(TM0),
    .I0(__971__),
    .O(__1774__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __5937__ (
    .I5(TM1),
    .I4(__1099__),
    .I3(__1035__),
    .I2(__1067__),
    .I1(__1003__),
    .I0(TM0),
    .O(__1775__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __5938__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__1775__),
    .I2(__1774__),
    .I1(__1773__),
    .I0(__1772__),
    .O(__1776__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __5939__ (
    .I5(TM0),
    .I4(__1082__),
    .I3(__1018__),
    .I2(__1050__),
    .I1(__1114__),
    .I0(__933__),
    .O(__1777__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __5940__ (
    .I5(TM0),
    .I4(__890__),
    .I3(__922__),
    .I2(__858__),
    .I1(__826__),
    .I0(__794__),
    .O(__1778__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __5941__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__1778__),
    .I0(__1777__),
    .O(__1779__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5942__ (
    .I1(RESET),
    .I0(__686__),
    .O(__1780__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5943__ (
    .I1(RESET),
    .I0(__14__),
    .O(__1781__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __5944__ (
    .I5(TM0),
    .I4(__894__),
    .I3(__862__),
    .I2(__830__),
    .I1(__926__),
    .I0(__737__),
    .O(__1782__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __5945__ (
    .I5(TM0),
    .I4(__702__),
    .I3(__670__),
    .I2(__638__),
    .I1(__734__),
    .I0(__606__),
    .O(__1783__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __5946__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__1783__),
    .I0(__1782__),
    .O(__1784__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5947__ (
    .I1(RESET),
    .I0(__1366__),
    .O(__1785__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __5948__ (
    .I2(RESET),
    .I1(__764__),
    .I0(__706__),
    .O(__1786__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5949__ (
    .I1(RESET),
    .I0(__1355__),
    .O(__1787__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5950__ (
    .I1(RESET),
    .I0(__81__),
    .O(__1788__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5951__ (
    .I1(RESET),
    .I0(__876__),
    .O(__1789__)
  );
  LUT5 #(
    .INIT(32'h14414114)
  ) __5952__ (
    .I4(__8__),
    .I3(__336__),
    .I2(__304__),
    .I1(__91__),
    .I0(TM0),
    .O(__1790__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __5953__ (
    .I5(TM0),
    .I4(__202__),
    .I3(__169__),
    .I2(__138__),
    .I1(__105__),
    .I0(__299__),
    .O(__1791__)
  );
  LUT6 #(
    .INIT(64'h00fff8f800000000)
  ) __5954__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__1791__),
    .I2(__1790__),
    .I1(TM0),
    .I0(__75__),
    .O(__1792__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __5955__ (
    .I2(RESET),
    .I1(__518__),
    .I0(__568__),
    .O(__1793__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5956__ (
    .I1(RESET),
    .I0(__783__),
    .O(__1794__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __5957__ (
    .I2(RESET),
    .I1(__102__),
    .I0(__154__),
    .O(__1795__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __5958__ (
    .I2(RESET),
    .I1(__196__),
    .I0(__117__),
    .O(__1796__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5959__ (
    .I1(RESET),
    .I0(__475__),
    .O(__1797__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __5960__ (
    .I1(RESET),
    .I0(__576__),
    .O(__1798__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5961__ (
    .I1(RESET),
    .I0(__672__),
    .O(__1799__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5962__ (
    .I1(RESET),
    .I0(__1065__),
    .O(__1800__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5963__ (
    .I1(RESET),
    .I0(__1631__),
    .O(__1801__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5964__ (
    .I1(RESET),
    .I0(__1374__),
    .O(__1802__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5965__ (
    .I1(RESET),
    .I0(__652__),
    .O(__1803__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5966__ (
    .I1(RESET),
    .I0(__612__),
    .O(__1804__)
  );
  LUT6 #(
    .INIT(64'h4bb4b44bb44b4bb4)
  ) __5967__ (
    .I5(__248__),
    .I4(__101__),
    .I3(__182__),
    .I2(__216__),
    .I1(TM0),
    .I0(__281__),
    .O(__1805__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5968__ (
    .I1(RESET),
    .I0(__452__),
    .O(__1806__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5969__ (
    .I1(RESET),
    .I0(__1400__),
    .O(__1807__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5970__ (
    .I1(RESET),
    .I0(__1070__),
    .O(__1808__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5971__ (
    .I1(RESET),
    .I0(__868__),
    .O(__1809__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5972__ (
    .I1(RESET),
    .I0(__1009__),
    .O(__1810__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5973__ (
    .I1(RESET),
    .I0(__216__),
    .O(__1811__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5974__ (
    .I1(RESET),
    .I0(__129__),
    .O(__1812__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5975__ (
    .I1(RESET),
    .I0(__599__),
    .O(__1813__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5976__ (
    .I1(RESET),
    .I0(__263__),
    .O(__1814__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5977__ (
    .I1(RESET),
    .I0(__603__),
    .O(__1815__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5978__ (
    .I1(TM0),
    .I0(__1141__),
    .O(__1816__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __5979__ (
    .I5(TM1),
    .I4(__1194__),
    .I3(__1258__),
    .I2(__1226__),
    .I1(__1290__),
    .I0(TM0),
    .O(__1817__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5980__ (
    .I1(TM0),
    .I0(__970__),
    .O(__1818__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __5981__ (
    .I5(TM1),
    .I4(__1066__),
    .I3(__1034__),
    .I2(__1002__),
    .I1(__1098__),
    .I0(TM0),
    .O(__1819__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __5982__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__1819__),
    .I2(__1818__),
    .I1(__1817__),
    .I0(__1816__),
    .O(__1820__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __5983__ (
    .I2(RESET),
    .I1(__535__),
    .I0(__551__),
    .O(__1821__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5984__ (
    .I1(RESET),
    .I0(__506__),
    .O(__1822__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5985__ (
    .I1(RESET),
    .I0(__455__),
    .O(__1823__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __5986__ (
    .I2(RESET),
    .I1(__1534__),
    .I0(__1472__),
    .O(__1824__)
  );
  LUT4 #(
    .INIT(16'h6900)
  ) __5987__ (
    .I3(RESET),
    .I2(__959__),
    .I1(__911__),
    .I0(__943__),
    .O(__1825__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5988__ (
    .I1(RESET),
    .I0(__666__),
    .O(__1826__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5989__ (
    .I1(RESET),
    .I0(__483__),
    .O(__1827__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5990__ (
    .I1(RESET),
    .I0(__1396__),
    .O(__1828__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __5991__ (
    .I2(RESET),
    .I1(__546__),
    .I0(__540__),
    .O(__1829__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5992__ (
    .I1(RESET),
    .I0(__664__),
    .O(__1830__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5993__ (
    .I1(RESET),
    .I0(__28__),
    .O(__1831__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __5994__ (
    .I2(RESET),
    .I1(__1720__),
    .I0(__1670__),
    .O(__1832__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5995__ (
    .I1(RESET),
    .I0(__1627__),
    .O(__1833__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5996__ (
    .I1(RESET),
    .I0(__1177__),
    .O(__1834__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5997__ (
    .I1(RESET),
    .I0(__42__),
    .O(__1835__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5998__ (
    .I1(RESET),
    .I0(__1220__),
    .O(__1836__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __5999__ (
    .I1(RESET),
    .I0(__487__),
    .O(__1837__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6000__ (
    .I1(RESET),
    .I0(__449__),
    .O(__1838__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6001__ (
    .I1(RESET),
    .I0(__485__),
    .O(__1839__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6002__ (
    .I1(RESET),
    .I0(__317__),
    .O(__1840__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6003__ (
    .I2(RESET),
    .I1(__767__),
    .I0(__735__),
    .O(__1841__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6004__ (
    .I1(RESET),
    .I0(__590__),
    .O(__1842__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6005__ (
    .I1(RESET),
    .I0(__1277__),
    .O(__1843__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6006__ (
    .I2(RESET),
    .I1(__1677__),
    .I0(__1713__),
    .O(__1844__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6007__ (
    .I1(RESET),
    .I0(__1268__),
    .O(__1845__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6008__ (
    .I2(RESET),
    .I1(__1124__),
    .I0(__1114__),
    .O(__1846__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6009__ (
    .I1(TM0),
    .I0(__1331__),
    .O(__1847__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6010__ (
    .I5(TM1),
    .I4(__1452__),
    .I3(__1420__),
    .I2(__1388__),
    .I1(__1484__),
    .I0(TM0),
    .O(__1848__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6011__ (
    .I1(TM0),
    .I0(__1164__),
    .O(__1849__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6012__ (
    .I5(TM1),
    .I4(__1292__),
    .I3(__1196__),
    .I2(__1260__),
    .I1(__1228__),
    .I0(TM0),
    .O(__1850__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __6013__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__1850__),
    .I2(__1849__),
    .I1(__1848__),
    .I0(__1847__),
    .O(__1851__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6014__ (
    .I1(RESET),
    .I0(__1158__),
    .O(__1852__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6015__ (
    .I1(RESET),
    .I0(__1397__),
    .O(__1853__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6016__ (
    .I1(RESET),
    .I0(__77__),
    .O(__1854__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6017__ (
    .I1(RESET),
    .I0(__486__),
    .O(__1855__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6018__ (
    .I1(RESET),
    .I0(__1272__),
    .O(__1856__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6019__ (
    .I1(RESET),
    .I0(__895__),
    .O(__1857__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6020__ (
    .I1(RESET),
    .I0(__775__),
    .O(__1858__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6021__ (
    .I1(RESET),
    .I0(__1603__),
    .O(__1859__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6022__ (
    .I1(TM0),
    .I0(__73__),
    .O(__1860__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6023__ (
    .I5(TM1),
    .I4(__302__),
    .I3(__34__),
    .I2(__87__),
    .I1(__334__),
    .I0(TM0),
    .O(__1861__)
  );
  LUT5 #(
    .INIT(32'h41141441)
  ) __6024__ (
    .I4(__140__),
    .I3(__171__),
    .I2(__204__),
    .I1(__107__),
    .I0(TM0),
    .O(__1862__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6025__ (
    .I1(TM0),
    .I0(__235__),
    .O(__1863__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __6026__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__1863__),
    .I2(__1862__),
    .I1(__1861__),
    .I0(__1860__),
    .O(__1864__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6027__ (
    .I1(TM0),
    .I0(__757__),
    .O(__1865__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6028__ (
    .I5(TM1),
    .I4(__874__),
    .I3(__842__),
    .I2(__810__),
    .I1(__906__),
    .I0(TM0),
    .O(__1866__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6029__ (
    .I1(TM0),
    .I0(__586__),
    .O(__1867__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6030__ (
    .I5(TM1),
    .I4(__682__),
    .I3(__650__),
    .I2(__618__),
    .I1(__714__),
    .I0(TM0),
    .O(__1868__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __6031__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__1868__),
    .I2(__1867__),
    .I1(__1866__),
    .I0(__1865__),
    .O(__1869__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6032__ (
    .I1(RESET),
    .I0(__405__),
    .O(__1870__)
  );
  LUT4 #(
    .INIT(16'h6900)
  ) __6033__ (
    .I3(RESET),
    .I2(__1151__),
    .I1(__1135__),
    .I0(__1103__),
    .O(__1871__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6034__ (
    .I1(RESET),
    .I0(__970__),
    .O(__1872__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6035__ (
    .I1(TM0),
    .I0(__1336__),
    .O(__1873__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6036__ (
    .I5(TM1),
    .I4(__1447__),
    .I3(__1415__),
    .I2(__1383__),
    .I1(__1479__),
    .I0(TM0),
    .O(__1874__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6037__ (
    .I1(TM0),
    .I0(__1159__),
    .O(__1875__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6038__ (
    .I5(TM1),
    .I4(__1255__),
    .I3(__1287__),
    .I2(__1223__),
    .I1(__1191__),
    .I0(TM0),
    .O(__1876__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __6039__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__1876__),
    .I2(__1875__),
    .I1(__1874__),
    .I0(__1873__),
    .O(__1877__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6040__ (
    .I1(RESET),
    .I0(__391__),
    .O(__1878__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6041__ (
    .I1(RESET),
    .I0(__795__),
    .O(__1879__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6042__ (
    .I1(RESET),
    .I0(__613__),
    .O(__1880__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6043__ (
    .I1(RESET),
    .I0(__243__),
    .O(__1881__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6044__ (
    .I5(TM0),
    .I4(__828__),
    .I3(__892__),
    .I2(__860__),
    .I1(__924__),
    .I0(__739__),
    .O(__1882__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6045__ (
    .I5(TM0),
    .I4(__668__),
    .I3(__732__),
    .I2(__700__),
    .I1(__636__),
    .I0(__604__),
    .O(__1883__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __6046__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__1883__),
    .I0(__1882__),
    .O(__1884__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6047__ (
    .I2(RESET),
    .I1(__514__),
    .I0(__572__),
    .O(__1885__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6048__ (
    .I1(RESET),
    .I0(__836__),
    .O(__1886__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6049__ (
    .I2(RESET),
    .I1(__1665__),
    .I0(__1725__),
    .O(__1887__)
  );
  LUT5 #(
    .INIT(32'h14414114)
  ) __6050__ (
    .I4(__309__),
    .I3(__23__),
    .I2(__4__),
    .I1(__341__),
    .I0(TM0),
    .O(__1888__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6051__ (
    .I5(TM0),
    .I4(__100__),
    .I3(__252__),
    .I2(__186__),
    .I1(__220__),
    .I0(__285__),
    .O(__1889__)
  );
  LUT6 #(
    .INIT(64'h00fff8f800000000)
  ) __6052__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__1889__),
    .I2(__1888__),
    .I1(TM0),
    .I0(__143__),
    .O(__1890__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6053__ (
    .I1(RESET),
    .I0(__1453__),
    .O(__1891__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6054__ (
    .I1(TM0),
    .I0(__269__),
    .O(__1892__)
  );
  LUT6 #(
    .INIT(64'h6996966996696996)
  ) __6055__ (
    .I5(TM1),
    .I4(__260__),
    .I3(__292__),
    .I2(__194__),
    .I1(__227__),
    .I0(__1892__),
    .O(__1893__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6056__ (
    .I2(RESET),
    .I1(__930__),
    .I0(__924__),
    .O(__1894__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6057__ (
    .I5(TM0),
    .I4(__1008__),
    .I3(__1040__),
    .I2(__1072__),
    .I1(__1104__),
    .I0(__943__),
    .O(__1895__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6058__ (
    .I5(TM0),
    .I4(__848__),
    .I3(__816__),
    .I2(__880__),
    .I1(__912__),
    .I0(__784__),
    .O(__1896__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __6059__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__1896__),
    .I0(__1895__),
    .O(__1897__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6060__ (
    .I2(RESET),
    .I1(__1516__),
    .I0(__1490__),
    .O(__1898__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6061__ (
    .I1(RESET),
    .I0(__806__),
    .O(__1899__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6062__ (
    .I5(TM0),
    .I4(__1465__),
    .I3(__1433__),
    .I2(__1401__),
    .I1(__1497__),
    .I0(__1318__),
    .O(__1900__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6063__ (
    .I5(TM0),
    .I4(__1209__),
    .I3(__1241__),
    .I2(__1273__),
    .I1(__1305__),
    .I0(__1177__),
    .O(__1901__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __6064__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__1901__),
    .I0(__1900__),
    .O(__1902__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6065__ (
    .I1(RESET),
    .I0(__1190__),
    .O(__1903__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6066__ (
    .I1(RESET),
    .I0(__229__),
    .O(__1904__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6067__ (
    .I1(RESET),
    .I0(__1575__),
    .O(__1905__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6068__ (
    .I1(TM0),
    .I0(__951__),
    .O(__1906__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6069__ (
    .I5(TM1),
    .I4(__1032__),
    .I3(__1000__),
    .I2(__1096__),
    .I1(__1064__),
    .I0(TM0),
    .O(__1907__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6070__ (
    .I1(TM0),
    .I0(__776__),
    .O(__1908__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6071__ (
    .I5(TM1),
    .I4(__872__),
    .I3(__904__),
    .I2(__840__),
    .I1(__808__),
    .I0(TM0),
    .O(__1909__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __6072__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__1909__),
    .I2(__1908__),
    .I1(__1907__),
    .I0(__1906__),
    .O(__1910__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6073__ (
    .I1(TM0),
    .I0(__567__),
    .O(__1911__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6074__ (
    .I5(TM1),
    .I4(__648__),
    .I3(__680__),
    .I2(__712__),
    .I1(__616__),
    .I0(TM0),
    .O(__1912__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6075__ (
    .I1(TM0),
    .I0(__392__),
    .O(__1913__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __6076__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__1913__),
    .I2(__1748__),
    .I1(__1912__),
    .I0(__1911__),
    .O(__1914__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6077__ (
    .I2(RESET),
    .I1(__1476__),
    .I0(__1530__),
    .O(__1915__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6078__ (
    .I1(RESET),
    .I0(__236__),
    .O(__1916__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6079__ (
    .I1(RESET),
    .I0(__1622__),
    .O(__1917__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6080__ (
    .I2(TM0),
    .I1(__1712__),
    .I0(DATA_0_16),
    .O(__1918__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6081__ (
    .I5(TM1),
    .I4(__1583__),
    .I3(__1647__),
    .I2(__1615__),
    .I1(__1679__),
    .I0(TM0),
    .O(__1919__)
  );
  LUT6 #(
    .INIT(64'hff88f0f000000000)
  ) __6082__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__1919__),
    .I2(__1918__),
    .I1(TM0),
    .I0(__1551__),
    .O(__1920__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6083__ (
    .I1(RESET),
    .I0(__1252__),
    .O(__1921__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6084__ (
    .I2(RESET),
    .I1(__558__),
    .I0(__528__),
    .O(__1922__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6085__ (
    .I5(TM0),
    .I4(__476__),
    .I3(__508__),
    .I2(__444__),
    .I1(__540__),
    .I0(__355__),
    .O(__1923__)
  );
  LUT5 #(
    .INIT(32'h14414114)
  ) __6086__ (
    .I4(__316__),
    .I3(__30__),
    .I2(__40__),
    .I1(__348__),
    .I0(TM0),
    .O(__1924__)
  );
  LUT6 #(
    .INIT(64'hff880f0f00000000)
  ) __6087__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__1924__),
    .I2(__1923__),
    .I1(TM0),
    .I0(__98__),
    .O(__1925__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6088__ (
    .I2(RESET),
    .I1(__195__),
    .I0(__118__),
    .O(__1926__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6089__ (
    .I2(RESET),
    .I1(__1723__),
    .I0(__1667__),
    .O(__1927__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6090__ (
    .I1(RESET),
    .I0(__1235__),
    .O(__1928__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6091__ (
    .I5(TM0),
    .I4(__1432__),
    .I3(__1464__),
    .I2(__1400__),
    .I1(__1496__),
    .I0(__1319__),
    .O(__1929__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6092__ (
    .I5(TM0),
    .I4(__1240__),
    .I3(__1208__),
    .I2(__1304__),
    .I1(__1272__),
    .I0(__1176__),
    .O(__1930__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __6093__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__1930__),
    .I0(__1929__),
    .O(__1931__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6094__ (
    .I1(RESET),
    .I0(__25__),
    .O(__1932__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6095__ (
    .I5(TM0),
    .I4(__1456__),
    .I3(__1424__),
    .I2(__1392__),
    .I1(__1488__),
    .I0(__1327__),
    .O(__1933__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6096__ (
    .I5(TM0),
    .I4(__1264__),
    .I3(__1232__),
    .I2(__1200__),
    .I1(__1296__),
    .I0(__1168__),
    .O(__1934__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __6097__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__1934__),
    .I0(__1933__),
    .O(__1935__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6098__ (
    .I1(RESET),
    .I0(__1437__),
    .O(__1936__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6099__ (
    .I1(RESET),
    .I0(__638__),
    .O(__1937__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6100__ (
    .I1(RESET),
    .I0(__303__),
    .O(__1938__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6101__ (
    .I2(RESET),
    .I1(__1293__),
    .I0(__1329__),
    .O(__1939__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6102__ (
    .I1(RESET),
    .I0(__5__),
    .O(__1940__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6103__ (
    .I1(RESET),
    .I0(__502__),
    .O(__1941__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6104__ (
    .I2(TM0),
    .I1(__1715__),
    .I0(DATA_0_19),
    .O(__1942__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6105__ (
    .I5(TM1),
    .I4(__1676__),
    .I3(__1644__),
    .I2(__1612__),
    .I1(__1580__),
    .I0(TM0),
    .O(__1943__)
  );
  LUT6 #(
    .INIT(64'hff88f0f000000000)
  ) __6106__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__1943__),
    .I2(__1942__),
    .I1(TM0),
    .I0(__1548__),
    .O(__1944__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6107__ (
    .I1(RESET),
    .I0(__459__),
    .O(__1945__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6108__ (
    .I1(RESET),
    .I0(__978__),
    .O(__1946__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6109__ (
    .I1(RESET),
    .I0(__800__),
    .O(__1947__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6110__ (
    .I2(RESET),
    .I1(__1477__),
    .I0(__1529__),
    .O(__1948__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6111__ (
    .I1(RESET),
    .I0(__244__),
    .O(__1949__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6112__ (
    .I1(TM0),
    .I0(__1339__),
    .O(__1950__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6113__ (
    .I5(TM1),
    .I4(__1444__),
    .I3(__1412__),
    .I2(__1380__),
    .I1(__1476__),
    .I0(TM0),
    .O(__1951__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6114__ (
    .I1(TM0),
    .I0(__1156__),
    .O(__1952__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6115__ (
    .I5(TM1),
    .I4(__1252__),
    .I3(__1220__),
    .I2(__1188__),
    .I1(__1284__),
    .I0(TM0),
    .O(__1953__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __6116__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__1953__),
    .I2(__1952__),
    .I1(__1951__),
    .I0(__1950__),
    .O(__1954__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6117__ (
    .I1(RESET),
    .I0(__597__),
    .O(__1955__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6118__ (
    .I1(RESET),
    .I0(__1075__),
    .O(__1956__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6119__ (
    .I1(RESET),
    .I0(__63__),
    .O(__1957__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6120__ (
    .I1(RESET),
    .I0(__967__),
    .O(__1958__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6121__ (
    .I2(TM0),
    .I1(__1716__),
    .I0(DATA_0_20),
    .O(__1959__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6122__ (
    .I5(TM1),
    .I4(__1643__),
    .I3(__1675__),
    .I2(__1579__),
    .I1(__1611__),
    .I0(TM0),
    .O(__1960__)
  );
  LUT6 #(
    .INIT(64'hff88f0f000000000)
  ) __6123__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__1960__),
    .I2(__1959__),
    .I1(TM0),
    .I0(__1547__),
    .O(__1961__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6124__ (
    .I5(TM0),
    .I4(__1278__),
    .I3(__1246__),
    .I2(__1214__),
    .I1(__1310__),
    .I0(__1121__),
    .O(__1962__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6125__ (
    .I5(TM0),
    .I4(__1118__),
    .I3(__1086__),
    .I2(__1022__),
    .I1(__1054__),
    .I0(__990__),
    .O(__1963__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __6126__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__1963__),
    .I0(__1962__),
    .O(__1964__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6127__ (
    .I1(RESET),
    .I0(__466__),
    .O(__1965__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6128__ (
    .I1(RESET),
    .I0(__26__),
    .O(__1966__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6129__ (
    .I1(RESET),
    .I0(__1001__),
    .O(__1967__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6130__ (
    .I2(RESET),
    .I1(__1523__),
    .I0(__1483__),
    .O(__1968__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6131__ (
    .I1(RESET),
    .I0(__1226__),
    .O(__1969__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6132__ (
    .I1(RESET),
    .I0(__889__),
    .O(__1970__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6133__ (
    .I2(RESET),
    .I1(__369__),
    .I0(__333__),
    .O(__1971__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6134__ (
    .I2(RESET),
    .I1(__1338__),
    .I0(__1284__),
    .O(__1972__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6135__ (
    .I1(RESET),
    .I0(__82__),
    .O(__1973__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6136__ (
    .I1(RESET),
    .I0(__1571__),
    .O(__1974__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6137__ (
    .I1(RESET),
    .I0(__116__),
    .O(__1975__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6138__ (
    .I1(RESET),
    .I0(__1234__),
    .O(__1976__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6139__ (
    .I1(RESET),
    .I0(__773__),
    .O(__1977__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6140__ (
    .I1(TM0),
    .I0(__1144__),
    .O(__1978__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6141__ (
    .I1(TM0),
    .I0(__967__),
    .O(__1979__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6142__ (
    .I5(TM1),
    .I4(__1063__),
    .I3(__1031__),
    .I2(__999__),
    .I1(__1095__),
    .I0(TM0),
    .O(__1980__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __6143__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__1980__),
    .I2(__1979__),
    .I1(__1876__),
    .I0(__1978__),
    .O(__1981__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6144__ (
    .I1(RESET),
    .I0(__307__),
    .O(__1982__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6145__ (
    .I1(TM0),
    .I0(__1526__),
    .O(__1983__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6146__ (
    .I5(TM1),
    .I4(__1609__),
    .I3(__1673__),
    .I2(__1641__),
    .I1(__1577__),
    .I0(TM0),
    .O(__1984__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6147__ (
    .I1(TM0),
    .I0(__1353__),
    .O(__1985__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6148__ (
    .I5(TM1),
    .I4(__1481__),
    .I3(__1417__),
    .I2(__1449__),
    .I1(__1385__),
    .I0(TM0),
    .O(__1986__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __6149__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__1986__),
    .I2(__1985__),
    .I1(__1984__),
    .I0(__1983__),
    .O(__1987__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6150__ (
    .I5(TM0),
    .I4(__692__),
    .I3(__660__),
    .I2(__628__),
    .I1(__724__),
    .I0(__555__),
    .O(__1988__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6151__ (
    .I5(TM0),
    .I4(__500__),
    .I3(__468__),
    .I2(__436__),
    .I1(__532__),
    .I0(__404__),
    .O(__1989__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __6152__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__1989__),
    .I0(__1988__),
    .O(__1990__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6153__ (
    .I2(RESET),
    .I1(__1328__),
    .I0(__1294__),
    .O(__1991__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6154__ (
    .I1(RESET),
    .I0(__310__),
    .O(__1992__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6155__ (
    .I1(RESET),
    .I0(__1176__),
    .O(__1993__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6156__ (
    .I1(RESET),
    .I0(__822__),
    .O(__1994__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6157__ (
    .I1(RESET),
    .I0(__780__),
    .O(__1995__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6158__ (
    .I1(RESET),
    .I0(__183__),
    .O(__1996__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6159__ (
    .I1(RESET),
    .I0(__141__),
    .O(__1997__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6160__ (
    .I1(RESET),
    .I0(__1544__),
    .O(__1998__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6161__ (
    .I1(RESET),
    .I0(__1619__),
    .O(__1999__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6162__ (
    .I2(RESET),
    .I1(__1125__),
    .I0(__1113__),
    .O(__2000__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6163__ (
    .I2(RESET),
    .I1(__1672__),
    .I0(__1718__),
    .O(__2001__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6164__ (
    .I1(RESET),
    .I0(__427__),
    .O(__2002__)
  );
  LUT5 #(
    .INIT(32'h14414114)
  ) __6165__ (
    .I4(__308__),
    .I3(__55__),
    .I2(__5__),
    .I1(__340__),
    .I0(TM0),
    .O(__2003__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6166__ (
    .I5(TM0),
    .I4(__248__),
    .I3(__101__),
    .I2(__182__),
    .I1(__216__),
    .I0(__281__),
    .O(__2004__)
  );
  LUT6 #(
    .INIT(64'h00fff8f800000000)
  ) __6167__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__2004__),
    .I2(__2003__),
    .I1(TM0),
    .I0(__154__),
    .O(__2005__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6168__ (
    .I2(TM0),
    .I1(__1721__),
    .I0(DATA_0_25),
    .O(__2006__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6169__ (
    .I5(TM1),
    .I4(__1638__),
    .I3(__1574__),
    .I2(__1606__),
    .I1(__1670__),
    .I0(TM0),
    .O(__2007__)
  );
  LUT6 #(
    .INIT(64'hff88f0f000000000)
  ) __6170__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__2007__),
    .I2(__2006__),
    .I1(TM0),
    .I0(__1542__),
    .O(__2008__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6171__ (
    .I1(RESET),
    .I0(__1199__),
    .O(__2009__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6172__ (
    .I1(RESET),
    .I0(__1427__),
    .O(__2010__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6173__ (
    .I5(TM0),
    .I4(__1398__),
    .I3(__1494__),
    .I2(__1462__),
    .I1(__1430__),
    .I0(__1321__),
    .O(__2011__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6174__ (
    .I5(TM0),
    .I4(__1270__),
    .I3(__1238__),
    .I2(__1302__),
    .I1(__1206__),
    .I0(__1174__),
    .O(__2012__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __6175__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__2012__),
    .I0(__2011__),
    .O(__2013__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6176__ (
    .I1(RESET),
    .I0(__882__),
    .O(__2014__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6177__ (
    .I1(RESET),
    .I0(__695__),
    .O(__2015__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6178__ (
    .I2(RESET),
    .I1(__944__),
    .I0(__910__),
    .O(__2016__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6179__ (
    .I1(RESET),
    .I0(__844__),
    .O(__2017__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6180__ (
    .I1(RESET),
    .I0(__621__),
    .O(__2018__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6181__ (
    .I1(RESET),
    .I0(__10__),
    .O(__2019__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6182__ (
    .I2(RESET),
    .I1(__1508__),
    .I0(__1498__),
    .O(__2020__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6183__ (
    .I1(RESET),
    .I0(__807__),
    .O(__2021__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6184__ (
    .I5(TM0),
    .I4(__1395__),
    .I3(__1459__),
    .I2(__1427__),
    .I1(__1491__),
    .I0(__1324__),
    .O(__2022__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6185__ (
    .I5(TM0),
    .I4(__1203__),
    .I3(__1267__),
    .I2(__1235__),
    .I1(__1299__),
    .I0(__1171__),
    .O(__2023__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __6186__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__2023__),
    .I0(__2022__),
    .O(__2024__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6187__ (
    .I1(TM0),
    .I0(__1148__),
    .O(__2025__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6188__ (
    .I5(TM1),
    .I4(__1251__),
    .I3(__1219__),
    .I2(__1187__),
    .I1(__1283__),
    .I0(TM0),
    .O(__2026__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6189__ (
    .I1(TM0),
    .I0(__963__),
    .O(__2027__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6190__ (
    .I5(TM1),
    .I4(__1059__),
    .I3(__1027__),
    .I2(__995__),
    .I1(__1091__),
    .I0(TM0),
    .O(__2028__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __6191__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__2028__),
    .I2(__2027__),
    .I1(__2026__),
    .I0(__2025__),
    .O(__2029__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6192__ (
    .I1(RESET),
    .I0(__687__),
    .O(__2030__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6193__ (
    .I1(RESET),
    .I0(__616__),
    .O(__2031__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6194__ (
    .I2(RESET),
    .I1(__536__),
    .I0(__550__),
    .O(__2032__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6195__ (
    .I1(RESET),
    .I0(__499__),
    .O(__2033__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6196__ (
    .I1(RESET),
    .I0(__259__),
    .O(__2034__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6197__ (
    .I1(RESET),
    .I0(__1195__),
    .O(__2035__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6198__ (
    .I1(RESET),
    .I0(__990__),
    .O(__2036__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6199__ (
    .I1(RESET),
    .I0(__582__),
    .O(__2037__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6200__ (
    .I1(RESET),
    .I0(__580__),
    .O(__2038__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6201__ (
    .I2(RESET),
    .I1(__713__),
    .I0(__757__),
    .O(__2039__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6202__ (
    .I1(RESET),
    .I0(__1202__),
    .O(__2040__)
  );
  LUT4 #(
    .INIT(16'h6900)
  ) __6203__ (
    .I3(RESET),
    .I2(__1322__),
    .I1(__1300__),
    .I0(__1343__),
    .O(__2041__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6204__ (
    .I1(RESET),
    .I0(__665__),
    .O(__2042__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6205__ (
    .I1(RESET),
    .I0(__821__),
    .O(__2043__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6206__ (
    .I1(TM0),
    .I0(__1521__),
    .O(__2044__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6207__ (
    .I5(TM1),
    .I4(__1614__),
    .I3(__1678__),
    .I2(__1582__),
    .I1(__1646__),
    .I0(TM0),
    .O(__2045__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6208__ (
    .I1(TM0),
    .I0(__1358__),
    .O(__2046__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6209__ (
    .I5(TM1),
    .I4(__1486__),
    .I3(__1390__),
    .I2(__1454__),
    .I1(__1422__),
    .I0(TM0),
    .O(__2047__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __6210__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__2047__),
    .I2(__2046__),
    .I1(__2045__),
    .I0(__2044__),
    .O(__2048__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6211__ (
    .I1(RESET),
    .I0(__1267__),
    .O(__2049__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6212__ (
    .I1(RESET),
    .I0(__1219__),
    .O(__2050__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6213__ (
    .I1(RESET),
    .I0(__577__),
    .O(__2051__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6214__ (
    .I1(RESET),
    .I0(__658__),
    .O(__2052__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6215__ (
    .I1(RESET),
    .I0(__1167__),
    .O(__2053__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6216__ (
    .I2(RESET),
    .I1(__348__),
    .I0(__354__),
    .O(__2054__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6217__ (
    .I1(RESET),
    .I0(__201__),
    .O(__2055__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6218__ (
    .I1(RESET),
    .I0(__982__),
    .O(__2056__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6219__ (
    .I1(RESET),
    .I0(__287__),
    .O(__2057__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6220__ (
    .I1(RESET),
    .I0(__1207__),
    .O(__2058__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6221__ (
    .I1(RESET),
    .I0(__788__),
    .O(__2059__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6222__ (
    .I1(RESET),
    .I0(__1543__),
    .O(__2060__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6223__ (
    .I1(RESET),
    .I0(__1015__),
    .O(__2061__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6224__ (
    .I1(RESET),
    .I0(__96__),
    .O(__2062__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6225__ (
    .I1(RESET),
    .I0(__1010__),
    .O(__2063__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6226__ (
    .I1(RESET),
    .I0(__812__),
    .O(__2064__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6227__ (
    .I1(RESET),
    .I0(__192__),
    .O(__2065__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6228__ (
    .I1(TM0),
    .I0(__767__),
    .O(__2066__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6229__ (
    .I5(TM1),
    .I4(__896__),
    .I3(__864__),
    .I2(__832__),
    .I1(__800__),
    .I0(TM0),
    .O(__2067__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6230__ (
    .I1(TM0),
    .I0(__576__),
    .O(__2068__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6231__ (
    .I5(TM1),
    .I4(__608__),
    .I3(__704__),
    .I2(__672__),
    .I1(__640__),
    .I0(TM0),
    .O(__2069__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __6232__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__2069__),
    .I2(__2068__),
    .I1(__2067__),
    .I0(__2066__),
    .O(__2070__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6233__ (
    .I1(RESET),
    .I0(__20__),
    .O(__2071__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6234__ (
    .I1(RESET),
    .I0(__802__),
    .O(__2072__)
  );
  LUT5 #(
    .INIT(32'h14414114)
  ) __6235__ (
    .I4(__52__),
    .I3(__349__),
    .I2(__317__),
    .I1(__62__),
    .I0(TM0),
    .O(__2073__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6236__ (
    .I5(TM0),
    .I4(__179__),
    .I3(__213__),
    .I2(__263__),
    .I1(__147__),
    .I0(__295__),
    .O(__2074__)
  );
  LUT6 #(
    .INIT(64'h00fff8f800000000)
  ) __6237__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__2074__),
    .I2(__2073__),
    .I1(TM0),
    .I0(__157__),
    .O(__2075__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6238__ (
    .I2(RESET),
    .I1(__1502__),
    .I0(__1504__),
    .O(__2076__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6239__ (
    .I1(RESET),
    .I0(__1462__),
    .O(__2077__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6240__ (
    .I2(RESET),
    .I1(__1664__),
    .I0(__1726__),
    .O(__2078__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6241__ (
    .I1(RESET),
    .I0(__1430__),
    .O(__2079__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6242__ (
    .I1(RESET),
    .I0(__611__),
    .O(__2080__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6243__ (
    .I1(RESET),
    .I0(__1028__),
    .O(__2081__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6244__ (
    .I1(RESET),
    .I0(__1380__),
    .O(__2082__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6245__ (
    .I5(TM0),
    .I4(__1402__),
    .I3(__1466__),
    .I2(__1434__),
    .I1(__1498__),
    .I0(__1317__),
    .O(__2083__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6246__ (
    .I5(TM0),
    .I4(__1274__),
    .I3(__1242__),
    .I2(__1210__),
    .I1(__1306__),
    .I0(__1178__),
    .O(__2084__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __6247__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__2084__),
    .I0(__2083__),
    .O(__2085__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6248__ (
    .I2(RESET),
    .I1(__177__),
    .I0(__114__),
    .O(__2086__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6249__ (
    .I1(RESET),
    .I0(__55__),
    .O(__2087__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6250__ (
    .I1(RESET),
    .I0(__779__),
    .O(__2088__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6251__ (
    .I1(RESET),
    .I0(__670__),
    .O(__2089__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6252__ (
    .I1(RESET),
    .I0(__44__),
    .O(__2090__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6253__ (
    .I1(RESET),
    .I0(__1621__),
    .O(__2091__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6254__ (
    .I1(RESET),
    .I0(__1200__),
    .O(__2092__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6255__ (
    .I1(TM0),
    .I0(__1529__),
    .O(__2093__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6256__ (
    .I1(TM0),
    .I0(__1350__),
    .O(__2094__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6257__ (
    .I5(TM1),
    .I4(__1382__),
    .I3(__1414__),
    .I2(__1446__),
    .I1(__1478__),
    .I0(TM0),
    .O(__2095__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __6258__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__2095__),
    .I2(__2094__),
    .I1(__2007__),
    .I0(__2093__),
    .O(__2096__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6259__ (
    .I2(RESET),
    .I1(__1097__),
    .I0(__1141__),
    .O(__2097__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6260__ (
    .I1(RESET),
    .I0(__308__),
    .O(__2098__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6261__ (
    .I2(RESET),
    .I1(__1692__),
    .I0(__1698__),
    .O(__2099__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6262__ (
    .I1(RESET),
    .I0(__1537__),
    .O(__2100__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6263__ (
    .I2(RESET),
    .I1(__728__),
    .I0(__742__),
    .O(__2101__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6264__ (
    .I1(RESET),
    .I0(__817__),
    .O(__2102__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6265__ (
    .I1(RESET),
    .I0(__1074__),
    .O(__2103__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6266__ (
    .I1(TM0),
    .I0(__268__),
    .O(__2104__)
  );
  LUT6 #(
    .INIT(64'h6996966996696996)
  ) __6267__ (
    .I5(TM1),
    .I4(__291__),
    .I3(__242__),
    .I2(__210__),
    .I1(__176__),
    .I0(__2104__),
    .O(__2105__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6268__ (
    .I2(TM0),
    .I1(__1723__),
    .I0(DATA_0_27),
    .O(__2106__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6269__ (
    .I5(TM1),
    .I4(__1604__),
    .I3(__1636__),
    .I2(__1572__),
    .I1(__1668__),
    .I0(TM0),
    .O(__2107__)
  );
  LUT6 #(
    .INIT(64'hff88f0f000000000)
  ) __6270__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__2107__),
    .I2(__2106__),
    .I1(TM0),
    .I0(__1540__),
    .O(__2108__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6271__ (
    .I1(RESET),
    .I0(__1428__),
    .O(__2109__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6272__ (
    .I1(RESET),
    .I0(__111__),
    .O(__2110__)
  );
  LUT6 #(
    .INIT(64'h4bb4b44bb44b4bb4)
  ) __6273__ (
    .I5(__100__),
    .I4(__252__),
    .I3(__186__),
    .I2(__220__),
    .I1(TM0),
    .I0(__285__),
    .O(__2111__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6274__ (
    .I1(RESET),
    .I0(__442__),
    .O(__2112__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6275__ (
    .I2(RESET),
    .I1(__1317__),
    .I0(__1305__),
    .O(__2113__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6276__ (
    .I2(RESET),
    .I1(__1104__),
    .I0(__1134__),
    .O(__2114__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6277__ (
    .I1(RESET),
    .I0(__120__),
    .O(__2115__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6278__ (
    .I1(RESET),
    .I0(__849__),
    .O(__2116__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6279__ (
    .I1(RESET),
    .I0(__273__),
    .O(__2117__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6280__ (
    .I1(TM0),
    .I0(__239__),
    .O(__2118__)
  );
  LUT6 #(
    .INIT(64'h6996966996696996)
  ) __6281__ (
    .I5(TM1),
    .I4(__208__),
    .I3(__175__),
    .I2(__225__),
    .I1(__201__),
    .I0(__2118__),
    .O(__2119__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6282__ (
    .I1(RESET),
    .I0(__230__),
    .O(__2120__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6283__ (
    .I1(TM0),
    .I0(__1334__),
    .O(__2121__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6284__ (
    .I1(TM0),
    .I0(__1161__),
    .O(__2122__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6285__ (
    .I5(TM1),
    .I4(__1289__),
    .I3(__1193__),
    .I2(__1225__),
    .I1(__1257__),
    .I0(TM0),
    .O(__2123__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __6286__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__2123__),
    .I2(__2122__),
    .I1(__1986__),
    .I0(__2121__),
    .O(__2124__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6287__ (
    .I5(TM0),
    .I4(__883__),
    .I3(__851__),
    .I2(__819__),
    .I1(__915__),
    .I0(__748__),
    .O(__2125__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6288__ (
    .I5(TM0),
    .I4(__659__),
    .I3(__691__),
    .I2(__627__),
    .I1(__723__),
    .I0(__595__),
    .O(__2126__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __6289__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__2126__),
    .I0(__2125__),
    .O(__2127__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6290__ (
    .I1(RESET),
    .I0(__1186__),
    .O(__2128__)
  );
  LUT6 #(
    .INIT(64'h4bb4b44bb44b4bb4)
  ) __6291__ (
    .I5(__202__),
    .I4(__169__),
    .I3(__138__),
    .I2(__105__),
    .I1(TM0),
    .I0(__299__),
    .O(__2129__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6292__ (
    .I5(TM0),
    .I4(__659__),
    .I3(__691__),
    .I2(__627__),
    .I1(__723__),
    .I0(__556__),
    .O(__2130__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6293__ (
    .I5(TM0),
    .I4(__499__),
    .I3(__467__),
    .I2(__435__),
    .I1(__531__),
    .I0(__403__),
    .O(__2131__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __6294__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__2131__),
    .I0(__2130__),
    .O(__2132__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6295__ (
    .I2(RESET),
    .I1(__722__),
    .I0(__748__),
    .O(__2133__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6296__ (
    .I2(RESET),
    .I1(__1136__),
    .I0(__1102__),
    .O(__2134__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6297__ (
    .I1(TM0),
    .I0(__759__),
    .O(__2135__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6298__ (
    .I1(TM0),
    .I0(__584__),
    .O(__2136__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __6299__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__2136__),
    .I2(__1912__),
    .I1(__1909__),
    .I0(__2135__),
    .O(__2137__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6300__ (
    .I2(RESET),
    .I1(__329__),
    .I0(__373__),
    .O(__2138__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6301__ (
    .I1(RESET),
    .I0(__655__),
    .O(__2139__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6302__ (
    .I1(RESET),
    .I0(__315__),
    .O(__2140__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6303__ (
    .I1(RESET),
    .I0(__1454__),
    .O(__2141__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6304__ (
    .I1(RESET),
    .I0(__884__),
    .O(__2142__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6305__ (
    .I1(TM0),
    .I0(__1328__),
    .O(__2143__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6306__ (
    .I5(TM1),
    .I4(__1455__),
    .I3(__1423__),
    .I2(__1391__),
    .I1(__1487__),
    .I0(TM0),
    .O(__2144__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6307__ (
    .I1(TM0),
    .I0(__1167__),
    .O(__2145__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6308__ (
    .I5(TM1),
    .I4(__1263__),
    .I3(__1231__),
    .I2(__1199__),
    .I1(__1295__),
    .I0(TM0),
    .O(__2146__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __6309__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__2146__),
    .I2(__2145__),
    .I1(__2144__),
    .I0(__2143__),
    .O(__2147__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6310__ (
    .I1(RESET),
    .I0(__1031__),
    .O(__2148__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6311__ (
    .I1(RESET),
    .I0(__1370__),
    .O(__2149__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6312__ (
    .I1(RESET),
    .I0(__1258__),
    .O(__2150__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6313__ (
    .I1(RESET),
    .I0(__385__),
    .O(__2151__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6314__ (
    .I1(RESET),
    .I0(__657__),
    .O(__2152__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6315__ (
    .I1(RESET),
    .I0(__856__),
    .O(__2153__)
  );
  LUT4 #(
    .INIT(16'h6900)
  ) __6316__ (
    .I3(RESET),
    .I2(__959__),
    .I1(__923__),
    .I0(__931__),
    .O(__2154__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6317__ (
    .I1(RESET),
    .I0(__1405__),
    .O(__2155__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6318__ (
    .I2(RESET),
    .I1(__1312__),
    .I0(__1310__),
    .O(__2156__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6319__ (
    .I2(RESET),
    .I1(__901__),
    .I0(__953__),
    .O(__2157__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6320__ (
    .I2(RESET),
    .I1(__190__),
    .I0(__133__),
    .O(__2158__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6321__ (
    .I5(TM0),
    .I4(__470__),
    .I3(__534__),
    .I2(__502__),
    .I1(__438__),
    .I0(__361__),
    .O(__2159__)
  );
  LUT5 #(
    .INIT(32'h14414114)
  ) __6322__ (
    .I4(__342__),
    .I3(__32__),
    .I2(__3__),
    .I1(__310__),
    .I0(TM0),
    .O(__2160__)
  );
  LUT6 #(
    .INIT(64'hff880f0f00000000)
  ) __6323__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__2160__),
    .I2(__2159__),
    .I1(TM0),
    .I0(__43__),
    .O(__2161__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6324__ (
    .I1(RESET),
    .I0(__467__),
    .O(__2162__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6325__ (
    .I1(TM0),
    .I0(__373__),
    .O(__2163__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6326__ (
    .I5(TM1),
    .I4(__426__),
    .I3(__522__),
    .I2(__490__),
    .I1(__458__),
    .I0(TM0),
    .O(__2164__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6327__ (
    .I1(TM0),
    .I0(__109__),
    .O(__2165__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6328__ (
    .I5(TM1),
    .I4(__25__),
    .I3(__10__),
    .I2(__77__),
    .I1(__330__),
    .I0(TM0),
    .O(__2166__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __6329__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__2166__),
    .I2(__2165__),
    .I1(__2164__),
    .I0(__2163__),
    .O(__2167__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6330__ (
    .I1(RESET),
    .I0(__1162__),
    .O(__2168__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6331__ (
    .I1(RESET),
    .I0(__1003__),
    .O(__2169__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6332__ (
    .I1(RESET),
    .I0(__1187__),
    .O(__2170__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6333__ (
    .I1(RESET),
    .I0(__1024__),
    .O(__2171__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6334__ (
    .I1(RESET),
    .I0(__445__),
    .O(__2172__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6335__ (
    .I1(RESET),
    .I0(__1168__),
    .O(__2173__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6336__ (
    .I1(RESET),
    .I0(__1363__),
    .O(__2174__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6337__ (
    .I1(TM0),
    .I0(__762__),
    .O(__2175__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6338__ (
    .I5(TM1),
    .I4(__869__),
    .I3(__837__),
    .I2(__805__),
    .I1(__901__),
    .I0(TM0),
    .O(__2176__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6339__ (
    .I1(TM0),
    .I0(__581__),
    .O(__2177__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6340__ (
    .I5(TM1),
    .I4(__645__),
    .I3(__677__),
    .I2(__613__),
    .I1(__709__),
    .I0(TM0),
    .O(__2178__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __6341__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__2178__),
    .I2(__2177__),
    .I1(__2176__),
    .I0(__2175__),
    .O(__2179__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6342__ (
    .I1(RESET),
    .I0(__1661__),
    .O(__2180__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6343__ (
    .I2(RESET),
    .I1(__1517__),
    .I0(__1489__),
    .O(__2181__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6344__ (
    .I1(RESET),
    .I0(__1359__),
    .O(__2182__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6345__ (
    .I1(TM0),
    .I0(__132__),
    .O(__2183__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6346__ (
    .I5(TM1),
    .I4(__79__),
    .I3(__323__),
    .I2(__60__),
    .I1(__50__),
    .I0(TM0),
    .O(__2184__)
  );
  LUT5 #(
    .INIT(32'h41141441)
  ) __6347__ (
    .I4(__293__),
    .I3(__228__),
    .I2(__261__),
    .I1(__195__),
    .I0(TM0),
    .O(__2185__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6348__ (
    .I1(TM0),
    .I0(__272__),
    .O(__2186__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __6349__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__2186__),
    .I2(__2185__),
    .I1(__2184__),
    .I0(__2183__),
    .O(__2187__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6350__ (
    .I1(TM0),
    .I0(__371__),
    .O(__2188__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6351__ (
    .I5(TM1),
    .I4(__428__),
    .I3(__460__),
    .I2(__492__),
    .I1(__524__),
    .I0(TM0),
    .O(__2189__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6352__ (
    .I1(TM0),
    .I0(__126__),
    .O(__2190__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6353__ (
    .I5(TM1),
    .I4(__300__),
    .I3(__57__),
    .I2(__93__),
    .I1(__332__),
    .I0(TM0),
    .O(__2191__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __6354__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__2191__),
    .I2(__2190__),
    .I1(__2189__),
    .I0(__2188__),
    .O(__2192__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6355__ (
    .I1(RESET),
    .I0(__1611__),
    .O(__2193__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6356__ (
    .I1(RESET),
    .I0(__431__),
    .O(__2194__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6357__ (
    .I1(RESET),
    .I0(__1178__),
    .O(__2195__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6358__ (
    .I1(RESET),
    .I0(__1613__),
    .O(__2196__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6359__ (
    .I1(RESET),
    .I0(__1541__),
    .O(__2197__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6360__ (
    .I1(RESET),
    .I0(__646__),
    .O(__2198__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6361__ (
    .I2(RESET),
    .I1(__1500__),
    .I0(__1506__),
    .O(__2199__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6362__ (
    .I1(RESET),
    .I0(__1221__),
    .O(__2200__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6363__ (
    .I1(RESET),
    .I0(__1231__),
    .O(__2201__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6364__ (
    .I2(RESET),
    .I1(__942__),
    .I0(__912__),
    .O(__2202__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6365__ (
    .I1(RESET),
    .I0(__1578__),
    .O(__2203__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6366__ (
    .I2(RESET),
    .I1(__1111__),
    .I0(__1127__),
    .O(__2204__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6367__ (
    .I1(RESET),
    .I0(__860__),
    .O(__2205__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6368__ (
    .I1(RESET),
    .I0(__633__),
    .O(__2206__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6369__ (
    .I1(RESET),
    .I0(__1648__),
    .O(__2207__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6370__ (
    .I2(RESET),
    .I1(__1299__),
    .I0(__1323__),
    .O(__2208__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6371__ (
    .I1(RESET),
    .I0(__826__),
    .O(__2209__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6372__ (
    .I1(RESET),
    .I0(__1615__),
    .O(__2210__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6373__ (
    .I1(RESET),
    .I0(__986__),
    .O(__2211__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6374__ (
    .I1(RESET),
    .I0(__435__),
    .O(__2212__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6375__ (
    .I1(RESET),
    .I0(__1233__),
    .O(__2213__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6376__ (
    .I1(RESET),
    .I0(__1068__),
    .O(__2214__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6377__ (
    .I1(TM0),
    .I0(__569__),
    .O(__2215__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6378__ (
    .I5(TM1),
    .I4(__678__),
    .I3(__646__),
    .I2(__614__),
    .I1(__710__),
    .I0(TM0),
    .O(__2216__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6379__ (
    .I1(TM0),
    .I0(__390__),
    .O(__2217__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6380__ (
    .I5(TM1),
    .I4(__486__),
    .I3(__454__),
    .I2(__422__),
    .I1(__518__),
    .I0(TM0),
    .O(__2218__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __6381__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__2218__),
    .I2(__2217__),
    .I1(__2216__),
    .I0(__2215__),
    .O(__2219__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6382__ (
    .I2(RESET),
    .I1(__104__),
    .I0(__158__),
    .O(__2220__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6383__ (
    .I1(RESET),
    .I0(__1353__),
    .O(__2221__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6384__ (
    .I1(RESET),
    .I0(__600__),
    .O(__2222__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6385__ (
    .I1(RESET),
    .I0(__50__),
    .O(__2223__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6386__ (
    .I1(RESET),
    .I0(__265__),
    .O(__2224__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6387__ (
    .I1(RESET),
    .I0(__586__),
    .O(__2225__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6388__ (
    .I1(RESET),
    .I0(__1172__),
    .O(__2226__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6389__ (
    .I1(RESET),
    .I0(__458__),
    .O(__2227__)
  );
  LUT4 #(
    .INIT(16'h6900)
  ) __6390__ (
    .I3(RESET),
    .I2(__554__),
    .I1(__575__),
    .I0(__532__),
    .O(__2228__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6391__ (
    .I1(RESET),
    .I0(__649__),
    .O(__2229__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6392__ (
    .I1(RESET),
    .I0(__402__),
    .O(__2230__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6393__ (
    .I1(RESET),
    .I0(__9__),
    .O(__2231__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6394__ (
    .I1(RESET),
    .I0(__266__),
    .O(__2232__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6395__ (
    .I1(RESET),
    .I0(__1061__),
    .O(__2233__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6396__ (
    .I1(RESET),
    .I0(__975__),
    .O(__2234__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6397__ (
    .I1(RESET),
    .I0(__1439__),
    .O(__2235__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6398__ (
    .I1(RESET),
    .I0(__1371__),
    .O(__2236__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6399__ (
    .I1(TM0),
    .I0(__753__),
    .O(__2237__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6400__ (
    .I5(TM1),
    .I4(__814__),
    .I3(__878__),
    .I2(__846__),
    .I1(__910__),
    .I0(TM0),
    .O(__2238__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6401__ (
    .I1(TM0),
    .I0(__590__),
    .O(__2239__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6402__ (
    .I5(TM1),
    .I4(__622__),
    .I3(__686__),
    .I2(__654__),
    .I1(__718__),
    .I0(TM0),
    .O(__2240__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __6403__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__2240__),
    .I2(__2239__),
    .I1(__2238__),
    .I0(__2237__),
    .O(__2241__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6404__ (
    .I1(RESET),
    .I0(__280__),
    .O(__2242__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6405__ (
    .I1(TM0),
    .I0(__380__),
    .O(__2243__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6406__ (
    .I5(TM1),
    .I4(__451__),
    .I3(__419__),
    .I2(__483__),
    .I1(__515__),
    .I0(TM0),
    .O(__2244__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6407__ (
    .I1(TM0),
    .I0(__129__),
    .O(__2245__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __6408__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__2245__),
    .I2(__2184__),
    .I1(__2244__),
    .I0(__2243__),
    .O(__2246__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6409__ (
    .I2(RESET),
    .I1(__531__),
    .I0(__555__),
    .O(__2247__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6410__ (
    .I1(RESET),
    .I0(__93__),
    .O(__2248__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6411__ (
    .I1(RESET),
    .I0(__1037__),
    .O(__2249__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6412__ (
    .I1(RESET),
    .I0(__200__),
    .O(__2250__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6413__ (
    .I1(RESET),
    .I0(__891__),
    .O(__2251__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6414__ (
    .I2(RESET),
    .I1(__1290__),
    .I0(__1332__),
    .O(__2252__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6415__ (
    .I1(RESET),
    .I0(__1663__),
    .O(__2253__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6416__ (
    .I1(RESET),
    .I0(__1456__),
    .O(__2254__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6417__ (
    .I2(RESET),
    .I1(__1131__),
    .I0(__1107__),
    .O(__2255__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6418__ (
    .I1(RESET),
    .I0(__1012__),
    .O(__2256__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6419__ (
    .I1(TM0),
    .I0(__113__),
    .O(__2257__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6420__ (
    .I5(TM1),
    .I4(__28__),
    .I3(__38__),
    .I2(__96__),
    .I1(__322__),
    .I0(TM0),
    .O(__2258__)
  );
  LUT5 #(
    .INIT(32'h41141441)
  ) __6421__ (
    .I4(__223__),
    .I3(__191__),
    .I2(__288__),
    .I1(__257__),
    .I0(TM0),
    .O(__2259__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6422__ (
    .I1(TM0),
    .I0(__273__),
    .O(__2260__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __6423__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__2260__),
    .I2(__2259__),
    .I1(__2258__),
    .I0(__2257__),
    .O(__2261__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6424__ (
    .I1(RESET),
    .I0(__1596__),
    .O(__2262__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6425__ (
    .I1(RESET),
    .I0(__241__),
    .O(__2263__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6426__ (
    .I2(RESET),
    .I1(__1339__),
    .I0(__1283__),
    .O(__2264__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6427__ (
    .I1(RESET),
    .I0(__203__),
    .O(__2265__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6428__ (
    .I2(RESET),
    .I1(__148__),
    .I0(__145__),
    .O(__2266__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6429__ (
    .I1(RESET),
    .I0(__19__),
    .O(__2267__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6430__ (
    .I1(RESET),
    .I0(__80__),
    .O(__2268__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6431__ (
    .I1(TM0),
    .I0(__1150__),
    .O(__2269__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6432__ (
    .I5(TM1),
    .I4(__1249__),
    .I3(__1281__),
    .I2(__1217__),
    .I1(__1185__),
    .I0(TM0),
    .O(__2270__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6433__ (
    .I1(TM0),
    .I0(__961__),
    .O(__2271__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6434__ (
    .I5(TM1),
    .I4(__1025__),
    .I3(__1089__),
    .I2(__1057__),
    .I1(__993__),
    .I0(TM0),
    .O(__2272__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __6435__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__2272__),
    .I2(__2271__),
    .I1(__2270__),
    .I0(__2269__),
    .O(__2273__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6436__ (
    .I1(TM0),
    .I0(__370__),
    .O(__2274__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6437__ (
    .I5(TM1),
    .I4(__493__),
    .I3(__461__),
    .I2(__429__),
    .I1(__525__),
    .I0(TM0),
    .O(__2275__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6438__ (
    .I1(TM0),
    .I0(__108__),
    .O(__2276__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6439__ (
    .I5(TM1),
    .I4(__301__),
    .I3(__76__),
    .I2(__9__),
    .I1(__333__),
    .I0(TM0),
    .O(__2277__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __6440__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__2277__),
    .I2(__2276__),
    .I1(__2275__),
    .I0(__2274__),
    .O(__2278__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6441__ (
    .I2(RESET),
    .I1(__188__),
    .I0(__71__),
    .O(__2279__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6442__ (
    .I2(RESET),
    .I1(__1336__),
    .I0(__1286__),
    .O(__2280__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6443__ (
    .I2(RESET),
    .I1(__538__),
    .I0(__548__),
    .O(__2281__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6444__ (
    .I1(RESET),
    .I0(__1358__),
    .O(__2282__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6445__ (
    .I2(RESET),
    .I1(__946__),
    .I0(__908__),
    .O(__2283__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6446__ (
    .I1(RESET),
    .I0(__396__),
    .O(__2284__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6447__ (
    .I2(TM0),
    .I1(__1719__),
    .I0(DATA_0_23),
    .O(__2285__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6448__ (
    .I5(TM1),
    .I4(__1608__),
    .I3(__1640__),
    .I2(__1576__),
    .I1(__1672__),
    .I0(TM0),
    .O(__2286__)
  );
  LUT6 #(
    .INIT(64'hff88f0f000000000)
  ) __6449__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__2286__),
    .I2(__2285__),
    .I1(TM0),
    .I0(__1544__),
    .O(__2287__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6450__ (
    .I5(TM0),
    .I4(__503__),
    .I3(__471__),
    .I2(__439__),
    .I1(__535__),
    .I0(__360__),
    .O(__2288__)
  );
  LUT5 #(
    .INIT(32'h14414114)
  ) __6451__ (
    .I4(__311__),
    .I3(__54__),
    .I2(__2__),
    .I1(__343__),
    .I0(TM0),
    .O(__2289__)
  );
  LUT6 #(
    .INIT(64'hff880f0f00000000)
  ) __6452__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__2289__),
    .I2(__2288__),
    .I1(TM0),
    .I0(__42__),
    .O(__2290__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6453__ (
    .I2(TM0),
    .I1(__1709__),
    .I0(DATA_0_13),
    .O(__2291__)
  );
  LUT5 #(
    .INIT(32'h14414114)
  ) __6454__ (
    .I4(__1586__),
    .I3(__1618__),
    .I2(__1650__),
    .I1(__1682__),
    .I0(TM0),
    .O(__2292__)
  );
  LUT6 #(
    .INIT(64'hff88f0f000000000)
  ) __6455__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__2292__),
    .I2(__2291__),
    .I1(TM0),
    .I0(__1554__),
    .O(__2293__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6456__ (
    .I1(RESET),
    .I0(__690__),
    .O(__2294__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6457__ (
    .I1(RESET),
    .I0(__503__),
    .O(__2295__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6458__ (
    .I2(RESET),
    .I1(__562__),
    .I0(__524__),
    .O(__2296__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6459__ (
    .I1(RESET),
    .I0(__298__),
    .O(__2297__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6460__ (
    .I1(RESET),
    .I0(__246__),
    .O(__2298__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6461__ (
    .I5(TM0),
    .I4(__530__),
    .I3(__498__),
    .I2(__434__),
    .I1(__466__),
    .I0(__365__),
    .O(__2299__)
  );
  LUT5 #(
    .INIT(32'h14414114)
  ) __6462__ (
    .I4(__24__),
    .I3(__7__),
    .I2(__306__),
    .I1(__338__),
    .I0(TM0),
    .O(__2300__)
  );
  LUT6 #(
    .INIT(64'hff880f0f00000000)
  ) __6463__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__2300__),
    .I2(__2299__),
    .I1(TM0),
    .I0(__47__),
    .O(__2301__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6464__ (
    .I1(RESET),
    .I0(__863__),
    .O(__2302__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6465__ (
    .I1(RESET),
    .I0(__1545__),
    .O(__2303__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6466__ (
    .I1(TM0),
    .I0(__240__),
    .O(__2304__)
  );
  LUT6 #(
    .INIT(64'h6996966996696996)
  ) __6467__ (
    .I5(TM1),
    .I4(__254__),
    .I3(__193__),
    .I2(__226__),
    .I1(__209__),
    .I0(__2304__),
    .O(__2305__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6468__ (
    .I1(RESET),
    .I0(__123__),
    .O(__2306__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6469__ (
    .I5(TM0),
    .I4(__1237__),
    .I3(__1301__),
    .I2(__1269__),
    .I1(__1205__),
    .I0(__1130__),
    .O(__2307__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6470__ (
    .I5(TM0),
    .I4(__1045__),
    .I3(__1013__),
    .I2(__1109__),
    .I1(__1077__),
    .I0(__981__),
    .O(__2308__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __6471__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__2308__),
    .I0(__2307__),
    .O(__2309__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6472__ (
    .I1(RESET),
    .I0(__623__),
    .O(__2310__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6473__ (
    .I1(TM0),
    .I0(__1332__),
    .O(__2311__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6474__ (
    .I5(TM1),
    .I4(__1387__),
    .I3(__1451__),
    .I2(__1419__),
    .I1(__1483__),
    .I0(TM0),
    .O(__2312__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6475__ (
    .I1(TM0),
    .I0(__1163__),
    .O(__2313__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __6476__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__2313__),
    .I2(__1773__),
    .I1(__2312__),
    .I0(__2311__),
    .O(__2314__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6477__ (
    .I1(TM0),
    .I0(__950__),
    .O(__2315__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6478__ (
    .I5(TM1),
    .I4(__1065__),
    .I3(__1033__),
    .I2(__1001__),
    .I1(__1097__),
    .I0(TM0),
    .O(__2316__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6479__ (
    .I1(TM0),
    .I0(__777__),
    .O(__2317__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6480__ (
    .I5(TM1),
    .I4(__873__),
    .I3(__841__),
    .I2(__809__),
    .I1(__905__),
    .I0(TM0),
    .O(__2318__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __6481__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__2318__),
    .I2(__2317__),
    .I1(__2316__),
    .I0(__2315__),
    .O(__2319__)
  );
  LUT5 #(
    .INIT(32'h14414114)
  ) __6482__ (
    .I4(__344__),
    .I3(__1__),
    .I2(__312__),
    .I1(__22__),
    .I0(TM0),
    .O(__2320__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6483__ (
    .I5(TM0),
    .I4(__185__),
    .I3(__219__),
    .I2(__251__),
    .I1(__153__),
    .I0(__284__),
    .O(__2321__)
  );
  LUT6 #(
    .INIT(64'h00fff8f800000000)
  ) __6484__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__2321__),
    .I2(__2320__),
    .I1(TM0),
    .I0(__144__),
    .O(__2322__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6485__ (
    .I5(TM0),
    .I4(__1110__),
    .I3(__1078__),
    .I2(__1046__),
    .I1(__1014__),
    .I0(__937__),
    .O(__2323__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6486__ (
    .I5(TM0),
    .I4(__854__),
    .I3(__886__),
    .I2(__822__),
    .I1(__918__),
    .I0(__790__),
    .O(__2324__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __6487__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__2324__),
    .I0(__2323__),
    .O(__2325__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6488__ (
    .I1(RESET),
    .I0(__1047__),
    .O(__2326__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6489__ (
    .I2(RESET),
    .I1(__372__),
    .I0(__330__),
    .O(__2327__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6490__ (
    .I2(TM0),
    .I1(__1722__),
    .I0(DATA_0_26),
    .O(__2328__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6491__ (
    .I5(TM1),
    .I4(__1669__),
    .I3(__1573__),
    .I2(__1605__),
    .I1(__1637__),
    .I0(TM0),
    .O(__2329__)
  );
  LUT6 #(
    .INIT(64'hff88f0f000000000)
  ) __6492__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__2329__),
    .I2(__2328__),
    .I1(TM0),
    .I0(__1541__),
    .O(__2330__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6493__ (
    .I1(RESET),
    .I0(__297__),
    .O(__2331__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6494__ (
    .I1(RESET),
    .I0(__628__),
    .O(__2332__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6495__ (
    .I1(RESET),
    .I0(__389__),
    .O(__2333__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6496__ (
    .I1(RESET),
    .I0(__1426__),
    .O(__2334__)
  );
  LUT4 #(
    .INIT(16'h6900)
  ) __6497__ (
    .I3(RESET),
    .I2(__1343__),
    .I1(__1295__),
    .I0(__1327__),
    .O(__2335__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6498__ (
    .I1(RESET),
    .I0(__490__),
    .O(__2336__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6499__ (
    .I1(RESET),
    .I0(__688__),
    .O(__2337__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6500__ (
    .I1(RESET),
    .I0(__264__),
    .O(__2338__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6501__ (
    .I1(RESET),
    .I0(__285__),
    .O(__2339__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6502__ (
    .I1(RESET),
    .I0(__1637__),
    .O(__2340__)
  );
  LUT5 #(
    .INIT(32'h14414114)
  ) __6503__ (
    .I4(__1594__),
    .I3(__1626__),
    .I2(__1690__),
    .I1(__1658__),
    .I0(TM0),
    .O(__2341__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6504__ (
    .I5(TM0),
    .I4(__1402__),
    .I3(__1466__),
    .I2(__1434__),
    .I1(__1498__),
    .I0(__1370__),
    .O(__2342__)
  );
  LUT6 #(
    .INIT(64'h00fff8f800000000)
  ) __6505__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__2342__),
    .I2(__2341__),
    .I1(TM0),
    .I0(__1509__),
    .O(__2343__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6506__ (
    .I1(RESET),
    .I0(__23__),
    .O(__2344__)
  );
  LUT4 #(
    .INIT(16'h6900)
  ) __6507__ (
    .I3(RESET),
    .I2(__347__),
    .I1(__383__),
    .I0(__355__),
    .O(__2345__)
  );
  LUT6 #(
    .INIT(64'h4bb4b44bb44b4bb4)
  ) __6508__ (
    .I5(__198__),
    .I4(__230__),
    .I3(__264__),
    .I2(__164__),
    .I1(TM0),
    .I0(__290__),
    .O(__2346__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6509__ (
    .I1(RESET),
    .I0(__810__),
    .O(__2347__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6510__ (
    .I1(RESET),
    .I0(__41__),
    .O(__2348__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6511__ (
    .I1(RESET),
    .I0(__685__),
    .O(__2349__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6512__ (
    .I1(RESET),
    .I0(__1180__),
    .O(__2350__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6513__ (
    .I1(RESET),
    .I0(__640__),
    .O(__2351__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6514__ (
    .I1(RESET),
    .I0(__870__),
    .O(__2352__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6515__ (
    .I1(RESET),
    .I0(__66__),
    .O(__2353__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6516__ (
    .I1(RESET),
    .I0(__47__),
    .O(__2354__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6517__ (
    .I5(TM0),
    .I4(__639__),
    .I3(__703__),
    .I2(__671__),
    .I1(__735__),
    .I0(__544__),
    .O(__2355__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6518__ (
    .I5(TM0),
    .I4(__479__),
    .I3(__447__),
    .I2(__511__),
    .I1(__543__),
    .I0(__415__),
    .O(__2356__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __6519__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__2356__),
    .I0(__2355__),
    .O(__2357__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6520__ (
    .I1(RESET),
    .I0(__1647__),
    .O(__2358__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6521__ (
    .I1(RESET),
    .I0(__456__),
    .O(__2359__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6522__ (
    .I2(RESET),
    .I1(__1674__),
    .I0(__1716__),
    .O(__2360__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6523__ (
    .I5(TM0),
    .I4(__890__),
    .I3(__922__),
    .I2(__858__),
    .I1(__826__),
    .I0(__741__),
    .O(__2361__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6524__ (
    .I5(TM0),
    .I4(__730__),
    .I3(__634__),
    .I2(__698__),
    .I1(__666__),
    .I0(__602__),
    .O(__2362__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __6525__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__2362__),
    .I0(__2361__),
    .O(__2363__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6526__ (
    .I5(TM0),
    .I4(__1118__),
    .I3(__1086__),
    .I2(__1022__),
    .I1(__1054__),
    .I0(__929__),
    .O(__2364__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6527__ (
    .I5(TM0),
    .I4(__894__),
    .I3(__862__),
    .I2(__830__),
    .I1(__926__),
    .I0(__798__),
    .O(__2365__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __6528__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__2365__),
    .I0(__2364__),
    .O(__2366__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6529__ (
    .I1(RESET),
    .I0(__488__),
    .O(__2367__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6530__ (
    .I1(RESET),
    .I0(__1206__),
    .O(__2368__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6531__ (
    .I1(RESET),
    .I0(__1033__),
    .O(__2369__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6532__ (
    .I1(TM0),
    .I0(__1143__),
    .O(__2370__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6533__ (
    .I5(TM1),
    .I4(__1256__),
    .I3(__1192__),
    .I2(__1224__),
    .I1(__1288__),
    .I0(TM0),
    .O(__2371__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6534__ (
    .I1(TM0),
    .I0(__968__),
    .O(__2372__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __6535__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__2372__),
    .I2(__1907__),
    .I1(__2371__),
    .I0(__2370__),
    .O(__2373__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6536__ (
    .I2(TM0),
    .I1(__1711__),
    .I0(DATA_0_15),
    .O(__2374__)
  );
  LUT5 #(
    .INIT(32'h14414114)
  ) __6537__ (
    .I4(__1648__),
    .I3(__1616__),
    .I2(__1584__),
    .I1(__1680__),
    .I0(TM0),
    .O(__2375__)
  );
  LUT6 #(
    .INIT(64'hff88f0f000000000)
  ) __6538__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__2375__),
    .I2(__2374__),
    .I1(TM0),
    .I0(__1552__),
    .O(__2376__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6539__ (
    .I1(RESET),
    .I0(__1154__),
    .O(__2377__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6540__ (
    .I1(RESET),
    .I0(__626__),
    .O(__2378__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6541__ (
    .I1(RESET),
    .I0(__793__),
    .O(__2379__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6542__ (
    .I1(RESET),
    .I0(__1589__),
    .O(__2380__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6543__ (
    .I1(RESET),
    .I0(__182__),
    .O(__2381__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6544__ (
    .I1(RESET),
    .I0(__1014__),
    .O(__2382__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6545__ (
    .I1(RESET),
    .I0(__1368__),
    .O(__2383__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6546__ (
    .I1(RESET),
    .I0(__124__),
    .O(__2384__)
  );
  LUT6 #(
    .INIT(64'h4bb4b44bb44b4bb4)
  ) __6547__ (
    .I5(__136__),
    .I4(__103__),
    .I3(__167__),
    .I2(__253__),
    .I1(TM0),
    .I0(__286__),
    .O(__2385__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6548__ (
    .I1(TM0),
    .I0(__1337__),
    .O(__2386__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6549__ (
    .I1(TM0),
    .I0(__1158__),
    .O(__2387__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6550__ (
    .I5(TM1),
    .I4(__1254__),
    .I3(__1222__),
    .I2(__1190__),
    .I1(__1286__),
    .I0(TM0),
    .O(__2388__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __6551__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__2388__),
    .I2(__2387__),
    .I1(__2095__),
    .I0(__2386__),
    .O(__2389__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6552__ (
    .I1(RESET),
    .I0(__979__),
    .O(__2390__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6553__ (
    .I2(RESET),
    .I1(__361__),
    .I0(__341__),
    .O(__2391__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6554__ (
    .I5(TM0),
    .I4(__500__),
    .I3(__468__),
    .I2(__436__),
    .I1(__532__),
    .I0(__363__),
    .O(__2392__)
  );
  LUT6 #(
    .INIT(64'hff880f0f00000000)
  ) __6555__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__2003__),
    .I2(__2392__),
    .I1(TM0),
    .I0(__45__),
    .O(__2393__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6556__ (
    .I1(TM0),
    .I0(__72__),
    .O(__2394__)
  );
  LUT5 #(
    .INIT(32'h41141441)
  ) __6557__ (
    .I4(__172__),
    .I3(__134__),
    .I2(__141__),
    .I1(__205__),
    .I0(TM0),
    .O(__2395__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6558__ (
    .I1(TM0),
    .I0(__236__),
    .O(__2396__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __6559__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__2396__),
    .I2(__2395__),
    .I1(__2277__),
    .I0(__2394__),
    .O(__2397__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6560__ (
    .I1(RESET),
    .I0(__771__),
    .O(__2398__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6561__ (
    .I1(TM0),
    .I0(__764__),
    .O(__2399__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6562__ (
    .I5(TM1),
    .I4(__899__),
    .I3(__835__),
    .I2(__867__),
    .I1(__803__),
    .I0(TM0),
    .O(__2400__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6563__ (
    .I1(TM0),
    .I0(__579__),
    .O(__2401__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6564__ (
    .I5(TM1),
    .I4(__675__),
    .I3(__643__),
    .I2(__611__),
    .I1(__707__),
    .I0(TM0),
    .O(__2402__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __6565__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__2402__),
    .I2(__2401__),
    .I1(__2400__),
    .I0(__2399__),
    .O(__2403__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6566__ (
    .I1(RESET),
    .I0(__845__),
    .O(__2404__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6567__ (
    .I1(RESET),
    .I0(__605__),
    .O(__2405__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6568__ (
    .I1(RESET),
    .I0(__414__),
    .O(__2406__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6569__ (
    .I1(TM0),
    .I0(__953__),
    .O(__2407__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6570__ (
    .I5(TM1),
    .I4(__1062__),
    .I3(__1094__),
    .I2(__998__),
    .I1(__1030__),
    .I0(TM0),
    .O(__2408__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6571__ (
    .I1(TM0),
    .I0(__774__),
    .O(__2409__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6572__ (
    .I5(TM1),
    .I4(__870__),
    .I3(__838__),
    .I2(__806__),
    .I1(__902__),
    .I0(TM0),
    .O(__2410__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __6573__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__2410__),
    .I2(__2409__),
    .I1(__2408__),
    .I0(__2407__),
    .O(__2411__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6574__ (
    .I5(TM0),
    .I4(__697__),
    .I3(__665__),
    .I2(__633__),
    .I1(__729__),
    .I0(__550__),
    .O(__2412__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6575__ (
    .I5(TM0),
    .I4(__505__),
    .I3(__473__),
    .I2(__441__),
    .I1(__537__),
    .I0(__409__),
    .O(__2413__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __6576__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__2413__),
    .I0(__2412__),
    .O(__2414__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6577__ (
    .I1(RESET),
    .I0(__1539__),
    .O(__2415__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6578__ (
    .I2(TM0),
    .I1(__1701__),
    .I0(DATA_0_5),
    .O(__2416__)
  );
  LUT6 #(
    .INIT(64'hff88f0f000000000)
  ) __6579__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__2341__),
    .I2(__2416__),
    .I1(TM0),
    .I0(__1562__),
    .O(__2417__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6580__ (
    .I2(RESET),
    .I1(__1485__),
    .I0(__1521__),
    .O(__2418__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6581__ (
    .I1(RESET),
    .I0(__306__),
    .O(__2419__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6582__ (
    .I1(RESET),
    .I0(__1083__),
    .O(__2420__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6583__ (
    .I1(TM0),
    .I0(__117__),
    .O(__2421__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6584__ (
    .I5(TM1),
    .I4(__84__),
    .I3(__321__),
    .I2(__13__),
    .I1(__19__),
    .I0(TM0),
    .O(__2422__)
  );
  LUT5 #(
    .INIT(32'h41141441)
  ) __6585__ (
    .I4(__277__),
    .I3(__178__),
    .I2(__212__),
    .I1(__244__),
    .I0(TM0),
    .O(__2423__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6586__ (
    .I1(TM0),
    .I0(__274__),
    .O(__2424__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __6587__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__2424__),
    .I2(__2423__),
    .I1(__2422__),
    .I0(__2421__),
    .O(__2425__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6588__ (
    .I1(RESET),
    .I0(__412__),
    .O(__2426__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6589__ (
    .I2(RESET),
    .I1(__928__),
    .I0(__926__),
    .O(__2427__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6590__ (
    .I1(RESET),
    .I0(__1191__),
    .O(__2428__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6591__ (
    .I1(RESET),
    .I0(__820__),
    .O(__2429__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6592__ (
    .I1(TM0),
    .I0(__945__),
    .O(__2430__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6593__ (
    .I5(TM1),
    .I4(__1006__),
    .I3(__1038__),
    .I2(__1070__),
    .I1(__1102__),
    .I0(TM0),
    .O(__2431__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6594__ (
    .I1(TM0),
    .I0(__782__),
    .O(__2432__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __6595__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__2432__),
    .I2(__2238__),
    .I1(__2431__),
    .I0(__2430__),
    .O(__2433__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6596__ (
    .I1(RESET),
    .I0(__1547__),
    .O(__2434__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6597__ (
    .I1(RESET),
    .I0(__1463__),
    .O(__2435__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6598__ (
    .I1(RESET),
    .I0(__1217__),
    .O(__2436__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6599__ (
    .I2(RESET),
    .I1(__708__),
    .I0(__762__),
    .O(__2437__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6600__ (
    .I1(RESET),
    .I0(__12__),
    .O(__2438__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6601__ (
    .I1(TM0),
    .I0(__563__),
    .O(__2439__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6602__ (
    .I5(TM1),
    .I4(__716__),
    .I3(__684__),
    .I2(__620__),
    .I1(__652__),
    .I0(TM0),
    .O(__2440__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6603__ (
    .I1(TM0),
    .I0(__396__),
    .O(__2441__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __6604__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__2441__),
    .I2(__2189__),
    .I1(__2440__),
    .I0(__2439__),
    .O(__2442__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6605__ (
    .I1(RESET),
    .I0(__1046__),
    .O(__2443__)
  );
  LUT4 #(
    .INIT(16'h6900)
  ) __6606__ (
    .I3(RESET),
    .I2(__1519__),
    .I1(__1487__),
    .I0(__1535__),
    .O(__2444__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6607__ (
    .I1(RESET),
    .I0(__511__),
    .O(__2445__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6608__ (
    .I1(TM0),
    .I0(__382__),
    .O(__2446__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6609__ (
    .I5(TM1),
    .I4(__481__),
    .I3(__417__),
    .I2(__449__),
    .I1(__513__),
    .I0(TM0),
    .O(__2447__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6610__ (
    .I1(TM0),
    .I0(__116__),
    .O(__2448__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __6611__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__2448__),
    .I2(__2422__),
    .I1(__2447__),
    .I0(__2446__),
    .O(__2449__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6612__ (
    .I2(RESET),
    .I1(__749__),
    .I0(__721__),
    .O(__2450__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6613__ (
    .I1(TM0),
    .I0(__1333__),
    .O(__2451__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6614__ (
    .I5(TM1),
    .I4(__1450__),
    .I3(__1418__),
    .I2(__1386__),
    .I1(__1482__),
    .I0(TM0),
    .O(__2452__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6615__ (
    .I1(TM0),
    .I0(__1162__),
    .O(__2453__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __6616__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__2453__),
    .I2(__1817__),
    .I1(__2452__),
    .I0(__2451__),
    .O(__2454__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6617__ (
    .I1(RESET),
    .I0(__1606__),
    .O(__2455__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6618__ (
    .I1(RESET),
    .I0(__1166__),
    .O(__2456__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6619__ (
    .I1(RESET),
    .I0(__786__),
    .O(__2457__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6620__ (
    .I1(RESET),
    .I0(__1228__),
    .O(__2458__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6621__ (
    .I5(TM0),
    .I4(__730__),
    .I3(__634__),
    .I2(__698__),
    .I1(__666__),
    .I0(__549__),
    .O(__2459__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6622__ (
    .I5(TM0),
    .I4(__506__),
    .I3(__474__),
    .I2(__442__),
    .I1(__538__),
    .I0(__410__),
    .O(__2460__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __6623__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__2460__),
    .I0(__2459__),
    .O(__2461__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __6624__ (
    .I1(RESET),
    .I0(__384__),
    .O(__2462__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6625__ (
    .I1(RESET),
    .I0(__631__),
    .O(__2463__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6626__ (
    .I1(RESET),
    .I0(__1388__),
    .O(__2464__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6627__ (
    .I1(RESET),
    .I0(__1352__),
    .O(__2465__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6628__ (
    .I5(TM0),
    .I4(__1458__),
    .I3(__1394__),
    .I2(__1426__),
    .I1(__1490__),
    .I0(__1325__),
    .O(__2466__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6629__ (
    .I5(TM0),
    .I4(__1298__),
    .I3(__1266__),
    .I2(__1234__),
    .I1(__1202__),
    .I0(__1170__),
    .O(__2467__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __6630__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__2467__),
    .I0(__2466__),
    .O(__2468__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6631__ (
    .I1(TM0),
    .I0(__1139__),
    .O(__2469__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6632__ (
    .I1(TM0),
    .I0(__972__),
    .O(__2470__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6633__ (
    .I5(TM1),
    .I4(__1036__),
    .I3(__1004__),
    .I2(__1100__),
    .I1(__1068__),
    .I0(TM0),
    .O(__2471__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __6634__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__2471__),
    .I2(__2470__),
    .I1(__1850__),
    .I0(__2469__),
    .O(__2472__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6635__ (
    .I1(RESET),
    .I0(__453__),
    .O(__2473__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6636__ (
    .I1(RESET),
    .I0(__585__),
    .O(__2474__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6637__ (
    .I1(RESET),
    .I0(__1224__),
    .O(__2475__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6638__ (
    .I2(TM0),
    .I1(__1710__),
    .I0(DATA_0_14),
    .O(__2476__)
  );
  LUT5 #(
    .INIT(32'h14414114)
  ) __6639__ (
    .I4(__1681__),
    .I3(__1585__),
    .I2(__1649__),
    .I1(__1617__),
    .I0(TM0),
    .O(__2477__)
  );
  LUT6 #(
    .INIT(64'hff88f0f000000000)
  ) __6640__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__2477__),
    .I2(__2476__),
    .I1(TM0),
    .I0(__1553__),
    .O(__2478__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6641__ (
    .I1(RESET),
    .I0(__411__),
    .O(__2479__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6642__ (
    .I1(RESET),
    .I0(__1279__),
    .O(__2480__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6643__ (
    .I2(RESET),
    .I1(__1095__),
    .I0(__1143__),
    .O(__2481__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6644__ (
    .I2(RESET),
    .I1(__537__),
    .I0(__549__),
    .O(__2482__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6645__ (
    .I1(RESET),
    .I0(__1081__),
    .O(__2483__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6646__ (
    .I1(TM0),
    .I0(__571__),
    .O(__2484__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6647__ (
    .I5(TM1),
    .I4(__676__),
    .I3(__644__),
    .I2(__612__),
    .I1(__708__),
    .I0(TM0),
    .O(__2485__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6648__ (
    .I1(TM0),
    .I0(__388__),
    .O(__2486__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6649__ (
    .I5(TM1),
    .I4(__420__),
    .I3(__484__),
    .I2(__452__),
    .I1(__516__),
    .I0(TM0),
    .O(__2487__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __6650__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__2487__),
    .I2(__2486__),
    .I1(__2485__),
    .I0(__2484__),
    .O(__2488__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6651__ (
    .I1(RESET),
    .I0(__827__),
    .O(__2489__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6652__ (
    .I2(RESET),
    .I1(__515__),
    .I0(__571__),
    .O(__2490__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6653__ (
    .I1(RESET),
    .I0(__126__),
    .O(__2491__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6654__ (
    .I1(RESET),
    .I0(__677__),
    .O(__2492__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6655__ (
    .I1(RESET),
    .I0(__987__),
    .O(__2493__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6656__ (
    .I2(RESET),
    .I1(__156__),
    .I0(__165__),
    .O(__2494__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6657__ (
    .I1(RESET),
    .I0(__394__),
    .O(__2495__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6658__ (
    .I1(RESET),
    .I0(__1452__),
    .O(__2496__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6659__ (
    .I1(RESET),
    .I0(__643__),
    .O(__2497__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6660__ (
    .I1(RESET),
    .I0(__227__),
    .O(__2498__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6661__ (
    .I1(TM0),
    .I0(__947__),
    .O(__2499__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6662__ (
    .I1(TM0),
    .I0(__780__),
    .O(__2500__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6663__ (
    .I5(TM1),
    .I4(__876__),
    .I3(__844__),
    .I2(__812__),
    .I1(__908__),
    .I0(TM0),
    .O(__2501__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __6664__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__2501__),
    .I2(__2500__),
    .I1(__2471__),
    .I0(__2499__),
    .O(__2502__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6665__ (
    .I1(RESET),
    .I0(__1419__),
    .O(__2503__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6666__ (
    .I1(TM0),
    .I0(__752__),
    .O(__2504__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6667__ (
    .I5(TM1),
    .I4(__815__),
    .I3(__879__),
    .I2(__847__),
    .I1(__911__),
    .I0(TM0),
    .O(__2505__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6668__ (
    .I1(TM0),
    .I0(__591__),
    .O(__2506__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6669__ (
    .I5(TM1),
    .I4(__687__),
    .I3(__655__),
    .I2(__623__),
    .I1(__719__),
    .I0(TM0),
    .O(__2507__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __6670__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__2507__),
    .I2(__2506__),
    .I1(__2505__),
    .I0(__2504__),
    .O(__2508__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6671__ (
    .I1(RESET),
    .I0(__994__),
    .O(__2509__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6672__ (
    .I1(TM0),
    .I0(__133__),
    .O(__2510__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6673__ (
    .I5(TM1),
    .I4(__95__),
    .I3(__59__),
    .I2(__49__),
    .I1(__326__),
    .I0(TM0),
    .O(__2511__)
  );
  LUT5 #(
    .INIT(32'h41141441)
  ) __6674__ (
    .I4(__260__),
    .I3(__292__),
    .I2(__194__),
    .I1(__227__),
    .I0(TM0),
    .O(__2512__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __6675__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__2512__),
    .I2(__1892__),
    .I1(__2511__),
    .I0(__2510__),
    .O(__2513__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6676__ (
    .I1(RESET),
    .I0(__1612__),
    .O(__2514__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6677__ (
    .I1(TM0),
    .I0(__68__),
    .O(__2515__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6678__ (
    .I5(TM1),
    .I4(__94__),
    .I3(__66__),
    .I2(__58__),
    .I1(__329__),
    .I0(TM0),
    .O(__2516__)
  );
  LUT5 #(
    .INIT(32'h41141441)
  ) __6679__ (
    .I4(__254__),
    .I3(__193__),
    .I2(__226__),
    .I1(__209__),
    .I0(TM0),
    .O(__2517__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __6680__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__2517__),
    .I2(__2304__),
    .I1(__2516__),
    .I0(__2515__),
    .O(__2518__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6681__ (
    .I1(RESET),
    .I0(__880__),
    .O(__2519__)
  );
  LUT6 #(
    .INIT(64'h6996966996696996)
  ) __6682__ (
    .I5(TM1),
    .I4(__277__),
    .I3(__178__),
    .I2(__212__),
    .I1(__244__),
    .I0(__2424__),
    .O(__2520__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6683__ (
    .I2(RESET),
    .I1(__747__),
    .I0(__723__),
    .O(__2521__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6684__ (
    .I1(RESET),
    .I0(__893__),
    .O(__2522__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6685__ (
    .I1(RESET),
    .I0(__1634__),
    .O(__2523__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6686__ (
    .I2(RESET),
    .I1(__343__),
    .I0(__359__),
    .O(__2524__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6687__ (
    .I1(RESET),
    .I0(__1422__),
    .O(__2525__)
  );
  LUT6 #(
    .INIT(64'h6996966996696996)
  ) __6688__ (
    .I5(TM1),
    .I4(__223__),
    .I3(__191__),
    .I2(__288__),
    .I1(__257__),
    .I0(__2260__),
    .O(__2526__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6689__ (
    .I5(TM0),
    .I4(__1458__),
    .I3(__1394__),
    .I2(__1426__),
    .I1(__1490__),
    .I0(__1362__),
    .O(__2527__)
  );
  LUT6 #(
    .INIT(64'h00fff8f800000000)
  ) __6690__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__2527__),
    .I2(__2292__),
    .I1(TM0),
    .I0(__1517__),
    .O(__2528__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6691__ (
    .I2(RESET),
    .I1(__900__),
    .I0(__954__),
    .O(__2529__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6692__ (
    .I1(RESET),
    .I0(__1064__),
    .O(__2530__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6693__ (
    .I2(RESET),
    .I1(__322__),
    .I0(__380__),
    .O(__2531__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6694__ (
    .I1(RESET),
    .I0(__1421__),
    .O(__2532__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6695__ (
    .I1(RESET),
    .I0(__299__),
    .O(__2533__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6696__ (
    .I5(TM0),
    .I4(__1045__),
    .I3(__1013__),
    .I2(__1109__),
    .I1(__1077__),
    .I0(__938__),
    .O(__2534__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6697__ (
    .I5(TM0),
    .I4(__917__),
    .I3(__853__),
    .I2(__885__),
    .I1(__821__),
    .I0(__789__),
    .O(__2535__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __6698__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__2535__),
    .I0(__2534__),
    .O(__2536__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6699__ (
    .I1(RESET),
    .I0(__139__),
    .O(__2537__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6700__ (
    .I1(RESET),
    .I0(__1546__),
    .O(__2538__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6701__ (
    .I2(RESET),
    .I1(__907__),
    .I0(__947__),
    .O(__2539__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6702__ (
    .I1(RESET),
    .I0(__656__),
    .O(__2540__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6703__ (
    .I1(RESET),
    .I0(__257__),
    .O(__2541__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6704__ (
    .I1(RESET),
    .I0(__1222__),
    .O(__2542__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6705__ (
    .I1(RESET),
    .I0(__1385__),
    .O(__2543__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6706__ (
    .I1(RESET),
    .I0(__818__),
    .O(__2544__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6707__ (
    .I1(RESET),
    .I0(__247__),
    .O(__2545__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6708__ (
    .I2(RESET),
    .I1(__383__),
    .I0(__351__),
    .O(__2546__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6709__ (
    .I1(RESET),
    .I0(__425__),
    .O(__2547__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6710__ (
    .I1(RESET),
    .I0(__1392__),
    .O(__2548__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6711__ (
    .I1(RESET),
    .I0(__1449__),
    .O(__2549__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6712__ (
    .I5(TM0),
    .I4(__1276__),
    .I3(__1308__),
    .I2(__1212__),
    .I1(__1244__),
    .I0(__1123__),
    .O(__2550__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6713__ (
    .I5(TM0),
    .I4(__1084__),
    .I3(__1020__),
    .I2(__1116__),
    .I1(__1052__),
    .I0(__988__),
    .O(__2551__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __6714__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__2551__),
    .I0(__2550__),
    .O(__2552__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6715__ (
    .I1(RESET),
    .I0(__1434__),
    .O(__2553__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6716__ (
    .I1(RESET),
    .I0(__1058__),
    .O(__2554__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6717__ (
    .I1(RESET),
    .I0(__1373__),
    .O(__2555__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6718__ (
    .I1(RESET),
    .I0(__213__),
    .O(__2556__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6719__ (
    .I5(TM0),
    .I4(__1049__),
    .I3(__1017__),
    .I2(__1081__),
    .I1(__1113__),
    .I0(__934__),
    .O(__2557__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6720__ (
    .I5(TM0),
    .I4(__857__),
    .I3(__825__),
    .I2(__889__),
    .I1(__921__),
    .I0(__793__),
    .O(__2558__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __6721__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__2558__),
    .I0(__2557__),
    .O(__2559__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6722__ (
    .I1(RESET),
    .I0(__62__),
    .O(__2560__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6723__ (
    .I2(RESET),
    .I1(__763__),
    .I0(__707__),
    .O(__2561__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6724__ (
    .I5(TM0),
    .I4(__1084__),
    .I3(__1020__),
    .I2(__1116__),
    .I1(__1052__),
    .I0(__931__),
    .O(__2562__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6725__ (
    .I5(TM0),
    .I4(__828__),
    .I3(__892__),
    .I2(__860__),
    .I1(__924__),
    .I0(__796__),
    .O(__2563__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __6726__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__2563__),
    .I0(__2562__),
    .O(__2564__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6727__ (
    .I1(RESET),
    .I0(__1651__),
    .O(__2565__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6728__ (
    .I1(TM0),
    .I0(__755__),
    .O(__2566__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6729__ (
    .I1(TM0),
    .I0(__588__),
    .O(__2567__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __6730__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__2567__),
    .I2(__2440__),
    .I1(__2501__),
    .I0(__2566__),
    .O(__2568__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6731__ (
    .I5(TM0),
    .I4(__694__),
    .I3(__662__),
    .I2(__726__),
    .I1(__630__),
    .I0(__553__),
    .O(__2569__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6732__ (
    .I5(TM0),
    .I4(__470__),
    .I3(__534__),
    .I2(__502__),
    .I1(__438__),
    .I0(__406__),
    .O(__2570__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __6733__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__2570__),
    .I0(__2569__),
    .O(__2571__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6734__ (
    .I1(RESET),
    .I0(__1417__),
    .O(__2572__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6735__ (
    .I1(RESET),
    .I0(__588__),
    .O(__2573__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6736__ (
    .I1(RESET),
    .I0(__1408__),
    .O(__2574__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6737__ (
    .I1(RESET),
    .I0(__1273__),
    .O(__2575__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6738__ (
    .I1(TM0),
    .I0(__241__),
    .O(__2576__)
  );
  LUT6 #(
    .INIT(64'h6996966996696996)
  ) __6739__ (
    .I5(TM1),
    .I4(__189__),
    .I3(__255__),
    .I2(__221__),
    .I1(__259__),
    .I0(__2576__),
    .O(__2577__)
  );
  LUT5 #(
    .INIT(32'h14414114)
  ) __6740__ (
    .I4(__318__),
    .I3(__20__),
    .I2(__14__),
    .I1(__350__),
    .I0(TM0),
    .O(__2578__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6741__ (
    .I5(TM0),
    .I4(__245__),
    .I3(__217__),
    .I2(__183__),
    .I1(__151__),
    .I0(__278__),
    .O(__2579__)
  );
  LUT6 #(
    .INIT(64'h00fff8f800000000)
  ) __6742__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__2579__),
    .I2(__2578__),
    .I1(TM0),
    .I0(__150__),
    .O(__2580__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6743__ (
    .I1(RESET),
    .I0(__1042__),
    .O(__2581__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6744__ (
    .I1(RESET),
    .I0(__496__),
    .O(__2582__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6745__ (
    .I1(RESET),
    .I0(__1188__),
    .O(__2583__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6746__ (
    .I1(RESET),
    .I0(__636__),
    .O(__2584__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6747__ (
    .I2(RESET),
    .I1(__521__),
    .I0(__565__),
    .O(__2585__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6748__ (
    .I2(RESET),
    .I1(__1708__),
    .I0(__1682__),
    .O(__2586__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6749__ (
    .I2(RESET),
    .I1(__1689__),
    .I0(__1701__),
    .O(__2587__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6750__ (
    .I1(RESET),
    .I0(__58__),
    .O(__2588__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6751__ (
    .I1(RESET),
    .I0(__1448__),
    .O(__2589__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6752__ (
    .I1(RESET),
    .I0(__1005__),
    .O(__2590__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6753__ (
    .I5(TM0),
    .I4(__1209__),
    .I3(__1241__),
    .I2(__1273__),
    .I1(__1305__),
    .I0(__1126__),
    .O(__2591__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6754__ (
    .I5(TM0),
    .I4(__1049__),
    .I3(__1017__),
    .I2(__1081__),
    .I1(__1113__),
    .I0(__985__),
    .O(__2592__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __6755__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__2592__),
    .I0(__2591__),
    .O(__2593__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6756__ (
    .I1(RESET),
    .I0(__1591__),
    .O(__2594__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6757__ (
    .I1(RESET),
    .I0(__1445__),
    .O(__2595__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6758__ (
    .I1(RESET),
    .I0(__769__),
    .O(__2596__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6759__ (
    .I1(RESET),
    .I0(__1264__),
    .O(__2597__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6760__ (
    .I1(RESET),
    .I0(__1156__),
    .O(__2598__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6761__ (
    .I1(RESET),
    .I0(__842__),
    .O(__2599__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6762__ (
    .I1(RESET),
    .I0(__1624__),
    .O(__2600__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6763__ (
    .I2(RESET),
    .I1(__1515__),
    .I0(__1491__),
    .O(__2601__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6764__ (
    .I1(RESET),
    .I0(__867__),
    .O(__2602__)
  );
  LUT4 #(
    .INIT(16'h6900)
  ) __6765__ (
    .I3(RESET),
    .I2(__1151__),
    .I1(__1115__),
    .I0(__1123__),
    .O(__2603__)
  );
  LUT6 #(
    .INIT(64'h4bb4b44bb44b4bb4)
  ) __6766__ (
    .I5(__245__),
    .I4(__217__),
    .I3(__183__),
    .I2(__151__),
    .I1(TM0),
    .I0(__278__),
    .O(__2604__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6767__ (
    .I1(RESET),
    .I0(__510__),
    .O(__2605__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6768__ (
    .I2(RESET),
    .I1(__758__),
    .I0(__712__),
    .O(__2606__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6769__ (
    .I2(RESET),
    .I1(__1117__),
    .I0(__1121__),
    .O(__2607__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6770__ (
    .I1(RESET),
    .I0(__251__),
    .O(__2608__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6771__ (
    .I2(TM0),
    .I1(__1702__),
    .I0(DATA_0_6),
    .O(__2609__)
  );
  LUT5 #(
    .INIT(32'h14414114)
  ) __6772__ (
    .I4(__1657__),
    .I3(__1625__),
    .I2(__1593__),
    .I1(__1689__),
    .I0(TM0),
    .O(__2610__)
  );
  LUT6 #(
    .INIT(64'hff88f0f000000000)
  ) __6773__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__2610__),
    .I2(__2609__),
    .I1(TM0),
    .I0(__1561__),
    .O(__2611__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6774__ (
    .I1(RESET),
    .I0(__217__),
    .O(__2612__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6775__ (
    .I1(TM0),
    .I0(__568__),
    .O(__2613__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6776__ (
    .I5(TM1),
    .I4(__679__),
    .I3(__647__),
    .I2(__615__),
    .I1(__711__),
    .I0(TM0),
    .O(__2614__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6777__ (
    .I1(TM0),
    .I0(__391__),
    .O(__2615__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6778__ (
    .I5(TM1),
    .I4(__487__),
    .I3(__455__),
    .I2(__423__),
    .I1(__519__),
    .I0(TM0),
    .O(__2616__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __6779__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__2616__),
    .I2(__2615__),
    .I1(__2614__),
    .I0(__2613__),
    .O(__2617__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6780__ (
    .I1(RESET),
    .I0(__1060__),
    .O(__2618__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6781__ (
    .I1(RESET),
    .I0(__1016__),
    .O(__2619__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6782__ (
    .I1(RESET),
    .I0(__90__),
    .O(__2620__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6783__ (
    .I1(RESET),
    .I0(__996__),
    .O(__2621__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6784__ (
    .I2(RESET),
    .I1(__1509__),
    .I0(__1497__),
    .O(__2622__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6785__ (
    .I1(RESET),
    .I0(__697__),
    .O(__2623__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6786__ (
    .I1(RESET),
    .I0(__999__),
    .O(__2624__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6787__ (
    .I1(RESET),
    .I0(__1652__),
    .O(__2625__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6788__ (
    .I1(RESET),
    .I0(__314__),
    .O(__2626__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6789__ (
    .I1(RESET),
    .I0(__1239__),
    .O(__2627__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6790__ (
    .I1(RESET),
    .I0(__1658__),
    .O(__2628__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6791__ (
    .I1(RESET),
    .I0(__15__),
    .O(__2629__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6792__ (
    .I1(RESET),
    .I0(__852__),
    .O(__2630__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6793__ (
    .I1(RESET),
    .I0(__778__),
    .O(__2631__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6794__ (
    .I5(TM0),
    .I4(__917__),
    .I3(__853__),
    .I2(__885__),
    .I1(__821__),
    .I0(__746__),
    .O(__2632__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6795__ (
    .I5(TM0),
    .I4(__693__),
    .I3(__629__),
    .I2(__725__),
    .I1(__661__),
    .I0(__597__),
    .O(__2633__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __6796__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__2633__),
    .I0(__2632__),
    .O(__2634__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6797__ (
    .I1(RESET),
    .I0(__472__),
    .O(__2635__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6798__ (
    .I1(RESET),
    .I0(__49__),
    .O(__2636__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6799__ (
    .I1(TM0),
    .I0(__118__),
    .O(__2637__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6800__ (
    .I5(TM1),
    .I4(__83__),
    .I3(__18__),
    .I2(__12__),
    .I1(__324__),
    .I0(TM0),
    .O(__2638__)
  );
  LUT5 #(
    .INIT(32'h41141441)
  ) __6801__ (
    .I4(__211__),
    .I3(__243__),
    .I2(__276__),
    .I1(__177__),
    .I0(TM0),
    .O(__2639__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6802__ (
    .I1(TM0),
    .I0(__271__),
    .O(__2640__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __6803__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__2640__),
    .I2(__2639__),
    .I1(__2638__),
    .I0(__2637__),
    .O(__2641__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6804__ (
    .I1(RESET),
    .I0(__1054__),
    .O(__2642__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6805__ (
    .I2(RESET),
    .I1(__718__),
    .I0(__752__),
    .O(__2643__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6806__ (
    .I1(RESET),
    .I0(__973__),
    .O(__2644__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6807__ (
    .I1(TM0),
    .I0(__754__),
    .O(__2645__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6808__ (
    .I5(TM1),
    .I4(__877__),
    .I3(__845__),
    .I2(__813__),
    .I1(__909__),
    .I0(TM0),
    .O(__2646__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6809__ (
    .I1(TM0),
    .I0(__589__),
    .O(__2647__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6810__ (
    .I5(TM1),
    .I4(__685__),
    .I3(__653__),
    .I2(__621__),
    .I1(__717__),
    .I0(TM0),
    .O(__2648__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __6811__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__2648__),
    .I2(__2647__),
    .I1(__2646__),
    .I0(__2645__),
    .O(__2649__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6812__ (
    .I2(RESET),
    .I1(__1482__),
    .I0(__1524__),
    .O(__2650__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6813__ (
    .I2(RESET),
    .I1(__542__),
    .I0(__544__),
    .O(__2651__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6814__ (
    .I1(RESET),
    .I0(__887__),
    .O(__2652__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6815__ (
    .I1(RESET),
    .I0(__35__),
    .O(__2653__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6816__ (
    .I1(RESET),
    .I0(__477__),
    .O(__2654__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6817__ (
    .I1(TM0),
    .I0(__1532__),
    .O(__2655__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6818__ (
    .I5(TM1),
    .I4(__1635__),
    .I3(__1603__),
    .I2(__1571__),
    .I1(__1667__),
    .I0(TM0),
    .O(__2656__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6819__ (
    .I1(TM0),
    .I0(__1347__),
    .O(__2657__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6820__ (
    .I5(TM1),
    .I4(__1475__),
    .I3(__1443__),
    .I2(__1379__),
    .I1(__1411__),
    .I0(TM0),
    .O(__2658__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __6821__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__2658__),
    .I2(__2657__),
    .I1(__2656__),
    .I0(__2655__),
    .O(__2659__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6822__ (
    .I1(RESET),
    .I0(__1067__),
    .O(__2660__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6823__ (
    .I1(RESET),
    .I0(__661__),
    .O(__2661__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6824__ (
    .I1(RESET),
    .I0(__99__),
    .O(__2662__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6825__ (
    .I1(RESET),
    .I0(__1218__),
    .O(__2663__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6826__ (
    .I1(RESET),
    .I0(__847__),
    .O(__2664__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6827__ (
    .I1(RESET),
    .I0(__964__),
    .O(__2665__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6828__ (
    .I2(RESET),
    .I1(__337__),
    .I0(__365__),
    .O(__2666__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6829__ (
    .I1(RESET),
    .I0(__1633__),
    .O(__2667__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6830__ (
    .I1(TM0),
    .I0(__1137__),
    .O(__2668__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6831__ (
    .I5(TM1),
    .I4(__1230__),
    .I3(__1198__),
    .I2(__1262__),
    .I1(__1294__),
    .I0(TM0),
    .O(__2669__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6832__ (
    .I1(TM0),
    .I0(__974__),
    .O(__2670__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __6833__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__2670__),
    .I2(__2431__),
    .I1(__2669__),
    .I0(__2668__),
    .O(__2671__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6834__ (
    .I1(TM0),
    .I0(__1340__),
    .O(__2672__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6835__ (
    .I1(TM0),
    .I0(__1155__),
    .O(__2673__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __6836__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__2673__),
    .I2(__2026__),
    .I1(__2658__),
    .I0(__2672__),
    .O(__2674__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6837__ (
    .I1(RESET),
    .I0(__1194__),
    .O(__2675__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6838__ (
    .I5(TM0),
    .I4(__1463__),
    .I3(__1431__),
    .I2(__1399__),
    .I1(__1495__),
    .I0(__1320__),
    .O(__2676__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6839__ (
    .I5(TM0),
    .I4(__1271__),
    .I3(__1239__),
    .I2(__1207__),
    .I1(__1303__),
    .I0(__1175__),
    .O(__2677__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __6840__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__2677__),
    .I0(__2676__),
    .O(__2678__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6841__ (
    .I1(TM0),
    .I0(__948__),
    .O(__2679__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6842__ (
    .I1(TM0),
    .I0(__779__),
    .O(__2680__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6843__ (
    .I5(TM1),
    .I4(__811__),
    .I3(__875__),
    .I2(__843__),
    .I1(__907__),
    .I0(TM0),
    .O(__2681__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __6844__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__2681__),
    .I2(__2680__),
    .I1(__1775__),
    .I0(__2679__),
    .O(__2682__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6845__ (
    .I1(RESET),
    .I0(__209__),
    .O(__2683__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6846__ (
    .I2(RESET),
    .I1(__1138__),
    .I0(__1100__),
    .O(__2684__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6847__ (
    .I1(RESET),
    .I0(__1649__),
    .O(__2685__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6848__ (
    .I1(RESET),
    .I0(__1471__),
    .O(__2686__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6849__ (
    .I1(RESET),
    .I0(__607__),
    .O(__2687__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6850__ (
    .I1(RESET),
    .I0(__1431__),
    .O(__2688__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6851__ (
    .I1(RESET),
    .I0(__1213__),
    .O(__2689__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6852__ (
    .I1(RESET),
    .I0(__813__),
    .O(__2690__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6853__ (
    .I1(TM0),
    .I0(__115__),
    .O(__2691__)
  );
  LUT5 #(
    .INIT(32'h41141441)
  ) __6854__ (
    .I4(__189__),
    .I3(__255__),
    .I2(__221__),
    .I1(__259__),
    .I0(TM0),
    .O(__2692__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __6855__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__2692__),
    .I2(__2576__),
    .I1(__1750__),
    .I0(__2691__),
    .O(__2693__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6856__ (
    .I1(RESET),
    .I0(__798__),
    .O(__2694__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6857__ (
    .I1(RESET),
    .I0(__1646__),
    .O(__2695__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6858__ (
    .I1(RESET),
    .I0(__1564__),
    .O(__2696__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6859__ (
    .I1(RESET),
    .I0(__641__),
    .O(__2697__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6860__ (
    .I2(RESET),
    .I1(__709__),
    .I0(__761__),
    .O(__2698__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6861__ (
    .I5(TM0),
    .I4(__690__),
    .I3(__658__),
    .I2(__626__),
    .I1(__722__),
    .I0(__557__),
    .O(__2699__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6862__ (
    .I5(TM0),
    .I4(__530__),
    .I3(__498__),
    .I2(__434__),
    .I1(__466__),
    .I0(__402__),
    .O(__2700__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __6863__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__2700__),
    .I0(__2699__),
    .O(__2701__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6864__ (
    .I1(RESET),
    .I0(__681__),
    .O(__2702__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6865__ (
    .I2(RESET),
    .I1(__711__),
    .I0(__759__),
    .O(__2703__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6866__ (
    .I1(RESET),
    .I0(__602__),
    .O(__2704__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6867__ (
    .I1(RESET),
    .I0(__969__),
    .O(__2705__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6868__ (
    .I2(RESET),
    .I1(__1495__),
    .I0(__1511__),
    .O(__2706__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6869__ (
    .I1(RESET),
    .I0(__583__),
    .O(__2707__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6870__ (
    .I1(TM0),
    .I0(__1145__),
    .O(__2708__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6871__ (
    .I1(TM0),
    .I0(__966__),
    .O(__2709__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __6872__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__2709__),
    .I2(__2408__),
    .I1(__2388__),
    .I0(__2708__),
    .O(__2710__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6873__ (
    .I1(RESET),
    .I0(__1425__),
    .O(__2711__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6874__ (
    .I2(RESET),
    .I1(__1106__),
    .I0(__1132__),
    .O(__2712__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6875__ (
    .I1(TM0),
    .I0(__564__),
    .O(__2713__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6876__ (
    .I5(TM1),
    .I4(__619__),
    .I3(__715__),
    .I2(__651__),
    .I1(__683__),
    .I0(TM0),
    .O(__2714__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6877__ (
    .I1(TM0),
    .I0(__395__),
    .O(__2715__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6878__ (
    .I5(TM1),
    .I4(__491__),
    .I3(__459__),
    .I2(__427__),
    .I1(__523__),
    .I0(TM0),
    .O(__2716__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __6879__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__2716__),
    .I2(__2715__),
    .I1(__2714__),
    .I0(__2713__),
    .O(__2717__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6880__ (
    .I2(RESET),
    .I1(__918__),
    .I0(__936__),
    .O(__2718__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6881__ (
    .I5(TM0),
    .I4(__1085__),
    .I3(__1053__),
    .I2(__1021__),
    .I1(__1117__),
    .I0(__930__),
    .O(__2719__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6882__ (
    .I5(TM0),
    .I4(__925__),
    .I3(__829__),
    .I2(__861__),
    .I1(__893__),
    .I0(__797__),
    .O(__2720__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __6883__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__2720__),
    .I0(__2719__),
    .O(__2721__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6884__ (
    .I1(RESET),
    .I0(__1004__),
    .O(__2722__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6885__ (
    .I2(RESET),
    .I1(__935__),
    .I0(__919__),
    .O(__2723__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6886__ (
    .I1(RESET),
    .I0(__1625__),
    .O(__2724__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6887__ (
    .I2(RESET),
    .I1(__557__),
    .I0(__529__),
    .O(__2725__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6888__ (
    .I1(RESET),
    .I0(__61__),
    .O(__2726__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __6889__ (
    .I2(TM0),
    .I1(__1717__),
    .I0(DATA_0_21),
    .O(__2727__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6890__ (
    .I5(TM1),
    .I4(__1642__),
    .I3(__1610__),
    .I2(__1578__),
    .I1(__1674__),
    .I0(TM0),
    .O(__2728__)
  );
  LUT6 #(
    .INIT(64'hff88f0f000000000)
  ) __6891__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__2728__),
    .I2(__2727__),
    .I1(TM0),
    .I0(__1546__),
    .O(__2729__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6892__ (
    .I1(RESET),
    .I0(__444__),
    .O(__2730__)
  );
  LUT6 #(
    .INIT(64'h4bb4b44bb44b4bb4)
  ) __6893__ (
    .I5(__218__),
    .I4(__250__),
    .I3(__152__),
    .I2(__184__),
    .I1(TM0),
    .I0(__283__),
    .O(__2731__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6894__ (
    .I5(TM0),
    .I4(__1073__),
    .I3(__1041__),
    .I2(__1009__),
    .I1(__1105__),
    .I0(__942__),
    .O(__2732__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6895__ (
    .I5(TM0),
    .I4(__881__),
    .I3(__849__),
    .I2(__817__),
    .I1(__913__),
    .I0(__785__),
    .O(__2733__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __6896__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__2733__),
    .I0(__2732__),
    .O(__2734__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6897__ (
    .I5(TM0),
    .I4(__895__),
    .I3(__863__),
    .I2(__831__),
    .I1(__927__),
    .I0(__736__),
    .O(__2735__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6898__ (
    .I5(TM0),
    .I4(__639__),
    .I3(__703__),
    .I2(__671__),
    .I1(__735__),
    .I0(__607__),
    .O(__2736__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __6899__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__2736__),
    .I0(__2735__),
    .O(__2737__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6900__ (
    .I1(RESET),
    .I0(__1617__),
    .O(__2738__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6901__ (
    .I2(RESET),
    .I1(__1505__),
    .I0(__1501__),
    .O(__2739__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6902__ (
    .I2(RESET),
    .I1(__734__),
    .I0(__736__),
    .O(__2740__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6903__ (
    .I1(RESET),
    .I0(__460__),
    .O(__2741__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6904__ (
    .I1(RESET),
    .I0(__1568__),
    .O(__2742__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6905__ (
    .I1(RESET),
    .I0(__296__),
    .O(__2743__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6906__ (
    .I1(RESET),
    .I0(__1410__),
    .O(__2744__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6907__ (
    .I2(RESET),
    .I1(__1122__),
    .I0(__1116__),
    .O(__2745__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6908__ (
    .I1(RESET),
    .I0(__484__),
    .O(__2746__)
  );
  LUT5 #(
    .INIT(32'h14414114)
  ) __6909__ (
    .I4(__1597__),
    .I3(__1693__),
    .I2(__1629__),
    .I1(__1661__),
    .I0(TM0),
    .O(__2747__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6910__ (
    .I5(TM0),
    .I4(__1469__),
    .I3(__1437__),
    .I2(__1405__),
    .I1(__1501__),
    .I0(__1373__),
    .O(__2748__)
  );
  LUT6 #(
    .INIT(64'h00fff8f800000000)
  ) __6911__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__2748__),
    .I2(__2747__),
    .I1(TM0),
    .I0(__1506__),
    .O(__2749__)
  );
  LUT6 #(
    .INIT(64'h4bb4b44bb44b4bb4)
  ) __6912__ (
    .I5(__215__),
    .I4(__149__),
    .I3(__181__),
    .I2(__247__),
    .I1(TM0),
    .I0(__280__),
    .O(__2750__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6913__ (
    .I1(TM0),
    .I0(__758__),
    .O(__2751__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6914__ (
    .I1(TM0),
    .I0(__585__),
    .O(__2752__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6915__ (
    .I5(TM1),
    .I4(__617__),
    .I3(__681__),
    .I2(__649__),
    .I1(__713__),
    .I0(TM0),
    .O(__2753__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __6916__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__2753__),
    .I2(__2752__),
    .I1(__2318__),
    .I0(__2751__),
    .O(__2754__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6917__ (
    .I1(RESET),
    .I0(__48__),
    .O(__2755__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6918__ (
    .I1(RESET),
    .I0(__1389__),
    .O(__2756__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6919__ (
    .I1(RESET),
    .I0(__1592__),
    .O(__2757__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6920__ (
    .I1(RESET),
    .I0(__584__),
    .O(__2758__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6921__ (
    .I1(RESET),
    .I0(__493__),
    .O(__2759__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6922__ (
    .I1(RESET),
    .I0(__1644__),
    .O(__2760__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6923__ (
    .I1(RESET),
    .I0(__1017__),
    .O(__2761__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6924__ (
    .I1(TM0),
    .I0(__119__),
    .O(__2762__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6925__ (
    .I5(TM1),
    .I4(__17__),
    .I3(__11__),
    .I2(__78__),
    .I1(__327__),
    .I0(TM0),
    .O(__2763__)
  );
  LUT5 #(
    .INIT(32'h41141441)
  ) __6926__ (
    .I4(__291__),
    .I3(__242__),
    .I2(__210__),
    .I1(__176__),
    .I0(TM0),
    .O(__2764__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __6927__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__2764__),
    .I2(__2104__),
    .I1(__2763__),
    .I0(__2762__),
    .O(__2765__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6928__ (
    .I1(RESET),
    .I0(__398__),
    .O(__2766__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6929__ (
    .I2(RESET),
    .I1(__513__),
    .I0(__573__),
    .O(__2767__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6930__ (
    .I1(RESET),
    .I0(__407__),
    .O(__2768__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6931__ (
    .I1(RESET),
    .I0(__1072__),
    .O(__2769__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6932__ (
    .I5(TM0),
    .I4(__624__),
    .I3(__688__),
    .I2(__656__),
    .I1(__720__),
    .I0(__559__),
    .O(__2770__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6933__ (
    .I5(TM0),
    .I4(__464__),
    .I3(__432__),
    .I2(__496__),
    .I1(__528__),
    .I0(__400__),
    .O(__2771__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __6934__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__2771__),
    .I0(__2770__),
    .O(__2772__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6935__ (
    .I1(RESET),
    .I0(__1424__),
    .O(__2773__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6936__ (
    .I1(TM0),
    .I0(__1533__),
    .O(__2774__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6937__ (
    .I5(TM1),
    .I4(__1570__),
    .I3(__1602__),
    .I2(__1666__),
    .I1(__1634__),
    .I0(TM0),
    .O(__2775__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6938__ (
    .I1(TM0),
    .I0(__1346__),
    .O(__2776__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6939__ (
    .I5(TM1),
    .I4(__1378__),
    .I3(__1474__),
    .I2(__1442__),
    .I1(__1410__),
    .I0(TM0),
    .O(__2777__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __6940__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__2777__),
    .I2(__2776__),
    .I1(__2775__),
    .I0(__2774__),
    .O(__2778__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6941__ (
    .I1(RESET),
    .I0(__441__),
    .O(__2779__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6942__ (
    .I1(RESET),
    .I0(__1593__),
    .O(__2780__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6943__ (
    .I1(RESET),
    .I0(__482__),
    .O(__2781__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6944__ (
    .I1(RESET),
    .I0(__770__),
    .O(__2782__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6945__ (
    .I5(TM0),
    .I4(__1393__),
    .I3(__1457__),
    .I2(__1425__),
    .I1(__1489__),
    .I0(__1361__),
    .O(__2783__)
  );
  LUT6 #(
    .INIT(64'h00fff8f800000000)
  ) __6946__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__2783__),
    .I2(__2477__),
    .I1(TM0),
    .I0(__1518__),
    .O(__2784__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6947__ (
    .I1(RESET),
    .I0(__595__),
    .O(__2785__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6948__ (
    .I1(RESET),
    .I0(__963__),
    .O(__2786__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6949__ (
    .I1(RESET),
    .I0(__1440__),
    .O(__2787__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6950__ (
    .I1(RESET),
    .I0(__980__),
    .O(__2788__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6951__ (
    .I1(RESET),
    .I0(__40__),
    .O(__2789__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6952__ (
    .I1(RESET),
    .I0(__1157__),
    .O(__2790__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6953__ (
    .I1(RESET),
    .I0(__1577__),
    .O(__2791__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6954__ (
    .I1(RESET),
    .I0(__589__),
    .O(__2792__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6955__ (
    .I1(RESET),
    .I0(__184__),
    .O(__2793__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6956__ (
    .I2(RESET),
    .I1(__382__),
    .I0(__320__),
    .O(__2794__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6957__ (
    .I1(RESET),
    .I0(__262__),
    .O(__2795__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6958__ (
    .I1(RESET),
    .I0(__1632__),
    .O(__2796__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6959__ (
    .I1(RESET),
    .I0(__13__),
    .O(__2797__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6960__ (
    .I1(RESET),
    .I0(__1223__),
    .O(__2798__)
  );
  LUT4 #(
    .INIT(16'h6900)
  ) __6961__ (
    .I3(RESET),
    .I2(__1727__),
    .I1(__1684__),
    .I0(__1706__),
    .O(__2799__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6962__ (
    .I1(RESET),
    .I0(__1540__),
    .O(__2800__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6963__ (
    .I2(RESET),
    .I1(__1528__),
    .I0(__1478__),
    .O(__2801__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6964__ (
    .I2(RESET),
    .I1(__959__),
    .I0(__927__),
    .O(__2802__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6965__ (
    .I2(RESET),
    .I1(__164__),
    .I0(__157__),
    .O(__2803__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6966__ (
    .I1(RESET),
    .I0(__1641__),
    .O(__2804__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6967__ (
    .I2(RESET),
    .I1(__949__),
    .I0(__905__),
    .O(__2805__)
  );
  LUT5 #(
    .INIT(32'h14414114)
  ) __6968__ (
    .I4(__307__),
    .I3(__33__),
    .I2(__6__),
    .I1(__339__),
    .I0(TM0),
    .O(__2806__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6969__ (
    .I5(TM0),
    .I4(__135__),
    .I3(__233__),
    .I2(__267__),
    .I1(__102__),
    .I0(__298__),
    .O(__2807__)
  );
  LUT6 #(
    .INIT(64'h00fff8f800000000)
  ) __6970__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__2807__),
    .I2(__2806__),
    .I1(TM0),
    .I0(__159__),
    .O(__2808__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6971__ (
    .I1(TM0),
    .I0(__1530__),
    .O(__2809__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6972__ (
    .I1(TM0),
    .I0(__1349__),
    .O(__2810__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6973__ (
    .I5(TM1),
    .I4(__1413__),
    .I3(__1381__),
    .I2(__1445__),
    .I1(__1477__),
    .I0(TM0),
    .O(__2811__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __6974__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__2811__),
    .I2(__2810__),
    .I1(__2329__),
    .I0(__2809__),
    .O(__2812__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6975__ (
    .I1(RESET),
    .I0(__1379__),
    .O(__2813__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6976__ (
    .I5(TM0),
    .I4(__1429__),
    .I3(__1461__),
    .I2(__1493__),
    .I1(__1397__),
    .I0(__1322__),
    .O(__2814__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6977__ (
    .I5(TM0),
    .I4(__1237__),
    .I3(__1301__),
    .I2(__1269__),
    .I1(__1205__),
    .I0(__1173__),
    .O(__2815__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __6978__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__2815__),
    .I0(__2814__),
    .O(__2816__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __6979__ (
    .I2(RESET),
    .I1(__364__),
    .I0(__338__),
    .O(__2817__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6980__ (
    .I1(RESET),
    .I0(__1183__),
    .O(__2818__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6981__ (
    .I1(RESET),
    .I0(__226__),
    .O(__2819__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6982__ (
    .I1(RESET),
    .I0(__87__),
    .O(__2820__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6983__ (
    .I1(RESET),
    .I0(__1185__),
    .O(__2821__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6984__ (
    .I1(RESET),
    .I0(__995__),
    .O(__2822__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6985__ (
    .I1(RESET),
    .I0(__701__),
    .O(__2823__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6986__ (
    .I1(RESET),
    .I0(__416__),
    .O(__2824__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6987__ (
    .I1(RESET),
    .I0(__1555__),
    .O(__2825__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6988__ (
    .I1(RESET),
    .I0(__965__),
    .O(__2826__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6989__ (
    .I1(RESET),
    .I0(__237__),
    .O(__2827__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6990__ (
    .I1(RESET),
    .I0(__653__),
    .O(__2828__)
  );
  LUT5 #(
    .INIT(32'h14414114)
  ) __6991__ (
    .I4(__1659__),
    .I3(__1627__),
    .I2(__1595__),
    .I1(__1691__),
    .I0(TM0),
    .O(__2829__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __6992__ (
    .I5(TM0),
    .I4(__1467__),
    .I3(__1435__),
    .I2(__1403__),
    .I1(__1499__),
    .I0(__1371__),
    .O(__2830__)
  );
  LUT6 #(
    .INIT(64'h00fff8f800000000)
  ) __6993__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__2830__),
    .I2(__2829__),
    .I1(TM0),
    .I0(__1508__),
    .O(__2831__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6994__ (
    .I1(RESET),
    .I0(__1271__),
    .O(__2832__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6995__ (
    .I1(RESET),
    .I0(__1161__),
    .O(__2833__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6996__ (
    .I1(RESET),
    .I0(__1260__),
    .O(__2834__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6997__ (
    .I1(TM0),
    .I0(__1343__),
    .O(__2835__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __6998__ (
    .I5(TM1),
    .I4(__1376__),
    .I3(__1440__),
    .I2(__1408__),
    .I1(__1472__),
    .I0(TM0),
    .O(__2836__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __6999__ (
    .I1(TM0),
    .I0(__1152__),
    .O(__2837__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __7000__ (
    .I5(TM1),
    .I4(__1248__),
    .I3(__1216__),
    .I2(__1184__),
    .I1(__1280__),
    .I0(TM0),
    .O(__2838__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __7001__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__2838__),
    .I2(__2837__),
    .I1(__2836__),
    .I0(__2835__),
    .O(__2839__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7002__ (
    .I1(RESET),
    .I0(__1386__),
    .O(__2840__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7003__ (
    .I1(TM0),
    .I0(__1341__),
    .O(__2841__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7004__ (
    .I1(TM0),
    .I0(__1154__),
    .O(__2842__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __7005__ (
    .I5(TM1),
    .I4(__1282__),
    .I3(__1250__),
    .I2(__1218__),
    .I1(__1186__),
    .I0(TM0),
    .O(__2843__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __7006__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__2843__),
    .I2(__2842__),
    .I1(__2777__),
    .I0(__2841__),
    .O(__2844__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7007__ (
    .I1(RESET),
    .I0(__167__),
    .O(__2845__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7008__ (
    .I2(TM0),
    .I1(__1703__),
    .I0(DATA_0_7),
    .O(__2846__)
  );
  LUT5 #(
    .INIT(32'h14414114)
  ) __7009__ (
    .I4(__1656__),
    .I3(__1624__),
    .I2(__1592__),
    .I1(__1688__),
    .I0(TM0),
    .O(__2847__)
  );
  LUT6 #(
    .INIT(64'hff88f0f000000000)
  ) __7010__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__2847__),
    .I2(__2846__),
    .I1(TM0),
    .I0(__1560__),
    .O(__2848__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7011__ (
    .I2(RESET),
    .I1(__1525__),
    .I0(__1481__),
    .O(__2849__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7012__ (
    .I1(RESET),
    .I0(__206__),
    .O(__2850__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7013__ (
    .I1(RESET),
    .I0(__1261__),
    .O(__2851__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7014__ (
    .I2(RESET),
    .I1(__903__),
    .I0(__951__),
    .O(__2852__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7015__ (
    .I1(TM0),
    .I0(__765__),
    .O(__2853__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __7016__ (
    .I5(TM1),
    .I4(__898__),
    .I3(__866__),
    .I2(__834__),
    .I1(__802__),
    .I0(TM0),
    .O(__2854__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7017__ (
    .I1(TM0),
    .I0(__578__),
    .O(__2855__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __7018__ (
    .I5(TM1),
    .I4(__642__),
    .I3(__610__),
    .I2(__674__),
    .I1(__706__),
    .I0(TM0),
    .O(__2856__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __7019__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__2856__),
    .I2(__2855__),
    .I1(__2854__),
    .I0(__2853__),
    .O(__2857__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7020__ (
    .I1(RESET),
    .I0(__993__),
    .O(__2858__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7021__ (
    .I1(RESET),
    .I0(__109__),
    .O(__2859__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7022__ (
    .I2(TM0),
    .I1(__1706__),
    .I0(DATA_0_10),
    .O(__2860__)
  );
  LUT5 #(
    .INIT(32'h14414114)
  ) __7023__ (
    .I4(__1653__),
    .I3(__1621__),
    .I2(__1589__),
    .I1(__1685__),
    .I0(TM0),
    .O(__2861__)
  );
  LUT6 #(
    .INIT(64'hff88f0f000000000)
  ) __7024__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__2861__),
    .I2(__2860__),
    .I1(TM0),
    .I0(__1557__),
    .O(__2862__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7025__ (
    .I1(RESET),
    .I0(__185__),
    .O(__2863__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7026__ (
    .I1(RESET),
    .I0(__290__),
    .O(__2864__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7027__ (
    .I1(RESET),
    .I0(__430__),
    .O(__2865__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7028__ (
    .I1(RESET),
    .I0(__428__),
    .O(__2866__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7029__ (
    .I1(RESET),
    .I0(__410__),
    .O(__2867__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7030__ (
    .I1(RESET),
    .I0(__495__),
    .O(__2868__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7031__ (
    .I2(RESET),
    .I1(__1092__),
    .I0(__1146__),
    .O(__2869__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7032__ (
    .I1(RESET),
    .I0(__1066__),
    .O(__2870__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7033__ (
    .I1(RESET),
    .I0(__1601__),
    .O(__2871__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7034__ (
    .I1(RESET),
    .I0(__1561__),
    .O(__2872__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7035__ (
    .I1(RESET),
    .I0(__1369__),
    .O(__2873__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7036__ (
    .I1(RESET),
    .I0(__214__),
    .O(__2874__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7037__ (
    .I1(RESET),
    .I0(__1409__),
    .O(__2875__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7038__ (
    .I1(TM0),
    .I0(__1329__),
    .O(__2876__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7039__ (
    .I1(TM0),
    .I0(__1166__),
    .O(__2877__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __7040__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__2877__),
    .I2(__2669__),
    .I1(__2047__),
    .I0(__2876__),
    .O(__2878__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7041__ (
    .I1(RESET),
    .I0(__858__),
    .O(__2879__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7042__ (
    .I1(RESET),
    .I0(__474__),
    .O(__2880__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7043__ (
    .I1(RESET),
    .I0(__316__),
    .O(__2881__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7044__ (
    .I1(RESET),
    .I0(__1403__),
    .O(__2882__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7045__ (
    .I1(RESET),
    .I0(__700__),
    .O(__2883__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7046__ (
    .I1(RESET),
    .I0(__274__),
    .O(__2884__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7047__ (
    .I2(RESET),
    .I1(__750__),
    .I0(__720__),
    .O(__2885__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7048__ (
    .I1(RESET),
    .I0(__974__),
    .O(__2886__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7049__ (
    .I2(RESET),
    .I1(__545__),
    .I0(__541__),
    .O(__2887__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7050__ (
    .I1(RESET),
    .I0(__122__),
    .O(__2888__)
  );
  LUT5 #(
    .INIT(32'h14414114)
  ) __7051__ (
    .I4(__314__),
    .I3(__53__),
    .I2(__63__),
    .I1(__346__),
    .I0(TM0),
    .O(__2889__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7052__ (
    .I5(TM0),
    .I4(__180__),
    .I3(__214__),
    .I2(__246__),
    .I1(__148__),
    .I0(__279__),
    .O(__2890__)
  );
  LUT6 #(
    .INIT(64'h00fff8f800000000)
  ) __7053__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__2890__),
    .I2(__2889__),
    .I1(TM0),
    .I0(__156__),
    .O(__2891__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7054__ (
    .I1(RESET),
    .I0(__1645__),
    .O(__2892__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7055__ (
    .I2(TM0),
    .I1(__1725__),
    .I0(DATA_0_29),
    .O(__2893__)
  );
  LUT6 #(
    .INIT(64'hff88f0f000000000)
  ) __7056__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__2775__),
    .I2(__2893__),
    .I1(TM0),
    .I0(__1538__),
    .O(__2894__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7057__ (
    .I2(RESET),
    .I1(__1142__),
    .I0(__1096__),
    .O(__2895__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7058__ (
    .I1(RESET),
    .I0(__1211__),
    .O(__2896__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7059__ (
    .I1(TM0),
    .I0(__575__),
    .O(__2897__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7060__ (
    .I1(TM0),
    .I0(__384__),
    .O(__2898__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __7061__ (
    .I5(TM1),
    .I4(__448__),
    .I3(__512__),
    .I2(__480__),
    .I1(__416__),
    .I0(TM0),
    .O(__2899__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __7062__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__2899__),
    .I2(__2898__),
    .I1(__2069__),
    .I0(__2897__),
    .O(__2900__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7063__ (
    .I1(RESET),
    .I0(__1274__),
    .O(__2901__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7064__ (
    .I1(RESET),
    .I0(__269__),
    .O(__2902__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7065__ (
    .I1(RESET),
    .I0(__1616__),
    .O(__2903__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7066__ (
    .I2(RESET),
    .I1(__1303__),
    .I0(__1319__),
    .O(__2904__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7067__ (
    .I5(TM0),
    .I4(__637__),
    .I3(__733__),
    .I2(__701__),
    .I1(__669__),
    .I0(__546__),
    .O(__2905__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7068__ (
    .I5(TM0),
    .I4(__509__),
    .I3(__477__),
    .I2(__445__),
    .I1(__541__),
    .I0(__413__),
    .O(__2906__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __7069__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__2906__),
    .I0(__2905__),
    .O(__2907__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7070__ (
    .I1(RESET),
    .I0(__1576__),
    .O(__2908__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7071__ (
    .I1(RESET),
    .I0(__267__),
    .O(__2909__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7072__ (
    .I1(RESET),
    .I0(__634__),
    .O(__2910__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7073__ (
    .I1(RESET),
    .I0(__1580__),
    .O(__2911__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7074__ (
    .I1(RESET),
    .I0(__1558__),
    .O(__2912__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7075__ (
    .I1(RESET),
    .I0(__239__),
    .O(__2913__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7076__ (
    .I1(TM0),
    .I0(__70__),
    .O(__2914__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __7077__ (
    .I5(TM1),
    .I4(__16__),
    .I3(__35__),
    .I2(__88__),
    .I1(__331__),
    .I0(TM0),
    .O(__2915__)
  );
  LUT5 #(
    .INIT(32'h41141441)
  ) __7078__ (
    .I4(__192__),
    .I3(__174__),
    .I2(__207__),
    .I1(__188__),
    .I0(TM0),
    .O(__2916__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7079__ (
    .I1(TM0),
    .I0(__238__),
    .O(__2917__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __7080__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__2917__),
    .I2(__2916__),
    .I1(__2915__),
    .I0(__2914__),
    .O(__2918__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7081__ (
    .I2(RESET),
    .I1(__1093__),
    .I0(__1145__),
    .O(__2919__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7082__ (
    .I1(RESET),
    .I0(__1020__),
    .O(__2920__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7083__ (
    .I1(RESET),
    .I0(__89__),
    .O(__2921__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7084__ (
    .I1(TM0),
    .I0(__572__),
    .O(__2922__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7085__ (
    .I1(TM0),
    .I0(__387__),
    .O(__2923__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __7086__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__2923__),
    .I2(__2244__),
    .I1(__2402__),
    .I0(__2922__),
    .O(__2924__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7087__ (
    .I1(RESET),
    .I0(__683__),
    .O(__2925__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7088__ (
    .I1(RESET),
    .I0(__4__),
    .O(__2926__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7089__ (
    .I1(TM0),
    .I0(__573__),
    .O(__2927__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7090__ (
    .I1(TM0),
    .I0(__386__),
    .O(__2928__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __7091__ (
    .I5(TM1),
    .I4(__482__),
    .I3(__450__),
    .I2(__418__),
    .I1(__514__),
    .I0(TM0),
    .O(__2929__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __7092__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__2929__),
    .I2(__2928__),
    .I1(__2856__),
    .I0(__2927__),
    .O(__2930__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7093__ (
    .I1(RESET),
    .I0(__1572__),
    .O(__2931__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7094__ (
    .I1(RESET),
    .I0(__803__),
    .O(__2932__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7095__ (
    .I1(RESET),
    .I0(__173__),
    .O(__2933__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7096__ (
    .I1(RESET),
    .I0(__465__),
    .O(__2934__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7097__ (
    .I1(RESET),
    .I0(__221__),
    .O(__2935__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7098__ (
    .I5(TM0),
    .I4(__1465__),
    .I3(__1433__),
    .I2(__1401__),
    .I1(__1497__),
    .I0(__1369__),
    .O(__2936__)
  );
  LUT6 #(
    .INIT(64'h00fff8f800000000)
  ) __7099__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__2936__),
    .I2(__2610__),
    .I1(TM0),
    .I0(__1510__),
    .O(__2937__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7100__ (
    .I1(RESET),
    .I0(__879__),
    .O(__2938__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7101__ (
    .I1(RESET),
    .I0(__423__),
    .O(__2939__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7102__ (
    .I1(RESET),
    .I0(__232__),
    .O(__2940__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7103__ (
    .I1(RESET),
    .I0(__406__),
    .O(__2941__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7104__ (
    .I1(TM0),
    .I0(__944__),
    .O(__2942__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __7105__ (
    .I5(TM1),
    .I4(__1039__),
    .I3(__1007__),
    .I2(__1071__),
    .I1(__1103__),
    .I0(TM0),
    .O(__2943__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7106__ (
    .I1(TM0),
    .I0(__783__),
    .O(__2944__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __7107__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__2944__),
    .I2(__2505__),
    .I1(__2943__),
    .I0(__2942__),
    .O(__2945__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7108__ (
    .I1(RESET),
    .I0(__1253__),
    .O(__2946__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7109__ (
    .I1(RESET),
    .I0(__855__),
    .O(__2947__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7110__ (
    .I2(RESET),
    .I1(__115__),
    .I0(__176__),
    .O(__2948__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7111__ (
    .I1(TM0),
    .I0(__574__),
    .O(__2949__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __7112__ (
    .I5(TM1),
    .I4(__673__),
    .I3(__705__),
    .I2(__641__),
    .I1(__609__),
    .I0(TM0),
    .O(__2950__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7113__ (
    .I1(TM0),
    .I0(__385__),
    .O(__2951__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __7114__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__2951__),
    .I2(__2447__),
    .I1(__2950__),
    .I0(__2949__),
    .O(__2952__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7115__ (
    .I2(RESET),
    .I1(__381__),
    .I0(__321__),
    .O(__2953__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7116__ (
    .I1(RESET),
    .I0(__1455__),
    .O(__2954__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7117__ (
    .I1(RESET),
    .I0(__1266__),
    .O(__2955__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7118__ (
    .I1(RESET),
    .I0(__88__),
    .O(__2956__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7119__ (
    .I1(RESET),
    .I0(__792__),
    .O(__2957__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7120__ (
    .I1(RESET),
    .I0(__1242__),
    .O(__2958__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7121__ (
    .I1(RESET),
    .I0(__434__),
    .O(__2959__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7122__ (
    .I1(RESET),
    .I0(__1155__),
    .O(__2960__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7123__ (
    .I1(RESET),
    .I0(__0__),
    .O(__2961__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7124__ (
    .I5(TM0),
    .I4(__464__),
    .I3(__432__),
    .I2(__496__),
    .I1(__528__),
    .I0(__367__),
    .O(__2962__)
  );
  LUT6 #(
    .INIT(64'hff880f0f00000000)
  ) __7125__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__1790__),
    .I2(__2962__),
    .I1(TM0),
    .I0(__67__),
    .O(__2963__)
  );
  LUT4 #(
    .INIT(16'h6900)
  ) __7126__ (
    .I3(RESET),
    .I2(__131__),
    .I1(__143__),
    .I0(__101__),
    .O(__2964__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7127__ (
    .I1(RESET),
    .I0(__961__),
    .O(__2965__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7128__ (
    .I1(RESET),
    .I0(__1059__),
    .O(__2966__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7129__ (
    .I1(RESET),
    .I0(__790__),
    .O(__2967__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7130__ (
    .I5(TM0),
    .I4(__1079__),
    .I3(__1047__),
    .I2(__1015__),
    .I1(__1111__),
    .I0(__936__),
    .O(__2968__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7131__ (
    .I5(TM0),
    .I4(__823__),
    .I3(__887__),
    .I2(__855__),
    .I1(__919__),
    .I0(__791__),
    .O(__2969__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __7132__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__2969__),
    .I0(__2968__),
    .O(__2970__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7133__ (
    .I1(RESET),
    .I0(__1569__),
    .O(__2971__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7134__ (
    .I1(RESET),
    .I0(__1566__),
    .O(__2972__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7135__ (
    .I1(RESET),
    .I0(__1057__),
    .O(__2973__)
  );
  LUT4 #(
    .INIT(16'h6900)
  ) __7136__ (
    .I3(RESET),
    .I2(__162__),
    .I1(__131__),
    .I0(__152__),
    .O(__2974__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7137__ (
    .I2(TM0),
    .I1(__1724__),
    .I0(DATA_0_28),
    .O(__2975__)
  );
  LUT6 #(
    .INIT(64'hff88f0f000000000)
  ) __7138__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__2656__),
    .I2(__2975__),
    .I1(TM0),
    .I0(__1539__),
    .O(__2976__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7139__ (
    .I1(RESET),
    .I0(__1160__),
    .O(__2977__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7140__ (
    .I2(RESET),
    .I1(__727__),
    .I0(__743__),
    .O(__2978__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7141__ (
    .I1(RESET),
    .I0(__674__),
    .O(__2979__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7142__ (
    .I1(TM0),
    .I0(__1330__),
    .O(__2980__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __7143__ (
    .I5(TM1),
    .I4(__1453__),
    .I3(__1421__),
    .I2(__1389__),
    .I1(__1485__),
    .I0(TM0),
    .O(__2981__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7144__ (
    .I1(TM0),
    .I0(__1165__),
    .O(__2982__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __7145__ (
    .I5(TM1),
    .I4(__1261__),
    .I3(__1229__),
    .I2(__1197__),
    .I1(__1293__),
    .I0(TM0),
    .O(__2983__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __7146__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__2983__),
    .I2(__2982__),
    .I1(__2981__),
    .I0(__2980__),
    .O(__2984__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7147__ (
    .I5(TM0),
    .I4(__625__),
    .I3(__689__),
    .I2(__657__),
    .I1(__721__),
    .I0(__558__),
    .O(__2985__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7148__ (
    .I5(TM0),
    .I4(__497__),
    .I3(__433__),
    .I2(__465__),
    .I1(__529__),
    .I0(__401__),
    .O(__2986__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __7149__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__2986__),
    .I0(__2985__),
    .O(__2987__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7150__ (
    .I5(TM0),
    .I4(__1407__),
    .I3(__1503__),
    .I2(__1471__),
    .I1(__1439__),
    .I0(__1312__),
    .O(__2988__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7151__ (
    .I5(TM0),
    .I4(__1247__),
    .I3(__1215__),
    .I2(__1279__),
    .I1(__1311__),
    .I0(__1183__),
    .O(__2989__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __7152__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__2989__),
    .I0(__2988__),
    .O(__2990__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7153__ (
    .I1(RESET),
    .I0(__478__),
    .O(__2991__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7154__ (
    .I1(RESET),
    .I0(__1550__),
    .O(__2992__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7155__ (
    .I1(RESET),
    .I0(__399__),
    .O(__2993__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7156__ (
    .I1(RESET),
    .I0(__174__),
    .O(__2994__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7157__ (
    .I5(TM0),
    .I4(__1083__),
    .I3(__1051__),
    .I2(__1019__),
    .I1(__1115__),
    .I0(__932__),
    .O(__2995__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7158__ (
    .I5(TM0),
    .I4(__859__),
    .I3(__891__),
    .I2(__827__),
    .I1(__923__),
    .I0(__795__),
    .O(__2996__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __7159__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__2996__),
    .I0(__2995__),
    .O(__2997__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7160__ (
    .I2(RESET),
    .I1(__740__),
    .I0(__730__),
    .O(__2998__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7161__ (
    .I5(TM0),
    .I4(__1468__),
    .I3(__1436__),
    .I2(__1404__),
    .I1(__1500__),
    .I0(__1315__),
    .O(__2999__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7162__ (
    .I5(TM0),
    .I4(__1276__),
    .I3(__1308__),
    .I2(__1212__),
    .I1(__1244__),
    .I0(__1180__),
    .O(__3000__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __7163__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__3000__),
    .I0(__2999__),
    .O(__3001__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7164__ (
    .I1(RESET),
    .I0(__1049__),
    .O(__3002__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7165__ (
    .I1(RESET),
    .I0(__594__),
    .O(__3003__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __7166__ (
    .I1(RESET),
    .I0(__1152__),
    .O(__3004__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7167__ (
    .I5(TM0),
    .I4(__848__),
    .I3(__816__),
    .I2(__880__),
    .I1(__912__),
    .I0(__751__),
    .O(__3005__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7168__ (
    .I5(TM0),
    .I4(__624__),
    .I3(__688__),
    .I2(__656__),
    .I1(__720__),
    .I0(__592__),
    .O(__3006__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __7169__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__3006__),
    .I0(__3005__),
    .O(__3007__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7170__ (
    .I1(RESET),
    .I0(__272__),
    .O(__3008__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7171__ (
    .I1(RESET),
    .I0(__675__),
    .O(__3009__)
  );
  LUT4 #(
    .INIT(16'h6900)
  ) __7172__ (
    .I3(RESET),
    .I2(__1499__),
    .I1(__1507__),
    .I0(__1535__),
    .O(__3010__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7173__ (
    .I1(RESET),
    .I0(__422__),
    .O(__3011__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7174__ (
    .I5(TM0),
    .I4(__1270__),
    .I3(__1238__),
    .I2(__1302__),
    .I1(__1206__),
    .I0(__1129__),
    .O(__3012__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7175__ (
    .I5(TM0),
    .I4(__1110__),
    .I3(__1078__),
    .I2(__1046__),
    .I1(__1014__),
    .I0(__982__),
    .O(__3013__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __7176__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__3013__),
    .I0(__3012__),
    .O(__3014__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7177__ (
    .I5(TM0),
    .I4(__497__),
    .I3(__433__),
    .I2(__465__),
    .I1(__529__),
    .I0(__366__),
    .O(__3015__)
  );
  LUT5 #(
    .INIT(32'h14414114)
  ) __7178__ (
    .I4(__64__),
    .I3(__65__),
    .I2(__305__),
    .I1(__337__),
    .I0(TM0),
    .O(__3016__)
  );
  LUT6 #(
    .INIT(64'hff880f0f00000000)
  ) __7179__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__3016__),
    .I2(__3015__),
    .I1(TM0),
    .I0(__48__),
    .O(__3017__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7180__ (
    .I2(RESET),
    .I1(__1719__),
    .I0(__1671__),
    .O(__3018__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7181__ (
    .I2(RESET),
    .I1(__729__),
    .I0(__741__),
    .O(__3019__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7182__ (
    .I1(RESET),
    .I0(__91__),
    .O(__3020__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7183__ (
    .I1(RESET),
    .I0(__1029__),
    .O(__3021__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7184__ (
    .I2(TM0),
    .I1(__1713__),
    .I0(DATA_0_17),
    .O(__3022__)
  );
  LUT6 #(
    .INIT(64'hff88f0f000000000)
  ) __7185__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__2045__),
    .I2(__3022__),
    .I1(TM0),
    .I0(__1550__),
    .O(__3023__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7186__ (
    .I1(RESET),
    .I0(__1459__),
    .O(__3024__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7187__ (
    .I1(RESET),
    .I0(__54__),
    .O(__3025__)
  );
  LUT4 #(
    .INIT(16'h6900)
  ) __7188__ (
    .I3(RESET),
    .I2(__719__),
    .I1(__767__),
    .I0(__751__),
    .O(__3026__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7189__ (
    .I1(RESET),
    .I0(__1438__),
    .O(__3027__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7190__ (
    .I2(RESET),
    .I1(__376__),
    .I0(__326__),
    .O(__3028__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7191__ (
    .I1(RESET),
    .I0(__871__),
    .O(__3029__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7192__ (
    .I2(RESET),
    .I1(__1700__),
    .I0(__1690__),
    .O(__3030__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7193__ (
    .I1(RESET),
    .I0(__830__),
    .O(__3031__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7194__ (
    .I1(TM0),
    .I0(__1136__),
    .O(__3032__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7195__ (
    .I1(TM0),
    .I0(__975__),
    .O(__3033__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __7196__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__3033__),
    .I2(__2943__),
    .I1(__2146__),
    .I0(__3032__),
    .O(__3034__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __7197__ (
    .I1(RESET),
    .I0(__275__),
    .O(__3035__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7198__ (
    .I1(RESET),
    .I0(__1175__),
    .O(__3036__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7199__ (
    .I1(RESET),
    .I0(__1000__),
    .O(__3037__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7200__ (
    .I1(RESET),
    .I0(__796__),
    .O(__3038__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7201__ (
    .I1(RESET),
    .I0(__1626__),
    .O(__3039__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7202__ (
    .I1(TM0),
    .I0(__959__),
    .O(__3040__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __7203__ (
    .I5(TM1),
    .I4(__1056__),
    .I3(__1024__),
    .I2(__992__),
    .I1(__1088__),
    .I0(TM0),
    .O(__3041__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7204__ (
    .I1(TM0),
    .I0(__768__),
    .O(__3042__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __7205__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__3042__),
    .I2(__2067__),
    .I1(__3041__),
    .I0(__3040__),
    .O(__3043__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7206__ (
    .I1(RESET),
    .I0(__1560__),
    .O(__3044__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7207__ (
    .I1(RESET),
    .I0(__424__),
    .O(__3045__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7208__ (
    .I1(RESET),
    .I0(__832__),
    .O(__3046__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7209__ (
    .I1(RESET),
    .I0(__680__),
    .O(__3047__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7210__ (
    .I1(RESET),
    .I0(__1173__),
    .O(__3048__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7211__ (
    .I1(RESET),
    .I0(__1022__),
    .O(__3049__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7212__ (
    .I1(RESET),
    .I0(__1600__),
    .O(__3050__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7213__ (
    .I1(RESET),
    .I0(__1246__),
    .O(__3051__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7214__ (
    .I2(RESET),
    .I1(__906__),
    .I0(__948__),
    .O(__3052__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7215__ (
    .I1(RESET),
    .I0(__36__),
    .O(__3053__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7216__ (
    .I1(RESET),
    .I0(__181__),
    .O(__3054__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7217__ (
    .I2(TM0),
    .I1(__1705__),
    .I0(DATA_0_9),
    .O(__3055__)
  );
  LUT5 #(
    .INIT(32'h14414114)
  ) __7218__ (
    .I4(__1654__),
    .I3(__1686__),
    .I2(__1590__),
    .I1(__1622__),
    .I0(TM0),
    .O(__3056__)
  );
  LUT6 #(
    .INIT(64'hff88f0f000000000)
  ) __7219__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__3056__),
    .I2(__3055__),
    .I1(TM0),
    .I0(__1558__),
    .O(__3057__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7220__ (
    .I1(RESET),
    .I0(__1549__),
    .O(__3058__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7221__ (
    .I1(RESET),
    .I0(__1450__),
    .O(__3059__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7222__ (
    .I2(RESET),
    .I1(__1320__),
    .I0(__1302__),
    .O(__3060__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7223__ (
    .I1(RESET),
    .I0(__808__),
    .O(__3061__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7224__ (
    .I1(RESET),
    .I0(__846__),
    .O(__3062__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7225__ (
    .I1(RESET),
    .I0(__18__),
    .O(__3063__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7226__ (
    .I1(RESET),
    .I0(__1356__),
    .O(__3064__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7227__ (
    .I2(RESET),
    .I1(__1688__),
    .I0(__1702__),
    .O(__3065__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7228__ (
    .I1(RESET),
    .I0(__1210__),
    .O(__3066__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7229__ (
    .I1(RESET),
    .I0(__644__),
    .O(__3067__)
  );
  LUT6 #(
    .INIT(64'h4bb4b44bb44b4bb4)
  ) __7230__ (
    .I5(__258__),
    .I4(__197__),
    .I3(__224__),
    .I2(__163__),
    .I1(TM0),
    .I0(__289__),
    .O(__3068__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7231__ (
    .I2(RESET),
    .I1(__756__),
    .I0(__714__),
    .O(__3069__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7232__ (
    .I1(RESET),
    .I0(__387__),
    .O(__3070__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7233__ (
    .I1(RESET),
    .I0(__1657__),
    .O(__3071__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7234__ (
    .I2(RESET),
    .I1(__1133__),
    .I0(__1105__),
    .O(__3072__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7235__ (
    .I1(RESET),
    .I0(__816__),
    .O(__3073__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7236__ (
    .I2(RESET),
    .I1(__1285__),
    .I0(__1337__),
    .O(__3074__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7237__ (
    .I1(RESET),
    .I0(__508__),
    .O(__3075__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7238__ (
    .I1(RESET),
    .I0(__288__),
    .O(__3076__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7239__ (
    .I1(RESET),
    .I0(__388__),
    .O(__3077__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7240__ (
    .I1(RESET),
    .I0(__197__),
    .O(__3078__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7241__ (
    .I1(RESET),
    .I0(__777__),
    .O(__3079__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7242__ (
    .I1(TM0),
    .I0(__383__),
    .O(__3080__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7243__ (
    .I1(TM0),
    .I0(__112__),
    .O(__3081__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __7244__ (
    .I5(TM1),
    .I4(__51__),
    .I3(__61__),
    .I2(__80__),
    .I1(__320__),
    .I0(TM0),
    .O(__3082__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __7245__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__3082__),
    .I2(__3081__),
    .I1(__2899__),
    .I0(__3080__),
    .O(__3083__)
  );
  LUT4 #(
    .INIT(16'h6900)
  ) __7246__ (
    .I3(RESET),
    .I2(__731__),
    .I1(__767__),
    .I0(__739__),
    .O(__3084__)
  );
  LUT5 #(
    .INIT(32'h14414114)
  ) __7247__ (
    .I4(__1695__),
    .I3(__1599__),
    .I2(__1663__),
    .I1(__1631__),
    .I0(TM0),
    .O(__3085__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7248__ (
    .I5(TM0),
    .I4(__1407__),
    .I3(__1503__),
    .I2(__1471__),
    .I1(__1439__),
    .I0(__1375__),
    .O(__3086__)
  );
  LUT6 #(
    .INIT(64'h00fff8f800000000)
  ) __7249__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__3086__),
    .I2(__3085__),
    .I1(TM0),
    .I0(__1504__),
    .O(__3087__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7250__ (
    .I2(RESET),
    .I1(__1724__),
    .I0(__1666__),
    .O(__3088__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7251__ (
    .I1(RESET),
    .I0(__1056__),
    .O(__3089__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7252__ (
    .I1(RESET),
    .I0(__1035__),
    .O(__3090__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7253__ (
    .I5(TM0),
    .I4(__859__),
    .I3(__891__),
    .I2(__827__),
    .I1(__923__),
    .I0(__740__),
    .O(__3091__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7254__ (
    .I5(TM0),
    .I4(__635__),
    .I3(__699__),
    .I2(__667__),
    .I1(__731__),
    .I0(__603__),
    .O(__3092__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __7255__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__3092__),
    .I0(__3091__),
    .O(__3093__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7256__ (
    .I1(TM0),
    .I0(__756__),
    .O(__3094__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7257__ (
    .I1(TM0),
    .I0(__587__),
    .O(__3095__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __7258__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__3095__),
    .I2(__2714__),
    .I1(__2681__),
    .I0(__3094__),
    .O(__3096__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7259__ (
    .I1(RESET),
    .I0(__831__),
    .O(__3097__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7260__ (
    .I1(RESET),
    .I0(__305__),
    .O(__3098__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7261__ (
    .I1(RESET),
    .I0(__419__),
    .O(__3099__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7262__ (
    .I1(RESET),
    .I0(__33__),
    .O(__3100__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7263__ (
    .I1(TM0),
    .I0(__368__),
    .O(__3101__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __7264__ (
    .I5(TM1),
    .I4(__463__),
    .I3(__527__),
    .I2(__495__),
    .I1(__431__),
    .I0(TM0),
    .O(__3102__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7265__ (
    .I1(TM0),
    .I0(__120__),
    .O(__3103__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __7266__ (
    .I5(TM1),
    .I4(__92__),
    .I3(__56__),
    .I2(__335__),
    .I1(__303__),
    .I0(TM0),
    .O(__3104__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __7267__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__3104__),
    .I2(__3103__),
    .I1(__3102__),
    .I0(__3101__),
    .O(__3105__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7268__ (
    .I1(RESET),
    .I0(__1466__),
    .O(__3106__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7269__ (
    .I1(RESET),
    .I0(__1350__),
    .O(__3107__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7270__ (
    .I1(RESET),
    .I0(__660__),
    .O(__3108__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7271__ (
    .I1(RESET),
    .I0(__1436__),
    .O(__3109__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7272__ (
    .I2(RESET),
    .I1(__1705__),
    .I0(__1685__),
    .O(__3110__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7273__ (
    .I5(TM0),
    .I4(__1398__),
    .I3(__1494__),
    .I2(__1462__),
    .I1(__1430__),
    .I0(__1366__),
    .O(__3111__)
  );
  LUT6 #(
    .INIT(64'h00fff8f800000000)
  ) __7274__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__3111__),
    .I2(__3056__),
    .I1(TM0),
    .I0(__1513__),
    .O(__3112__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7275__ (
    .I5(TM0),
    .I4(__1469__),
    .I3(__1437__),
    .I2(__1405__),
    .I1(__1501__),
    .I0(__1314__),
    .O(__3113__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7276__ (
    .I5(TM0),
    .I4(__1245__),
    .I3(__1277__),
    .I2(__1213__),
    .I1(__1309__),
    .I0(__1181__),
    .O(__3114__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __7277__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__3114__),
    .I0(__3113__),
    .O(__3115__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7278__ (
    .I5(TM0),
    .I4(__1247__),
    .I3(__1215__),
    .I2(__1279__),
    .I1(__1311__),
    .I0(__1120__),
    .O(__3116__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7279__ (
    .I5(TM0),
    .I4(__1055__),
    .I3(__1023__),
    .I2(__1087__),
    .I1(__1119__),
    .I0(__991__),
    .O(__3117__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __7280__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__3117__),
    .I0(__3116__),
    .O(__3118__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7281__ (
    .I1(RESET),
    .I0(__1442__),
    .O(__3119__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7282__ (
    .I1(RESET),
    .I0(__843__),
    .O(__3120__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7283__ (
    .I2(RESET),
    .I1(__570__),
    .I0(__516__),
    .O(__3121__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7284__ (
    .I2(RESET),
    .I1(__1296__),
    .I0(__1326__),
    .O(__3122__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7285__ (
    .I1(RESET),
    .I0(__224__),
    .O(__3123__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7286__ (
    .I1(RESET),
    .I0(__1457__),
    .O(__3124__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7287__ (
    .I1(RESET),
    .I0(__1265__),
    .O(__3125__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7288__ (
    .I2(RESET),
    .I1(__153__),
    .I0(__161__),
    .O(__3126__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7289__ (
    .I1(RESET),
    .I0(__1364__),
    .O(__3127__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7290__ (
    .I1(RESET),
    .I0(__859__),
    .O(__3128__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7291__ (
    .I5(TM0),
    .I4(__509__),
    .I3(__477__),
    .I2(__445__),
    .I1(__541__),
    .I0(__354__),
    .O(__3129__)
  );
  LUT6 #(
    .INIT(64'hff880f0f00000000)
  ) __7292__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__2073__),
    .I2(__3129__),
    .I1(TM0),
    .I0(__81__),
    .O(__3130__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7293__ (
    .I1(RESET),
    .I0(__1021__),
    .O(__3131__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7294__ (
    .I1(RESET),
    .I0(__121__),
    .O(__3132__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7295__ (
    .I1(TM0),
    .I0(__1142__),
    .O(__3133__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7296__ (
    .I1(TM0),
    .I0(__969__),
    .O(__3134__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __7297__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__3134__),
    .I2(__2316__),
    .I1(__2123__),
    .I0(__3133__),
    .O(__3135__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __7298__ (
    .I1(RESET),
    .I0(__960__),
    .O(__3136__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7299__ (
    .I2(RESET),
    .I1(__1316__),
    .I0(__1306__),
    .O(__3137__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7300__ (
    .I1(RESET),
    .I0(__1215__),
    .O(__3138__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7301__ (
    .I2(RESET),
    .I1(__1313__),
    .I0(__1309__),
    .O(__3139__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7302__ (
    .I1(RESET),
    .I0(__1556__),
    .O(__3140__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7303__ (
    .I1(RESET),
    .I0(__480__),
    .O(__3141__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7304__ (
    .I1(RESET),
    .I0(__881__),
    .O(__3142__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7305__ (
    .I1(RESET),
    .I0(__1153__),
    .O(__3143__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7306__ (
    .I1(RESET),
    .I0(__1030__),
    .O(__3144__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7307__ (
    .I1(RESET),
    .I0(__219__),
    .O(__3145__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7308__ (
    .I5(TM0),
    .I4(__1460__),
    .I3(__1428__),
    .I2(__1396__),
    .I1(__1492__),
    .I0(__1323__),
    .O(__3146__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7309__ (
    .I5(TM0),
    .I4(__1236__),
    .I3(__1268__),
    .I2(__1204__),
    .I1(__1300__),
    .I0(__1172__),
    .O(__3147__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __7310__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__3147__),
    .I0(__3146__),
    .O(__3148__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7311__ (
    .I1(RESET),
    .I0(__1590__),
    .O(__3149__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7312__ (
    .I1(RESET),
    .I0(__1542__),
    .O(__3150__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7313__ (
    .I1(RESET),
    .I0(__1399__),
    .O(__3151__)
  );
  LUT5 #(
    .INIT(32'h14414114)
  ) __7314__ (
    .I4(__1587__),
    .I3(__1651__),
    .I2(__1619__),
    .I1(__1683__),
    .I0(TM0),
    .O(__3152__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7315__ (
    .I5(TM0),
    .I4(__1395__),
    .I3(__1459__),
    .I2(__1427__),
    .I1(__1491__),
    .I0(__1363__),
    .O(__3153__)
  );
  LUT6 #(
    .INIT(64'h00fff8f800000000)
  ) __7316__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__3153__),
    .I2(__3152__),
    .I1(TM0),
    .I0(__1516__),
    .O(__3154__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7317__ (
    .I1(RESET),
    .I0(__1557__),
    .O(__3155__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7318__ (
    .I1(RESET),
    .I0(__1170__),
    .O(__3156__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7319__ (
    .I1(TM0),
    .I0(__1524__),
    .O(__3157__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7320__ (
    .I1(TM0),
    .I0(__1355__),
    .O(__3158__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __7321__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__3158__),
    .I2(__2312__),
    .I1(__1960__),
    .I0(__3157__),
    .O(__3159__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7322__ (
    .I5(TM0),
    .I4(__693__),
    .I3(__629__),
    .I2(__725__),
    .I1(__661__),
    .I0(__554__),
    .O(__3160__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7323__ (
    .I5(TM0),
    .I4(__533__),
    .I3(__469__),
    .I2(__501__),
    .I1(__437__),
    .I0(__405__),
    .O(__3161__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __7324__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__3161__),
    .I0(__3160__),
    .O(__3162__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7325__ (
    .I2(RESET),
    .I1(__1325__),
    .I0(__1297__),
    .O(__3163__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7326__ (
    .I1(RESET),
    .I0(__1579__),
    .O(__3164__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7327__ (
    .I1(RESET),
    .I0(__819__),
    .O(__3165__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7328__ (
    .I1(RESET),
    .I0(__669__),
    .O(__3166__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7329__ (
    .I1(RESET),
    .I0(__1605__),
    .O(__3167__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7330__ (
    .I1(RESET),
    .I0(__1086__),
    .O(__3168__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7331__ (
    .I2(RESET),
    .I1(__150__),
    .I0(__147__),
    .O(__3169__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7332__ (
    .I1(RESET),
    .I0(__233__),
    .O(__3170__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7333__ (
    .I2(RESET),
    .I1(__745__),
    .I0(__725__),
    .O(__3171__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7334__ (
    .I1(RESET),
    .I0(__629__),
    .O(__3172__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7335__ (
    .I1(RESET),
    .I0(__1196__),
    .O(__3173__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7336__ (
    .I1(RESET),
    .I0(__689__),
    .O(__3174__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7337__ (
    .I5(TM0),
    .I4(__1076__),
    .I3(__1044__),
    .I2(__1012__),
    .I1(__1108__),
    .I0(__939__),
    .O(__3175__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7338__ (
    .I5(TM0),
    .I4(__884__),
    .I3(__852__),
    .I2(__820__),
    .I1(__916__),
    .I0(__788__),
    .O(__3176__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __7339__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__3176__),
    .I0(__3175__),
    .O(__3177__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7340__ (
    .I1(RESET),
    .I0(__1650__),
    .O(__3178__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7341__ (
    .I1(TM0),
    .I0(__1335__),
    .O(__3179__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __7342__ (
    .I5(TM1),
    .I4(__1480__),
    .I3(__1384__),
    .I2(__1448__),
    .I1(__1416__),
    .I0(TM0),
    .O(__3180__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7343__ (
    .I1(TM0),
    .I0(__1160__),
    .O(__3181__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __7344__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__3181__),
    .I2(__2371__),
    .I1(__3180__),
    .I0(__3179__),
    .O(__3182__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7345__ (
    .I1(RESET),
    .I0(__409__),
    .O(__3183__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7346__ (
    .I1(RESET),
    .I0(__1174__),
    .O(__3184__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7347__ (
    .I2(RESET),
    .I1(__552__),
    .I0(__534__),
    .O(__3185__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7348__ (
    .I2(RESET),
    .I1(__945__),
    .I0(__909__),
    .O(__3186__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7349__ (
    .I2(TM0),
    .I1(__1718__),
    .I0(DATA_0_22),
    .O(__3187__)
  );
  LUT6 #(
    .INIT(64'hff88f0f000000000)
  ) __7350__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__1984__),
    .I2(__3187__),
    .I1(TM0),
    .I0(__1545__),
    .O(__3188__)
  );
  LUT4 #(
    .INIT(16'h6900)
  ) __7351__ (
    .I3(RESET),
    .I2(__724__),
    .I1(__767__),
    .I0(__746__),
    .O(__3189__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7352__ (
    .I1(TM0),
    .I0(__565__),
    .O(__3190__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7353__ (
    .I1(TM0),
    .I0(__394__),
    .O(__3191__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __7354__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__3191__),
    .I2(__2164__),
    .I1(__1868__),
    .I0(__3190__),
    .O(__3192__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7355__ (
    .I5(TM0),
    .I4(__505__),
    .I3(__473__),
    .I2(__441__),
    .I1(__537__),
    .I0(__358__),
    .O(__3193__)
  );
  LUT5 #(
    .INIT(32'h14414114)
  ) __7356__ (
    .I4(__31__),
    .I3(__345__),
    .I2(__313__),
    .I1(__0__),
    .I0(TM0),
    .O(__3194__)
  );
  LUT6 #(
    .INIT(64'hff880f0f00000000)
  ) __7357__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__3194__),
    .I2(__3193__),
    .I1(TM0),
    .I0(__99__),
    .O(__3195__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7358__ (
    .I1(RESET),
    .I0(__1367__),
    .O(__3196__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7359__ (
    .I1(RESET),
    .I0(__238__),
    .O(__3197__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7360__ (
    .I1(RESET),
    .I0(__1349__),
    .O(__3198__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7361__ (
    .I2(RESET),
    .I1(__1704__),
    .I0(__1686__),
    .O(__3199__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7362__ (
    .I1(RESET),
    .I0(__2__),
    .O(__3200__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7363__ (
    .I1(RESET),
    .I0(__304__),
    .O(__3201__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7364__ (
    .I1(TM0),
    .I0(__74__),
    .O(__3202__)
  );
  LUT5 #(
    .INIT(32'h41141441)
  ) __7365__ (
    .I4(__139__),
    .I3(__170__),
    .I2(__203__),
    .I1(__106__),
    .I0(TM0),
    .O(__3203__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7366__ (
    .I1(TM0),
    .I0(__234__),
    .O(__3204__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __7367__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__3204__),
    .I2(__3203__),
    .I1(__3104__),
    .I0(__3202__),
    .O(__3205__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7368__ (
    .I1(RESET),
    .I0(__1034__),
    .O(__3206__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7369__ (
    .I1(RESET),
    .I0(__1662__),
    .O(__3207__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7370__ (
    .I5(TM0),
    .I4(__668__),
    .I3(__732__),
    .I2(__700__),
    .I1(__636__),
    .I0(__547__),
    .O(__3208__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7371__ (
    .I5(TM0),
    .I4(__476__),
    .I3(__508__),
    .I2(__444__),
    .I1(__540__),
    .I0(__412__),
    .O(__3209__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __7372__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__3209__),
    .I0(__3208__),
    .O(__3210__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7373__ (
    .I1(RESET),
    .I0(__1159__),
    .O(__3211__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7374__ (
    .I1(RESET),
    .I0(__78__),
    .O(__3212__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7375__ (
    .I1(RESET),
    .I0(__220__),
    .O(__3213__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7376__ (
    .I2(RESET),
    .I1(__119__),
    .I0(__194__),
    .O(__3214__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7377__ (
    .I1(RESET),
    .I0(__51__),
    .O(__3215__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7378__ (
    .I1(RESET),
    .I0(__1573__),
    .O(__3216__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7379__ (
    .I1(RESET),
    .I0(__851__),
    .O(__3217__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7380__ (
    .I1(RESET),
    .I0(__234__),
    .O(__3218__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7381__ (
    .I1(RESET),
    .I0(__1582__),
    .O(__3219__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7382__ (
    .I1(RESET),
    .I0(__1080__),
    .O(__3220__)
  );
  LUT6 #(
    .INIT(64'h4bb4b44bb44b4bb4)
  ) __7383__ (
    .I5(__168__),
    .I4(__249__),
    .I3(__137__),
    .I2(__104__),
    .I1(TM0),
    .I0(__282__),
    .O(__3221__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7384__ (
    .I1(RESET),
    .I0(__1053__),
    .O(__3222__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7385__ (
    .I1(RESET),
    .I0(__848__),
    .O(__3223__)
  );
  LUT6 #(
    .INIT(64'h4bb4b44bb44b4bb4)
  ) __7386__ (
    .I5(__135__),
    .I4(__233__),
    .I3(__267__),
    .I2(__102__),
    .I1(TM0),
    .I0(__298__),
    .O(__3224__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7387__ (
    .I2(RESET),
    .I1(__1112__),
    .I0(__1126__),
    .O(__3225__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7388__ (
    .I1(RESET),
    .I0(__1247__),
    .O(__3226__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7389__ (
    .I1(RESET),
    .I0(__866__),
    .O(__3227__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7390__ (
    .I1(RESET),
    .I0(__1347__),
    .O(__3228__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7391__ (
    .I2(TM0),
    .I1(__1696__),
    .I0(DATA_0_0),
    .O(__3229__)
  );
  LUT6 #(
    .INIT(64'hff88f0f000000000)
  ) __7392__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__3085__),
    .I2(__3229__),
    .I1(TM0),
    .I0(__1567__),
    .O(__3230__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7393__ (
    .I1(RESET),
    .I0(__1051__),
    .O(__3231__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7394__ (
    .I1(RESET),
    .I0(__989__),
    .O(__3232__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7395__ (
    .I1(RESET),
    .I0(__1468__),
    .O(__3233__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7396__ (
    .I1(RESET),
    .I0(__1656__),
    .O(__3234__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7397__ (
    .I1(RESET),
    .I0(__598__),
    .O(__3235__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7398__ (
    .I1(TM0),
    .I0(__275__),
    .O(__3236__)
  );
  LUT6 #(
    .INIT(64'h6996966996696996)
  ) __7399__ (
    .I5(TM1),
    .I4(__229__),
    .I3(__262__),
    .I2(__294__),
    .I1(__196__),
    .I0(__3236__),
    .O(__3237__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7400__ (
    .I2(RESET),
    .I1(__378__),
    .I0(__324__),
    .O(__3238__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7401__ (
    .I1(RESET),
    .I0(__838__),
    .O(__3239__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7402__ (
    .I2(RESET),
    .I1(__1527__),
    .I0(__1479__),
    .O(__3240__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7403__ (
    .I1(RESET),
    .I0(__1077__),
    .O(__3241__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7404__ (
    .I1(RESET),
    .I0(__869__),
    .O(__3242__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7405__ (
    .I1(RESET),
    .I0(__253__),
    .O(__3243__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7406__ (
    .I1(TM0),
    .I0(__1527__),
    .O(__3244__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7407__ (
    .I1(TM0),
    .I0(__1352__),
    .O(__3245__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __7408__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__3245__),
    .I2(__3180__),
    .I1(__2286__),
    .I0(__3244__),
    .O(__3246__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7409__ (
    .I1(RESET),
    .I0(__1585__),
    .O(__3247__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7410__ (
    .I5(TM0),
    .I4(__1240__),
    .I3(__1208__),
    .I2(__1304__),
    .I1(__1272__),
    .I0(__1127__),
    .O(__3248__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7411__ (
    .I5(TM0),
    .I4(__1080__),
    .I3(__1048__),
    .I2(__1016__),
    .I1(__1112__),
    .I0(__984__),
    .O(__3249__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __7412__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__3249__),
    .I0(__3248__),
    .O(__3250__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7413__ (
    .I1(RESET),
    .I0(__38__),
    .O(__3251__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7414__ (
    .I2(RESET),
    .I1(__1717__),
    .I0(__1673__),
    .O(__3252__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7415__ (
    .I1(RESET),
    .I0(__454__),
    .O(__3253__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7416__ (
    .I1(TM0),
    .I0(__958__),
    .O(__3254__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7417__ (
    .I1(TM0),
    .I0(__769__),
    .O(__3255__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __7418__ (
    .I5(TM1),
    .I4(__897__),
    .I3(__865__),
    .I2(__801__),
    .I1(__833__),
    .I0(TM0),
    .O(__3256__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __7419__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__3256__),
    .I2(__3255__),
    .I1(__2272__),
    .I0(__3254__),
    .O(__3257__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7420__ (
    .I2(RESET),
    .I1(__1318__),
    .I0(__1304__),
    .O(__3258__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7421__ (
    .I1(RESET),
    .I0(__1660__),
    .O(__3259__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7422__ (
    .I1(RESET),
    .I0(__433__),
    .O(__3260__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7423__ (
    .I5(TM0),
    .I4(__200__),
    .I3(__232__),
    .I2(__266__),
    .I1(__166__),
    .I0(__297__),
    .O(__3261__)
  );
  LUT6 #(
    .INIT(64'h00fff8f800000000)
  ) __7424__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__3261__),
    .I2(__2160__),
    .I1(TM0),
    .I0(__160__),
    .O(__3262__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7425__ (
    .I5(TM0),
    .I4(__1429__),
    .I3(__1461__),
    .I2(__1493__),
    .I1(__1397__),
    .I0(__1365__),
    .O(__3263__)
  );
  LUT6 #(
    .INIT(64'h00fff8f800000000)
  ) __7426__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__3263__),
    .I2(__2861__),
    .I1(TM0),
    .I0(__1514__),
    .O(__3264__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7427__ (
    .I1(RESET),
    .I0(__393__),
    .O(__3265__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7428__ (
    .I1(TM0),
    .I0(__114__),
    .O(__3266__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __7429__ (
    .I5(TM1),
    .I4(__27__),
    .I3(__37__),
    .I2(__90__),
    .I1(__325__),
    .I0(TM0),
    .O(__3267__)
  );
  LUT5 #(
    .INIT(32'h41141441)
  ) __7430__ (
    .I4(__222__),
    .I3(__256__),
    .I2(__287__),
    .I1(__190__),
    .I0(TM0),
    .O(__3268__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7431__ (
    .I1(TM0),
    .I0(__270__),
    .O(__3269__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __7432__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__3269__),
    .I2(__3268__),
    .I1(__3267__),
    .I0(__3266__),
    .O(__3270__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7433__ (
    .I1(RESET),
    .I0(__128__),
    .O(__3271__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7434__ (
    .I1(RESET),
    .I0(__805__),
    .O(__3272__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7435__ (
    .I1(RESET),
    .I0(__250__),
    .O(__3273__)
  );
  LUT4 #(
    .INIT(16'h6900)
  ) __7436__ (
    .I3(RESET),
    .I2(__916__),
    .I1(__959__),
    .I0(__938__),
    .O(__3274__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7437__ (
    .I1(RESET),
    .I0(__1087__),
    .O(__3275__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7438__ (
    .I1(TM0),
    .I0(__379__),
    .O(__3276__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7439__ (
    .I1(TM0),
    .I0(__111__),
    .O(__3277__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __7440__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__3277__),
    .I2(__2638__),
    .I1(__2487__),
    .I0(__3276__),
    .O(__3278__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7441__ (
    .I1(RESET),
    .I0(__663__),
    .O(__3279__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7442__ (
    .I1(RESET),
    .I0(__1184__),
    .O(__3280__)
  );
  LUT4 #(
    .INIT(16'h6900)
  ) __7443__ (
    .I3(RESET),
    .I2(__1151__),
    .I1(__1130__),
    .I0(__1108__),
    .O(__3281__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7444__ (
    .I1(RESET),
    .I0(__988__),
    .O(__3282__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7445__ (
    .I1(RESET),
    .I0(__1584__),
    .O(__3283__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7446__ (
    .I1(RESET),
    .I0(__667__),
    .O(__3284__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7447__ (
    .I1(RESET),
    .I0(__86__),
    .O(__3285__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7448__ (
    .I2(RESET),
    .I1(__331__),
    .I0(__371__),
    .O(__3286__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7449__ (
    .I2(RESET),
    .I1(__760__),
    .I0(__710__),
    .O(__3287__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7450__ (
    .I2(RESET),
    .I1(__566__),
    .I0(__520__),
    .O(__3288__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7451__ (
    .I1(RESET),
    .I0(__1640__),
    .O(__3289__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7452__ (
    .I1(RESET),
    .I0(__1412__),
    .O(__3290__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7453__ (
    .I1(RESET),
    .I0(__417__),
    .O(__3291__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7454__ (
    .I1(RESET),
    .I0(__837__),
    .O(__3292__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7455__ (
    .I1(RESET),
    .I0(__473__),
    .O(__3293__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7456__ (
    .I1(RESET),
    .I0(__302__),
    .O(__3294__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7457__ (
    .I2(RESET),
    .I1(__332__),
    .I0(__370__),
    .O(__3295__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7458__ (
    .I1(RESET),
    .I0(__432__),
    .O(__3296__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7459__ (
    .I1(RESET),
    .I0(__877__),
    .O(__3297__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7460__ (
    .I2(RESET),
    .I1(__1151__),
    .I0(__1119__),
    .O(__3298__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7461__ (
    .I1(RESET),
    .I0(__1464__),
    .O(__3299__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7462__ (
    .I2(RESET),
    .I1(__575__),
    .I0(__543__),
    .O(__3300__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7463__ (
    .I5(TM0),
    .I4(__136__),
    .I3(__103__),
    .I2(__167__),
    .I1(__253__),
    .I0(__286__),
    .O(__3301__)
  );
  LUT6 #(
    .INIT(64'h00fff8f800000000)
  ) __7464__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__3301__),
    .I2(__2300__),
    .I1(TM0),
    .I0(__158__),
    .O(__3302__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7465__ (
    .I1(RESET),
    .I0(__509__),
    .O(__3303__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7466__ (
    .I1(TM0),
    .I0(__1535__),
    .O(__3304__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __7467__ (
    .I5(TM1),
    .I4(__1632__),
    .I3(__1600__),
    .I2(__1568__),
    .I1(__1664__),
    .I0(TM0),
    .O(__3305__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7468__ (
    .I1(TM0),
    .I0(__1344__),
    .O(__3306__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __7469__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__3306__),
    .I2(__2836__),
    .I1(__3305__),
    .I0(__3304__),
    .O(__3307__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7470__ (
    .I2(TM0),
    .I1(__1698__),
    .I0(DATA_0_2),
    .O(__3308__)
  );
  LUT6 #(
    .INIT(64'hff88f0f000000000)
  ) __7471__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__2747__),
    .I2(__3308__),
    .I1(TM0),
    .I0(__1565__),
    .O(__3309__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7472__ (
    .I2(TM0),
    .I1(__1714__),
    .I0(DATA_0_18),
    .O(__3310__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __7473__ (
    .I5(TM1),
    .I4(__1645__),
    .I3(__1613__),
    .I2(__1581__),
    .I1(__1677__),
    .I0(TM0),
    .O(__3311__)
  );
  LUT6 #(
    .INIT(64'hff88f0f000000000)
  ) __7474__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__3311__),
    .I2(__3310__),
    .I1(TM0),
    .I0(__1549__),
    .O(__3312__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7475__ (
    .I1(RESET),
    .I0(__1229__),
    .O(__3313__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7476__ (
    .I5(TM0),
    .I4(__1470__),
    .I3(__1438__),
    .I2(__1406__),
    .I1(__1502__),
    .I0(__1313__),
    .O(__3314__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7477__ (
    .I5(TM0),
    .I4(__1278__),
    .I3(__1246__),
    .I2(__1214__),
    .I1(__1310__),
    .I0(__1182__),
    .O(__3315__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __7478__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__3315__),
    .I0(__3314__),
    .O(__3316__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7479__ (
    .I1(RESET),
    .I0(__888__),
    .O(__3317__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7480__ (
    .I1(RESET),
    .I0(__1192__),
    .O(__3318__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7481__ (
    .I1(RESET),
    .I0(__647__),
    .O(__3319__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7482__ (
    .I1(RESET),
    .I0(__874__),
    .O(__3320__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7483__ (
    .I2(RESET),
    .I1(__353__),
    .I0(__349__),
    .O(__3321__)
  );
  LUT6 #(
    .INIT(64'h4bb4b44bb44b4bb4)
  ) __7484__ (
    .I5(__179__),
    .I4(__213__),
    .I3(__263__),
    .I2(__147__),
    .I1(TM0),
    .I0(__295__),
    .O(__3322__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7485__ (
    .I1(RESET),
    .I0(__614__),
    .O(__3323__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7486__ (
    .I1(RESET),
    .I0(__1189__),
    .O(__3324__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7487__ (
    .I1(RESET),
    .I0(__451__),
    .O(__3325__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7488__ (
    .I1(RESET),
    .I0(__1263__),
    .O(__3326__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7489__ (
    .I1(RESET),
    .I0(__671__),
    .O(__3327__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7490__ (
    .I1(RESET),
    .I0(__85__),
    .O(__3328__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7491__ (
    .I1(RESET),
    .I0(__632__),
    .O(__3329__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7492__ (
    .I1(RESET),
    .I0(__294__),
    .O(__3330__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7493__ (
    .I1(RESET),
    .I0(__1391__),
    .O(__3331__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7494__ (
    .I1(RESET),
    .I0(__1048__),
    .O(__3332__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7495__ (
    .I1(RESET),
    .I0(__3__),
    .O(__3333__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7496__ (
    .I2(RESET),
    .I1(__766__),
    .I0(__704__),
    .O(__3334__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7497__ (
    .I1(RESET),
    .I0(__1078__),
    .O(__3335__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7498__ (
    .I1(RESET),
    .I0(__794__),
    .O(__3336__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7499__ (
    .I1(RESET),
    .I0(__505__),
    .O(__3337__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7500__ (
    .I1(RESET),
    .I0(__1365__),
    .O(__3338__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7501__ (
    .I1(RESET),
    .I0(__1443__),
    .O(__3339__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7502__ (
    .I2(RESET),
    .I1(__69__),
    .I0(__193__),
    .O(__3340__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7503__ (
    .I1(RESET),
    .I0(__1588__),
    .O(__3341__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7504__ (
    .I1(RESET),
    .I0(__462__),
    .O(__3342__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7505__ (
    .I5(TM0),
    .I4(__1393__),
    .I3(__1457__),
    .I2(__1425__),
    .I1(__1489__),
    .I0(__1326__),
    .O(__3343__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7506__ (
    .I5(TM0),
    .I4(__1201__),
    .I3(__1265__),
    .I2(__1233__),
    .I1(__1297__),
    .I0(__1169__),
    .O(__3344__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __7507__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__3344__),
    .I0(__3343__),
    .O(__3345__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7508__ (
    .I5(TM0),
    .I4(__1274__),
    .I3(__1242__),
    .I2(__1210__),
    .I1(__1306__),
    .I0(__1125__),
    .O(__3346__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7509__ (
    .I5(TM0),
    .I4(__1082__),
    .I3(__1018__),
    .I2(__1050__),
    .I1(__1114__),
    .I0(__986__),
    .O(__3347__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __7510__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__3347__),
    .I0(__3346__),
    .O(__3348__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7511__ (
    .I1(RESET),
    .I0(__1362__),
    .O(__3349__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7512__ (
    .I1(RESET),
    .I0(__1384__),
    .O(__3350__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7513__ (
    .I2(RESET),
    .I1(__1098__),
    .I0(__1140__),
    .O(__3351__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7514__ (
    .I1(RESET),
    .I0(__1594__),
    .O(__3352__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7515__ (
    .I1(RESET),
    .I0(__436__),
    .O(__3353__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7516__ (
    .I1(RESET),
    .I0(__268__),
    .O(__3354__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7517__ (
    .I1(RESET),
    .I0(__1019__),
    .O(__3355__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7518__ (
    .I1(RESET),
    .I0(__60__),
    .O(__3356__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7519__ (
    .I1(RESET),
    .I0(__57__),
    .O(__3357__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7520__ (
    .I5(TM0),
    .I4(__231__),
    .I3(__199__),
    .I2(__265__),
    .I1(__165__),
    .I0(__296__),
    .O(__3358__)
  );
  LUT6 #(
    .INIT(64'h00fff8f800000000)
  ) __7521__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__3358__),
    .I2(__3194__),
    .I1(TM0),
    .I0(__161__),
    .O(__3359__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7522__ (
    .I1(RESET),
    .I0(__1470__),
    .O(__3360__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7523__ (
    .I2(RESET),
    .I1(__921__),
    .I0(__933__),
    .O(__3361__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7524__ (
    .I1(RESET),
    .I0(__34__),
    .O(__3362__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7525__ (
    .I1(RESET),
    .I0(__471__),
    .O(__3363__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7526__ (
    .I1(RESET),
    .I0(__199__),
    .O(__3364__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7527__ (
    .I1(RESET),
    .I0(__651__),
    .O(__3365__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7528__ (
    .I1(RESET),
    .I0(__627__),
    .O(__3366__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7529__ (
    .I2(RESET),
    .I1(__517__),
    .I0(__569__),
    .O(__3367__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7530__ (
    .I2(TM0),
    .I1(__1704__),
    .I0(DATA_0_8),
    .O(__3368__)
  );
  LUT5 #(
    .INIT(32'h14414114)
  ) __7531__ (
    .I4(__1655__),
    .I3(__1623__),
    .I2(__1591__),
    .I1(__1687__),
    .I0(TM0),
    .O(__3369__)
  );
  LUT6 #(
    .INIT(64'hff88f0f000000000)
  ) __7532__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__3369__),
    .I2(__3368__),
    .I1(TM0),
    .I0(__1559__),
    .O(__3370__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7533__ (
    .I1(RESET),
    .I0(__615__),
    .O(__3371__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7534__ (
    .I5(TM0),
    .I4(__854__),
    .I3(__886__),
    .I2(__822__),
    .I1(__918__),
    .I0(__745__),
    .O(__3372__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7535__ (
    .I5(TM0),
    .I4(__694__),
    .I3(__662__),
    .I2(__726__),
    .I1(__630__),
    .I0(__598__),
    .O(__3373__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __7536__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__3373__),
    .I0(__3372__),
    .O(__3374__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7537__ (
    .I1(RESET),
    .I0(__579__),
    .O(__3375__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7538__ (
    .I1(RESET),
    .I0(__22__),
    .O(__3376__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7539__ (
    .I2(RESET),
    .I1(__1149__),
    .I0(__1089__),
    .O(__3377__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7540__ (
    .I1(RESET),
    .I0(__1076__),
    .O(__3378__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7541__ (
    .I2(RESET),
    .I1(__125__),
    .I0(__105__),
    .O(__3379__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7542__ (
    .I1(RESET),
    .I0(__809__),
    .O(__3380__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7543__ (
    .I5(TM0),
    .I4(__1245__),
    .I3(__1277__),
    .I2(__1213__),
    .I1(__1309__),
    .I0(__1122__),
    .O(__3381__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7544__ (
    .I5(TM0),
    .I4(__1085__),
    .I3(__1053__),
    .I2(__1021__),
    .I1(__1117__),
    .I0(__989__),
    .O(__3382__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __7545__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__3382__),
    .I0(__3381__),
    .O(__3383__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7546__ (
    .I1(RESET),
    .I0(__397__),
    .O(__3384__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7547__ (
    .I1(RESET),
    .I0(__1085__),
    .O(__3385__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7548__ (
    .I1(RESET),
    .I0(__498__),
    .O(__3386__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7549__ (
    .I1(RESET),
    .I0(__255__),
    .O(__3387__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7550__ (
    .I1(RESET),
    .I0(__7__),
    .O(__3388__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7551__ (
    .I1(TM0),
    .I0(__374__),
    .O(__3389__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __7552__ (
    .I5(TM1),
    .I4(__489__),
    .I3(__457__),
    .I2(__425__),
    .I1(__521__),
    .I0(TM0),
    .O(__3390__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7553__ (
    .I1(TM0),
    .I0(__127__),
    .O(__3391__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __7554__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__3391__),
    .I2(__2516__),
    .I1(__3390__),
    .I0(__3389__),
    .O(__3392__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7555__ (
    .I1(RESET),
    .I0(__1623__),
    .O(__3393__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7556__ (
    .I1(RESET),
    .I0(__135__),
    .O(__3394__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7557__ (
    .I1(RESET),
    .I0(__864__),
    .O(__3395__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7558__ (
    .I2(RESET),
    .I1(__1101__),
    .I0(__1137__),
    .O(__3396__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7559__ (
    .I1(RESET),
    .I0(__1618__),
    .O(__3397__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7560__ (
    .I2(RESET),
    .I1(__556__),
    .I0(__530__),
    .O(__3398__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7561__ (
    .I1(RESET),
    .I0(__390__),
    .O(__3399__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7562__ (
    .I1(RESET),
    .I0(__1554__),
    .O(__3400__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7563__ (
    .I1(RESET),
    .I0(__587__),
    .O(__3401__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7564__ (
    .I5(TM0),
    .I4(__440__),
    .I3(__504__),
    .I2(__472__),
    .I1(__536__),
    .I0(__359__),
    .O(__3402__)
  );
  LUT6 #(
    .INIT(64'hff880f0f00000000)
  ) __7565__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__2320__),
    .I2(__3402__),
    .I1(TM0),
    .I0(__41__),
    .O(__3403__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7566__ (
    .I1(RESET),
    .I0(__799__),
    .O(__3404__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7567__ (
    .I5(TM0),
    .I4(__824__),
    .I3(__888__),
    .I2(__856__),
    .I1(__920__),
    .I0(__743__),
    .O(__3405__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7568__ (
    .I5(TM0),
    .I4(__696__),
    .I3(__664__),
    .I2(__632__),
    .I1(__728__),
    .I0(__600__),
    .O(__3406__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __7569__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__3406__),
    .I0(__3405__),
    .O(__3407__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7570__ (
    .I2(RESET),
    .I1(__131__),
    .I0(__163__),
    .O(__3408__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7571__ (
    .I2(RESET),
    .I1(__1707__),
    .I0(__1683__),
    .O(__3409__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7572__ (
    .I1(RESET),
    .I0(__1406__),
    .O(__3410__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7573__ (
    .I2(RESET),
    .I1(__920__),
    .I0(__934__),
    .O(__3411__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7574__ (
    .I1(RESET),
    .I0(__279__),
    .O(__3412__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7575__ (
    .I1(RESET),
    .I0(__1599__),
    .O(__3413__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7576__ (
    .I1(RESET),
    .I0(__596__),
    .O(__3414__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7577__ (
    .I5(TM0),
    .I4(__857__),
    .I3(__825__),
    .I2(__889__),
    .I1(__921__),
    .I0(__742__),
    .O(__3415__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7578__ (
    .I5(TM0),
    .I4(__697__),
    .I3(__665__),
    .I2(__633__),
    .I1(__729__),
    .I0(__601__),
    .O(__3416__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __7579__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__3416__),
    .I0(__3415__),
    .O(__3417__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7580__ (
    .I5(TM0),
    .I4(__1201__),
    .I3(__1265__),
    .I2(__1233__),
    .I1(__1297__),
    .I0(__1134__),
    .O(__3418__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7581__ (
    .I5(TM0),
    .I4(__1073__),
    .I3(__1041__),
    .I2(__1009__),
    .I1(__1105__),
    .I0(__977__),
    .O(__3419__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __7582__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__3419__),
    .I0(__3418__),
    .O(__3420__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7583__ (
    .I1(RESET),
    .I0(__1256__),
    .O(__3421__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7584__ (
    .I1(RESET),
    .I0(__171__),
    .O(__3422__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7585__ (
    .I2(RESET),
    .I1(__339__),
    .I0(__363__),
    .O(__3423__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7586__ (
    .I1(TM0),
    .I0(__1528__),
    .O(__3424__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7587__ (
    .I1(TM0),
    .I0(__1351__),
    .O(__3425__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __7588__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__3425__),
    .I2(__1874__),
    .I1(__1762__),
    .I0(__3424__),
    .O(__3426__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7589__ (
    .I2(RESET),
    .I1(__939__),
    .I0(__915__),
    .O(__3427__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7590__ (
    .I1(RESET),
    .I0(__862__),
    .O(__3428__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7591__ (
    .I1(RESET),
    .I0(__386__),
    .O(__3429__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7592__ (
    .I1(RESET),
    .I0(__841__),
    .O(__3430__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7593__ (
    .I1(RESET),
    .I0(__1071__),
    .O(__3431__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7594__ (
    .I1(RESET),
    .I0(__281__),
    .O(__3432__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7595__ (
    .I5(TM0),
    .I4(__1080__),
    .I3(__1048__),
    .I2(__1016__),
    .I1(__1112__),
    .I0(__935__),
    .O(__3433__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7596__ (
    .I5(TM0),
    .I4(__824__),
    .I3(__888__),
    .I2(__856__),
    .I1(__920__),
    .I0(__792__),
    .O(__3434__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __7597__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__3434__),
    .I0(__3433__),
    .O(__3435__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7598__ (
    .I2(RESET),
    .I1(__132__),
    .I0(__191__),
    .O(__3436__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7599__ (
    .I1(TM0),
    .I0(__1338__),
    .O(__3437__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7600__ (
    .I1(TM0),
    .I0(__1157__),
    .O(__3438__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __7601__ (
    .I5(TM1),
    .I4(__1253__),
    .I3(__1221__),
    .I2(__1189__),
    .I1(__1285__),
    .I0(TM0),
    .O(__3439__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __7602__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__3439__),
    .I2(__3438__),
    .I1(__2811__),
    .I0(__3437__),
    .O(__3440__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7603__ (
    .I5(TM0),
    .I4(__1043__),
    .I3(__1075__),
    .I2(__1011__),
    .I1(__1107__),
    .I0(__940__),
    .O(__3441__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7604__ (
    .I5(TM0),
    .I4(__883__),
    .I3(__851__),
    .I2(__819__),
    .I1(__915__),
    .I0(__787__),
    .O(__3442__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __7605__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__3442__),
    .I0(__3441__),
    .O(__3443__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7606__ (
    .I1(RESET),
    .I0(__1574__),
    .O(__3444__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7607__ (
    .I1(RESET),
    .I0(__76__),
    .O(__3445__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7608__ (
    .I1(RESET),
    .I0(__1232__),
    .O(__3446__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7609__ (
    .I1(RESET),
    .I0(__1079__),
    .O(__3447__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7610__ (
    .I2(RESET),
    .I1(__1512__),
    .I0(__1494__),
    .O(__3448__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7611__ (
    .I5(TM0),
    .I4(__168__),
    .I3(__249__),
    .I2(__137__),
    .I1(__104__),
    .I0(__282__),
    .O(__3449__)
  );
  LUT6 #(
    .INIT(64'h00fff8f800000000)
  ) __7612__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__3449__),
    .I2(__3016__),
    .I1(TM0),
    .I0(__125__),
    .O(__3450__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7613__ (
    .I1(RESET),
    .I0(__1244__),
    .O(__3451__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7614__ (
    .I1(RESET),
    .I0(__170__),
    .O(__3452__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7615__ (
    .I2(RESET),
    .I1(__1709__),
    .I0(__1681__),
    .O(__3453__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7616__ (
    .I1(RESET),
    .I0(__1390__),
    .O(__3454__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7617__ (
    .I1(RESET),
    .I0(__439__),
    .O(__3455__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7618__ (
    .I1(RESET),
    .I0(__1581__),
    .O(__3456__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7619__ (
    .I1(RESET),
    .I0(__1420__),
    .O(__3457__)
  );
  LUT4 #(
    .INIT(16'h6900)
  ) __7620__ (
    .I3(RESET),
    .I2(__1727__),
    .I1(__1711__),
    .I0(__1679__),
    .O(__3458__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7621__ (
    .I2(TM0),
    .I1(__1726__),
    .I0(DATA_0_30),
    .O(__3459__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __7622__ (
    .I5(TM1),
    .I4(__1633__),
    .I3(__1601__),
    .I2(__1569__),
    .I1(__1665__),
    .I0(TM0),
    .O(__3460__)
  );
  LUT6 #(
    .INIT(64'hff88f0f000000000)
  ) __7623__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__3460__),
    .I2(__3459__),
    .I1(TM0),
    .I0(__1537__),
    .O(__3461__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7624__ (
    .I1(RESET),
    .I0(__1567__),
    .O(__3462__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7625__ (
    .I1(RESET),
    .I0(__1171__),
    .O(__3463__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7626__ (
    .I1(RESET),
    .I0(__1038__),
    .O(__3464__)
  );
  LUT4 #(
    .INIT(16'h6900)
  ) __7627__ (
    .I3(RESET),
    .I2(__106__),
    .I1(__131__),
    .I0(__75__),
    .O(__3465__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7628__ (
    .I1(RESET),
    .I0(__418__),
    .O(__3466__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7629__ (
    .I1(RESET),
    .I0(__205__),
    .O(__3467__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7630__ (
    .I1(RESET),
    .I0(__504__),
    .O(__3468__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __7631__ (
    .I1(RESET),
    .I0(__768__),
    .O(__3469__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7632__ (
    .I1(RESET),
    .I0(__815__),
    .O(__3470__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7633__ (
    .I1(RESET),
    .I0(__591__),
    .O(__3471__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7634__ (
    .I2(RESET),
    .I1(__1526__),
    .I0(__1480__),
    .O(__3472__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7635__ (
    .I2(RESET),
    .I1(__1535__),
    .I0(__1503__),
    .O(__3473__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7636__ (
    .I1(TM0),
    .I0(__766__),
    .O(__3474__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7637__ (
    .I1(TM0),
    .I0(__577__),
    .O(__3475__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __7638__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__3475__),
    .I2(__2950__),
    .I1(__3256__),
    .I0(__3474__),
    .O(__3476__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7639__ (
    .I2(RESET),
    .I1(__379__),
    .I0(__323__),
    .O(__3477__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7640__ (
    .I1(RESET),
    .I0(__261__),
    .O(__3478__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7641__ (
    .I1(RESET),
    .I0(__878__),
    .O(__3479__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7642__ (
    .I1(RESET),
    .I0(__892__),
    .O(__3480__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7643__ (
    .I1(RESET),
    .I0(__1595__),
    .O(__3481__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7644__ (
    .I5(TM0),
    .I4(__1055__),
    .I3(__1023__),
    .I2(__1087__),
    .I1(__1119__),
    .I0(__928__),
    .O(__3482__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7645__ (
    .I5(TM0),
    .I4(__895__),
    .I3(__863__),
    .I2(__831__),
    .I1(__927__),
    .I0(__799__),
    .O(__3483__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __7646__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__3483__),
    .I0(__3482__),
    .O(__3484__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7647__ (
    .I1(RESET),
    .I0(__65__),
    .O(__3485__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7648__ (
    .I1(RESET),
    .I0(__1041__),
    .O(__3486__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7649__ (
    .I2(RESET),
    .I1(__932__),
    .I0(__922__),
    .O(__3487__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7650__ (
    .I1(RESET),
    .I0(__1620__),
    .O(__3488__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7651__ (
    .I1(RESET),
    .I0(__1383__),
    .O(__3489__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7652__ (
    .I2(RESET),
    .I1(__1150__),
    .I0(__1088__),
    .O(__3490__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7653__ (
    .I1(RESET),
    .I0(__1204__),
    .O(__3491__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7654__ (
    .I1(RESET),
    .I0(__32__),
    .O(__3492__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7655__ (
    .I2(RESET),
    .I1(__327__),
    .I0(__375__),
    .O(__3493__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7656__ (
    .I1(RESET),
    .I0(__610__),
    .O(__3494__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7657__ (
    .I5(TM0),
    .I4(__479__),
    .I3(__447__),
    .I2(__511__),
    .I1(__543__),
    .I0(__352__),
    .O(__3495__)
  );
  LUT5 #(
    .INIT(32'h14414114)
  ) __7658__ (
    .I4(__29__),
    .I3(__319__),
    .I2(__39__),
    .I1(__351__),
    .I0(TM0),
    .O(__3496__)
  );
  LUT6 #(
    .INIT(64'hff880f0f00000000)
  ) __7659__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__3496__),
    .I2(__3495__),
    .I1(TM0),
    .I0(__97__),
    .O(__3497__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7660__ (
    .I1(RESET),
    .I0(__699__),
    .O(__3498__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7661__ (
    .I1(RESET),
    .I0(__840__),
    .O(__3499__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7662__ (
    .I1(RESET),
    .I0(__461__),
    .O(__3500__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7663__ (
    .I1(RESET),
    .I0(__283__),
    .O(__3501__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7664__ (
    .I2(RESET),
    .I1(__68__),
    .I0(__189__),
    .O(__3502__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7665__ (
    .I1(RESET),
    .I0(__797__),
    .O(__3503__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7666__ (
    .I2(RESET),
    .I1(__1473__),
    .I0(__1533__),
    .O(__3504__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7667__ (
    .I2(RESET),
    .I1(__1335__),
    .I0(__1287__),
    .O(__3505__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7668__ (
    .I1(TM0),
    .I0(__377__),
    .O(__3506__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7669__ (
    .I1(TM0),
    .I0(__128__),
    .O(__3507__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __7670__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__3507__),
    .I2(__2511__),
    .I1(__2218__),
    .I0(__3506__),
    .O(__3508__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7671__ (
    .I1(RESET),
    .I0(__1404__),
    .O(__3509__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7672__ (
    .I2(RESET),
    .I1(__755__),
    .I0(__715__),
    .O(__3510__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7673__ (
    .I1(RESET),
    .I0(__1602__),
    .O(__3511__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7674__ (
    .I2(TM0),
    .I1(__1708__),
    .I0(DATA_0_12),
    .O(__3512__)
  );
  LUT6 #(
    .INIT(64'hff88f0f000000000)
  ) __7675__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__3152__),
    .I2(__3512__),
    .I1(TM0),
    .I0(__1555__),
    .O(__3513__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7676__ (
    .I1(RESET),
    .I0(__1423__),
    .O(__3514__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7677__ (
    .I1(RESET),
    .I0(__654__),
    .O(__3515__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7678__ (
    .I1(RESET),
    .I0(__254__),
    .O(__3516__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7679__ (
    .I2(RESET),
    .I1(__1715__),
    .I0(__1675__),
    .O(__3517__)
  );
  LUT6 #(
    .INIT(64'h4bb4b44bb44b4bb4)
  ) __7680__ (
    .I5(__231__),
    .I4(__199__),
    .I3(__265__),
    .I2(__165__),
    .I1(TM0),
    .I0(__296__),
    .O(__3518__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7681__ (
    .I5(TM0),
    .I4(__1298__),
    .I3(__1266__),
    .I2(__1234__),
    .I1(__1202__),
    .I0(__1133__),
    .O(__3519__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7682__ (
    .I5(TM0),
    .I4(__1074__),
    .I3(__1042__),
    .I2(__1010__),
    .I1(__1106__),
    .I0(__978__),
    .O(__3520__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __7683__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__3520__),
    .I0(__3519__),
    .O(__3521__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7684__ (
    .I1(RESET),
    .I0(__620__),
    .O(__3522__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7685__ (
    .I2(RESET),
    .I1(__564__),
    .I0(__522__),
    .O(__3523__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7686__ (
    .I5(TM0),
    .I4(__925__),
    .I3(__829__),
    .I2(__861__),
    .I1(__893__),
    .I0(__738__),
    .O(__3524__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7687__ (
    .I5(TM0),
    .I4(__637__),
    .I3(__733__),
    .I2(__701__),
    .I1(__669__),
    .I0(__605__),
    .O(__3525__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __7688__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__3525__),
    .I0(__3524__),
    .O(__3526__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7689__ (
    .I1(RESET),
    .I0(__1346__),
    .O(__3527__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7690__ (
    .I1(RESET),
    .I0(__962__),
    .O(__3528__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7691__ (
    .I2(RESET),
    .I1(__1727__),
    .I0(__1695__),
    .O(__3529__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7692__ (
    .I1(RESET),
    .I0(__833__),
    .O(__3530__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7693__ (
    .I1(RESET),
    .I0(__1257__),
    .O(__3531__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7694__ (
    .I2(RESET),
    .I1(__1139__),
    .I0(__1099__),
    .O(__3532__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7695__ (
    .I1(RESET),
    .I0(__784__),
    .O(__3533__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7696__ (
    .I1(RESET),
    .I0(__108__),
    .O(__3534__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7697__ (
    .I1(RESET),
    .I0(__1643__),
    .O(__3535__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __7698__ (
    .I1(RESET),
    .I0(__1536__),
    .O(__3536__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7699__ (
    .I1(RESET),
    .I0(__271__),
    .O(__3537__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7700__ (
    .I2(RESET),
    .I1(__155__),
    .I0(__166__),
    .O(__3538__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7701__ (
    .I1(RESET),
    .I0(__702__),
    .O(__3539__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7702__ (
    .I5(TM0),
    .I4(__258__),
    .I3(__197__),
    .I2(__224__),
    .I1(__163__),
    .I0(__289__),
    .O(__3540__)
  );
  LUT6 #(
    .INIT(64'h00fff8f800000000)
  ) __7703__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__3540__),
    .I2(__3496__),
    .I1(TM0),
    .I0(__146__),
    .O(__3541__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7704__ (
    .I1(RESET),
    .I0(__45__),
    .O(__3542__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7705__ (
    .I1(RESET),
    .I0(__1451__),
    .O(__3543__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7706__ (
    .I2(RESET),
    .I1(__958__),
    .I0(__896__),
    .O(__3544__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7707__ (
    .I1(RESET),
    .I0(__998__),
    .O(__3545__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7708__ (
    .I1(RESET),
    .I0(__1551__),
    .O(__3546__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7709__ (
    .I1(RESET),
    .I0(__1241__),
    .O(__3547__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7710__ (
    .I1(RESET),
    .I0(__97__),
    .O(__3548__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7711__ (
    .I1(RESET),
    .I0(__1248__),
    .O(__3549__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7712__ (
    .I2(RESET),
    .I1(__574__),
    .I0(__512__),
    .O(__3550__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7713__ (
    .I1(RESET),
    .I0(__1225__),
    .O(__3551__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7714__ (
    .I1(RESET),
    .I0(__1435__),
    .O(__3552__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7715__ (
    .I1(RESET),
    .I0(__222__),
    .O(__3553__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7716__ (
    .I1(RESET),
    .I0(__1629__),
    .O(__3554__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7717__ (
    .I1(RESET),
    .I0(__186__),
    .O(__3555__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7718__ (
    .I1(RESET),
    .I0(__1238__),
    .O(__3556__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7719__ (
    .I2(RESET),
    .I1(__1090__),
    .I0(__1148__),
    .O(__3557__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7720__ (
    .I2(RESET),
    .I1(__913__),
    .I0(__941__),
    .O(__3558__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7721__ (
    .I1(RESET),
    .I0(__59__),
    .O(__3559__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7722__ (
    .I1(RESET),
    .I0(__248__),
    .O(__3560__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7723__ (
    .I2(RESET),
    .I1(__366__),
    .I0(__336__),
    .O(__3561__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7724__ (
    .I1(RESET),
    .I0(__1208__),
    .O(__3562__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7725__ (
    .I1(TM0),
    .I0(__1520__),
    .O(__3563__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7726__ (
    .I1(TM0),
    .I0(__1359__),
    .O(__3564__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __7727__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__3564__),
    .I2(__2144__),
    .I1(__1919__),
    .I0(__3563__),
    .O(__3565__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7728__ (
    .I1(TM0),
    .I0(__1342__),
    .O(__3566__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __7729__ (
    .I5(TM1),
    .I4(__1377__),
    .I3(__1441__),
    .I2(__1409__),
    .I1(__1473__),
    .I0(TM0),
    .O(__3567__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7730__ (
    .I1(TM0),
    .I0(__1153__),
    .O(__3568__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __7731__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__3568__),
    .I2(__2270__),
    .I1(__3567__),
    .I0(__3566__),
    .O(__3569__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7732__ (
    .I1(RESET),
    .I0(__630__),
    .O(__3570__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7733__ (
    .I2(RESET),
    .I1(__360__),
    .I0(__342__),
    .O(__3571__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7734__ (
    .I1(RESET),
    .I0(__578__),
    .O(__3572__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7735__ (
    .I1(RESET),
    .I0(__130__),
    .O(__3573__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7736__ (
    .I1(RESET),
    .I0(__138__),
    .O(__3574__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7737__ (
    .I1(RESET),
    .I0(__249__),
    .O(__3575__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7738__ (
    .I2(RESET),
    .I1(__1331__),
    .I0(__1291__),
    .O(__3576__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7739__ (
    .I2(RESET),
    .I1(__952__),
    .I0(__902__),
    .O(__3577__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7740__ (
    .I2(RESET),
    .I1(__950__),
    .I0(__904__),
    .O(__3578__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7741__ (
    .I2(RESET),
    .I1(__1341__),
    .I0(__1281__),
    .O(__3579__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7742__ (
    .I1(RESET),
    .I0(__1552__),
    .O(__3580__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7743__ (
    .I2(RESET),
    .I1(__1091__),
    .I0(__1147__),
    .O(__3581__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7744__ (
    .I1(RESET),
    .I0(__1441__),
    .O(__3582__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7745__ (
    .I1(RESET),
    .I0(__1179__),
    .O(__3583__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7746__ (
    .I1(RESET),
    .I0(__1050__),
    .O(__3584__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7747__ (
    .I1(RESET),
    .I0(__207__),
    .O(__3585__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7748__ (
    .I1(RESET),
    .I0(__17__),
    .O(__3586__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __7749__ (
    .I2(TM0),
    .I1(__1699__),
    .I0(DATA_0_3),
    .O(__3587__)
  );
  LUT5 #(
    .INIT(32'h14414114)
  ) __7750__ (
    .I4(__1660__),
    .I3(__1628__),
    .I2(__1596__),
    .I1(__1692__),
    .I0(TM0),
    .O(__3588__)
  );
  LUT6 #(
    .INIT(64'hff88f0f000000000)
  ) __7751__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__3588__),
    .I2(__3587__),
    .I1(TM0),
    .I0(__1564__),
    .O(__3589__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7752__ (
    .I1(RESET),
    .I0(__997__),
    .O(__3590__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7753__ (
    .I1(RESET),
    .I0(__476__),
    .O(__3591__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7754__ (
    .I1(RESET),
    .I0(__885__),
    .O(__3592__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7755__ (
    .I1(RESET),
    .I0(__1401__),
    .O(__3593__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7756__ (
    .I1(RESET),
    .I0(__1562__),
    .O(__3594__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7757__ (
    .I1(RESET),
    .I0(__1069__),
    .O(__3595__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7758__ (
    .I1(RESET),
    .I0(__886__),
    .O(__3596__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7759__ (
    .I1(TM0),
    .I0(__946__),
    .O(__3597__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __7760__ (
    .I5(TM1),
    .I4(__1069__),
    .I3(__1037__),
    .I2(__1005__),
    .I1(__1101__),
    .I0(TM0),
    .O(__3598__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7761__ (
    .I1(TM0),
    .I0(__781__),
    .O(__3599__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __7762__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__3599__),
    .I2(__2646__),
    .I1(__3598__),
    .I0(__3597__),
    .O(__3600__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __7763__ (
    .I1(RESET),
    .I0(__112__),
    .O(__3601__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7764__ (
    .I1(TM0),
    .I0(__761__),
    .O(__3602__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7765__ (
    .I1(TM0),
    .I0(__582__),
    .O(__3603__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __7766__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__3603__),
    .I2(__2216__),
    .I1(__2410__),
    .I0(__3602__),
    .O(__3604__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7767__ (
    .I1(RESET),
    .I0(__1006__),
    .O(__3605__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7768__ (
    .I1(TM0),
    .I0(__560__),
    .O(__3606__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7769__ (
    .I1(TM0),
    .I0(__399__),
    .O(__3607__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __7770__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__3607__),
    .I2(__3102__),
    .I1(__2507__),
    .I0(__3606__),
    .O(__3608__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7771__ (
    .I1(RESET),
    .I0(__420__),
    .O(__3609__)
  );
  LUT6 #(
    .INIT(64'h6996966996696996)
  ) __7772__ (
    .I5(TM1),
    .I4(__172__),
    .I3(__134__),
    .I2(__141__),
    .I1(__205__),
    .I0(__2396__),
    .O(__3610__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7773__ (
    .I1(RESET),
    .I0(__1630__),
    .O(__3611__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7774__ (
    .I1(RESET),
    .I0(__1255__),
    .O(__3612__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7775__ (
    .I2(RESET),
    .I1(__738__),
    .I0(__732__),
    .O(__3613__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7776__ (
    .I1(TM0),
    .I0(__566__),
    .O(__3614__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7777__ (
    .I1(TM0),
    .I0(__393__),
    .O(__3615__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __7778__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__3615__),
    .I2(__3390__),
    .I1(__2753__),
    .I0(__3614__),
    .O(__3616__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7779__ (
    .I1(RESET),
    .I0(__853__),
    .O(__3617__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7780__ (
    .I1(RESET),
    .I0(__413__),
    .O(__3618__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7781__ (
    .I1(RESET),
    .I0(__684__),
    .O(__3619__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7782__ (
    .I1(RESET),
    .I0(__1387__),
    .O(__3620__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7783__ (
    .I2(RESET),
    .I1(__1697__),
    .I0(__1693__),
    .O(__3621__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7784__ (
    .I5(TM0),
    .I4(__533__),
    .I3(__469__),
    .I2(__501__),
    .I1(__437__),
    .I0(__362__),
    .O(__3622__)
  );
  LUT6 #(
    .INIT(64'hff880f0f00000000)
  ) __7785__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__1888__),
    .I2(__3622__),
    .I1(TM0),
    .I0(__44__),
    .O(__3623__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7786__ (
    .I1(RESET),
    .I0(__850__),
    .O(__3624__)
  );
  LUT4 #(
    .INIT(16'h6900)
  ) __7787__ (
    .I3(RESET),
    .I2(__575__),
    .I1(__559__),
    .I0(__527__),
    .O(__3625__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7788__ (
    .I1(RESET),
    .I0(__1227__),
    .O(__3626__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7789__ (
    .I1(RESET),
    .I0(__1193__),
    .O(__3627__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7790__ (
    .I1(RESET),
    .I0(__617__),
    .O(__3628__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7791__ (
    .I1(RESET),
    .I0(__606__),
    .O(__3629__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7792__ (
    .I1(RESET),
    .I0(__1259__),
    .O(__3630__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7793__ (
    .I1(RESET),
    .I0(__971__),
    .O(__3631__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7794__ (
    .I1(RESET),
    .I0(__312__),
    .O(__3632__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7795__ (
    .I1(RESET),
    .I0(__1553__),
    .O(__3633__)
  );
  LUT6 #(
    .INIT(64'h6996966996696996)
  ) __7796__ (
    .I5(TM1),
    .I4(__293__),
    .I3(__228__),
    .I2(__261__),
    .I1(__195__),
    .I0(__2186__),
    .O(__3634__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7797__ (
    .I1(TM0),
    .I0(__952__),
    .O(__3635__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7798__ (
    .I1(TM0),
    .I0(__775__),
    .O(__3636__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __7799__ (
    .I5(TM1),
    .I4(__839__),
    .I3(__871__),
    .I2(__807__),
    .I1(__903__),
    .I0(TM0),
    .O(__3637__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __7800__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__3637__),
    .I2(__3636__),
    .I1(__1980__),
    .I0(__3635__),
    .O(__3638__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7801__ (
    .I1(RESET),
    .I0(__668__),
    .O(__3639__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7802__ (
    .I1(RESET),
    .I0(__1654__),
    .O(__3640__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7803__ (
    .I2(RESET),
    .I1(__717__),
    .I0(__753__),
    .O(__3641__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7804__ (
    .I1(RESET),
    .I0(__619__),
    .O(__3642__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7805__ (
    .I1(RESET),
    .I0(__1036__),
    .O(__3643__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7806__ (
    .I1(RESET),
    .I0(__169__),
    .O(__3644__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7807__ (
    .I1(RESET),
    .I0(__1063__),
    .O(__3645__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7808__ (
    .I1(RESET),
    .I0(__1025__),
    .O(__3646__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7809__ (
    .I1(RESET),
    .I0(__43__),
    .O(__3647__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7810__ (
    .I1(RESET),
    .I0(__992__),
    .O(__3648__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7811__ (
    .I1(RESET),
    .I0(__83__),
    .O(__3649__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7812__ (
    .I1(RESET),
    .I0(__976__),
    .O(__3650__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7813__ (
    .I1(RESET),
    .I0(__276__),
    .O(__3651__)
  );
  LUT4 #(
    .INIT(16'h6900)
  ) __7814__ (
    .I3(RESET),
    .I2(__1727__),
    .I1(__1691__),
    .I0(__1699__),
    .O(__3652__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7815__ (
    .I1(RESET),
    .I0(__1011__),
    .O(__3653__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7816__ (
    .I1(RESET),
    .I0(__180__),
    .O(__3654__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7817__ (
    .I1(RESET),
    .I0(__284__),
    .O(__3655__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7818__ (
    .I1(RESET),
    .I0(__225__),
    .O(__3656__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7819__ (
    .I1(RESET),
    .I0(__223__),
    .O(__3657__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7820__ (
    .I1(TM0),
    .I0(__561__),
    .O(__3658__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7821__ (
    .I1(TM0),
    .I0(__398__),
    .O(__3659__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __7822__ (
    .I5(TM1),
    .I4(__494__),
    .I3(__462__),
    .I2(__430__),
    .I1(__526__),
    .I0(TM0),
    .O(__3660__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __7823__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__3660__),
    .I2(__3659__),
    .I1(__2240__),
    .I0(__3658__),
    .O(__3661__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7824__ (
    .I1(RESET),
    .I0(__1460__),
    .O(__3662__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7825__ (
    .I5(TM0),
    .I4(__1203__),
    .I3(__1267__),
    .I2(__1235__),
    .I1(__1299__),
    .I0(__1132__),
    .O(__3663__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7826__ (
    .I5(TM0),
    .I4(__1043__),
    .I3(__1075__),
    .I2(__1011__),
    .I1(__1107__),
    .I0(__979__),
    .O(__3664__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __7827__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__3664__),
    .I0(__3663__),
    .O(__3665__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7828__ (
    .I2(RESET),
    .I1(__346__),
    .I0(__356__),
    .O(__3666__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7829__ (
    .I1(RESET),
    .I0(__1044__),
    .O(__3667__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7830__ (
    .I1(RESET),
    .I0(__696__),
    .O(__3668__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7831__ (
    .I2(RESET),
    .I1(__744__),
    .I0(__726__),
    .O(__3669__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7832__ (
    .I1(TM0),
    .I0(__954__),
    .O(__3670__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __7833__ (
    .I5(TM1),
    .I4(__1061__),
    .I3(__1029__),
    .I2(__997__),
    .I1(__1093__),
    .I0(TM0),
    .O(__3671__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7834__ (
    .I1(TM0),
    .I0(__773__),
    .O(__3672__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __7835__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__3672__),
    .I2(__2176__),
    .I1(__3671__),
    .I0(__3670__),
    .O(__3673__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7836__ (
    .I5(TM0),
    .I4(__696__),
    .I3(__664__),
    .I2(__632__),
    .I1(__728__),
    .I0(__551__),
    .O(__3674__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7837__ (
    .I5(TM0),
    .I4(__440__),
    .I3(__504__),
    .I2(__472__),
    .I1(__536__),
    .I0(__408__),
    .O(__3675__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __7838__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__3675__),
    .I0(__3674__),
    .O(__3676__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7839__ (
    .I2(RESET),
    .I1(__1522__),
    .I0(__1484__),
    .O(__3677__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7840__ (
    .I1(RESET),
    .I0(__39__),
    .O(__3678__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7841__ (
    .I1(RESET),
    .I0(__1638__),
    .O(__3679__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7842__ (
    .I1(RESET),
    .I0(__1250__),
    .O(__3680__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7843__ (
    .I5(TM0),
    .I4(__1264__),
    .I3(__1232__),
    .I2(__1200__),
    .I1(__1296__),
    .I0(__1135__),
    .O(__3681__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7844__ (
    .I5(TM0),
    .I4(__1008__),
    .I3(__1040__),
    .I2(__1072__),
    .I1(__1104__),
    .I0(__976__),
    .O(__3682__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __7845__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__3682__),
    .I0(__3681__),
    .O(__3683__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7846__ (
    .I1(RESET),
    .I0(__16__),
    .O(__3684__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7847__ (
    .I1(RESET),
    .I0(__212__),
    .O(__3685__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7848__ (
    .I1(RESET),
    .I0(__968__),
    .O(__3686__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7849__ (
    .I2(RESET),
    .I1(__107__),
    .I0(__74__),
    .O(__3687__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7850__ (
    .I1(RESET),
    .I0(__292__),
    .O(__3688__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7851__ (
    .I2(RESET),
    .I1(__765__),
    .I0(__705__),
    .O(__3689__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7852__ (
    .I1(RESET),
    .I0(__673__),
    .O(__3690__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7853__ (
    .I1(RESET),
    .I0(__52__),
    .O(__3691__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7854__ (
    .I1(RESET),
    .I0(__825__),
    .O(__3692__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7855__ (
    .I1(TM0),
    .I0(__1534__),
    .O(__3693__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7856__ (
    .I1(TM0),
    .I0(__1345__),
    .O(__3694__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __7857__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__3694__),
    .I2(__3567__),
    .I1(__3460__),
    .I0(__3693__),
    .O(__3695__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7858__ (
    .I1(RESET),
    .I0(__1182__),
    .O(__3696__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7859__ (
    .I1(RESET),
    .I0(__440__),
    .O(__3697__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7860__ (
    .I1(RESET),
    .I0(__1212__),
    .O(__3698__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7861__ (
    .I1(TM0),
    .I0(__1146__),
    .O(__3699__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7862__ (
    .I1(TM0),
    .I0(__965__),
    .O(__3700__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __7863__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__3700__),
    .I2(__3671__),
    .I1(__3439__),
    .I0(__3699__),
    .O(__3701__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7864__ (
    .I1(RESET),
    .I0(__834__),
    .O(__3702__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7865__ (
    .I1(RESET),
    .I0(__278__),
    .O(__3703__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7866__ (
    .I2(RESET),
    .I1(__73__),
    .I0(__134__),
    .O(__3704__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7867__ (
    .I2(RESET),
    .I1(__1496__),
    .I0(__1510__),
    .O(__3705__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7868__ (
    .I1(RESET),
    .I0(__1467__),
    .O(__3706__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7869__ (
    .I1(TM0),
    .I0(__1523__),
    .O(__3707__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7870__ (
    .I1(TM0),
    .I0(__1356__),
    .O(__3708__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __7871__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__3708__),
    .I2(__1848__),
    .I1(__1943__),
    .I0(__3707__),
    .O(__3709__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7872__ (
    .I1(RESET),
    .I0(__1628__),
    .O(__3710__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7873__ (
    .I1(RESET),
    .I0(__791__),
    .O(__3711__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7874__ (
    .I2(RESET),
    .I1(__159__),
    .I0(__103__),
    .O(__3712__)
  );
  LUT4 #(
    .INIT(16'h6900)
  ) __7875__ (
    .I3(RESET),
    .I2(__367__),
    .I1(__383__),
    .I0(__335__),
    .O(__3713__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7876__ (
    .I1(RESET),
    .I0(__1377__),
    .O(__3714__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7877__ (
    .I1(RESET),
    .I0(__1559__),
    .O(__3715__)
  );
  LUT6 #(
    .INIT(64'h4bb4b44bb44b4bb4)
  ) __7878__ (
    .I5(__200__),
    .I4(__232__),
    .I3(__266__),
    .I2(__166__),
    .I1(TM0),
    .I0(__297__),
    .O(__3716__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7879__ (
    .I1(RESET),
    .I0(__650__),
    .O(__3717__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7880__ (
    .I1(RESET),
    .I0(__592__),
    .O(__3718__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7881__ (
    .I1(RESET),
    .I0(__231__),
    .O(__3719__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7882__ (
    .I1(RESET),
    .I0(__1394__),
    .O(__3720__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7883__ (
    .I1(RESET),
    .I0(__1262__),
    .O(__3721__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7884__ (
    .I1(RESET),
    .I0(__1357__),
    .O(__3722__)
  );
  LUT4 #(
    .INIT(16'h6900)
  ) __7885__ (
    .I3(RESET),
    .I2(__1315__),
    .I1(__1307__),
    .I0(__1343__),
    .O(__3723__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7886__ (
    .I1(RESET),
    .I0(__1205__),
    .O(__3724__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7887__ (
    .I1(RESET),
    .I0(__127__),
    .O(__3725__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7888__ (
    .I1(RESET),
    .I0(__1023__),
    .O(__3726__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7889__ (
    .I1(RESET),
    .I0(__774__),
    .O(__3727__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7890__ (
    .I1(RESET),
    .I0(__1381__),
    .O(__3728__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7891__ (
    .I2(RESET),
    .I1(__525__),
    .I0(__561__),
    .O(__3729__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7892__ (
    .I1(RESET),
    .I0(__313__),
    .O(__3730__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7893__ (
    .I2(RESET),
    .I1(__1129__),
    .I0(__1109__),
    .O(__3731__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7894__ (
    .I1(RESET),
    .I0(__6__),
    .O(__3732__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7895__ (
    .I1(RESET),
    .I0(__1197__),
    .O(__3733__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7896__ (
    .I1(RESET),
    .I0(__776__),
    .O(__3734__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7897__ (
    .I5(TM0),
    .I4(__1236__),
    .I3(__1268__),
    .I2(__1204__),
    .I1(__1300__),
    .I0(__1131__),
    .O(__3735__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7898__ (
    .I5(TM0),
    .I4(__1076__),
    .I3(__1044__),
    .I2(__1012__),
    .I1(__1108__),
    .I0(__980__),
    .O(__3736__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __7899__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__3736__),
    .I0(__3735__),
    .O(__3737__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7900__ (
    .I1(RESET),
    .I0(__1446__),
    .O(__3738__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7901__ (
    .I1(RESET),
    .I0(__1013__),
    .O(__3739__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7902__ (
    .I1(RESET),
    .I0(__1032__),
    .O(__3740__)
  );
  LUT5 #(
    .INIT(32'h14414114)
  ) __7903__ (
    .I4(__1598__),
    .I3(__1662__),
    .I2(__1630__),
    .I1(__1694__),
    .I0(TM0),
    .O(__3741__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7904__ (
    .I5(TM0),
    .I4(__1470__),
    .I3(__1438__),
    .I2(__1406__),
    .I1(__1502__),
    .I0(__1374__),
    .O(__3742__)
  );
  LUT6 #(
    .INIT(64'h00fff8f800000000)
  ) __7905__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__3742__),
    .I2(__3741__),
    .I1(TM0),
    .I0(__1505__),
    .O(__3743__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7906__ (
    .I2(RESET),
    .I1(__113__),
    .I0(__178__),
    .O(__3744__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7907__ (
    .I1(RESET),
    .I0(__245__),
    .O(__3745__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7908__ (
    .I1(RESET),
    .I0(__991__),
    .O(__3746__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7909__ (
    .I1(RESET),
    .I0(__1278__),
    .O(__3747__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7910__ (
    .I5(TM0),
    .I4(__510__),
    .I3(__478__),
    .I2(__446__),
    .I1(__542__),
    .I0(__353__),
    .O(__3748__)
  );
  LUT6 #(
    .INIT(64'hff880f0f00000000)
  ) __7911__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__2578__),
    .I2(__3748__),
    .I1(TM0),
    .I0(__85__),
    .O(__3749__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7912__ (
    .I1(RESET),
    .I0(__1639__),
    .O(__3750__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7913__ (
    .I1(RESET),
    .I0(__1597__),
    .O(__3751__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7914__ (
    .I1(RESET),
    .I0(__1444__),
    .O(__3752__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7915__ (
    .I2(RESET),
    .I1(__325__),
    .I0(__377__),
    .O(__3753__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7916__ (
    .I5(TM0),
    .I4(__499__),
    .I3(__467__),
    .I2(__435__),
    .I1(__531__),
    .I0(__364__),
    .O(__3754__)
  );
  LUT6 #(
    .INIT(64'hff880f0f00000000)
  ) __7917__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__2806__),
    .I2(__3754__),
    .I1(TM0),
    .I0(__46__),
    .O(__3755__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7918__ (
    .I2(RESET),
    .I1(__1333__),
    .I0(__1289__),
    .O(__3756__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7919__ (
    .I1(RESET),
    .I0(__622__),
    .O(__3757__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7920__ (
    .I1(RESET),
    .I0(__497__),
    .O(__3758__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7921__ (
    .I1(RESET),
    .I0(__1084__),
    .O(__3759__)
  );
  LUT4 #(
    .INIT(16'h6900)
  ) __7922__ (
    .I3(RESET),
    .I2(__539__),
    .I1(__547__),
    .I0(__575__),
    .O(__3760__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7923__ (
    .I1(RESET),
    .I0(__494__),
    .O(__3761__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7924__ (
    .I1(RESET),
    .I0(__1007__),
    .O(__3762__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7925__ (
    .I1(RESET),
    .I0(__703__),
    .O(__3763__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7926__ (
    .I1(RESET),
    .I0(__801__),
    .O(__3764__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7927__ (
    .I2(RESET),
    .I1(__737__),
    .I0(__733__),
    .O(__3765__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7928__ (
    .I1(RESET),
    .I0(__1251__),
    .O(__3766__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7929__ (
    .I1(RESET),
    .I0(__604__),
    .O(__3767__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7930__ (
    .I1(RESET),
    .I0(__676__),
    .O(__3768__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7931__ (
    .I1(RESET),
    .I0(__1565__),
    .O(__3769__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7932__ (
    .I1(RESET),
    .I0(__293__),
    .O(__3770__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7933__ (
    .I1(RESET),
    .I0(__1055__),
    .O(__3771__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7934__ (
    .I1(TM0),
    .I0(__760__),
    .O(__3772__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7935__ (
    .I1(TM0),
    .I0(__583__),
    .O(__3773__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __7936__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__3773__),
    .I2(__2614__),
    .I1(__3637__),
    .I0(__3772__),
    .O(__3774__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7937__ (
    .I5(TM0),
    .I4(__823__),
    .I3(__887__),
    .I2(__855__),
    .I1(__919__),
    .I0(__744__),
    .O(__3775__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7938__ (
    .I5(TM0),
    .I4(__695__),
    .I3(__663__),
    .I2(__631__),
    .I1(__727__),
    .I0(__599__),
    .O(__3776__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __7939__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__3776__),
    .I0(__3775__),
    .O(__3777__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7940__ (
    .I1(RESET),
    .I0(__501__),
    .O(__3778__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7941__ (
    .I1(RESET),
    .I0(__37__),
    .O(__3779__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7942__ (
    .I2(RESET),
    .I1(__1712__),
    .I0(__1678__),
    .O(__3780__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7943__ (
    .I5(TM0),
    .I4(__1275__),
    .I3(__1243__),
    .I2(__1211__),
    .I1(__1307__),
    .I0(__1124__),
    .O(__3781__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7944__ (
    .I5(TM0),
    .I4(__1083__),
    .I3(__1051__),
    .I2(__1019__),
    .I1(__1115__),
    .I0(__987__),
    .O(__3782__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __7945__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__3782__),
    .I0(__3781__),
    .O(__3783__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7946__ (
    .I5(TM0),
    .I4(__1432__),
    .I3(__1464__),
    .I2(__1400__),
    .I1(__1496__),
    .I0(__1368__),
    .O(__3784__)
  );
  LUT6 #(
    .INIT(64'h00fff8f800000000)
  ) __7947__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__3784__),
    .I2(__2847__),
    .I1(TM0),
    .I0(__1511__),
    .O(__3785__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7948__ (
    .I2(RESET),
    .I1(__1324__),
    .I0(__1298__),
    .O(__3786__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7949__ (
    .I1(RESET),
    .I0(__781__),
    .O(__3787__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7950__ (
    .I1(TM0),
    .I0(__69__),
    .O(__3788__)
  );
  LUT5 #(
    .INIT(32'h41141441)
  ) __7951__ (
    .I4(__208__),
    .I3(__175__),
    .I2(__225__),
    .I1(__201__),
    .I0(TM0),
    .O(__3789__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __7952__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__3789__),
    .I2(__2118__),
    .I1(__2166__),
    .I0(__3788__),
    .O(__3790__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7953__ (
    .I2(RESET),
    .I1(__1680__),
    .I0(__1710__),
    .O(__3791__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7954__ (
    .I1(TM0),
    .I0(__1149__),
    .O(__3792__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7955__ (
    .I1(TM0),
    .I0(__962__),
    .O(__3793__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __7956__ (
    .I5(TM1),
    .I4(__1058__),
    .I3(__1026__),
    .I2(__994__),
    .I1(__1090__),
    .I0(TM0),
    .O(__3794__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __7957__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__3794__),
    .I2(__3793__),
    .I1(__2843__),
    .I0(__3792__),
    .O(__3795__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7958__ (
    .I1(RESET),
    .I0(__447__),
    .O(__3796__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7959__ (
    .I1(TM0),
    .I0(__131__),
    .O(__3797__)
  );
  LUT5 #(
    .INIT(32'h41141441)
  ) __7960__ (
    .I4(__229__),
    .I3(__262__),
    .I2(__294__),
    .I1(__196__),
    .I0(TM0),
    .O(__3798__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __7961__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__3798__),
    .I2(__3236__),
    .I1(__3082__),
    .I0(__3797__),
    .O(__3799__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7962__ (
    .I1(RESET),
    .I0(__1607__),
    .O(__3800__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7963__ (
    .I1(RESET),
    .I0(__985__),
    .O(__3801__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7964__ (
    .I1(RESET),
    .I0(__64__),
    .O(__3802__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7965__ (
    .I1(RESET),
    .I0(__469__),
    .O(__3803__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7966__ (
    .I1(RESET),
    .I0(__1018__),
    .O(__3804__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7967__ (
    .I1(RESET),
    .I0(__581__),
    .O(__3805__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7968__ (
    .I1(RESET),
    .I0(__981__),
    .O(__3806__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7969__ (
    .I1(RESET),
    .I0(__662__),
    .O(__3807__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7970__ (
    .I1(RESET),
    .I0(__204__),
    .O(__3808__)
  );
  LUT6 #(
    .INIT(64'h4bb4b44bb44b4bb4)
  ) __7971__ (
    .I5(__185__),
    .I4(__219__),
    .I3(__251__),
    .I2(__153__),
    .I1(TM0),
    .I0(__284__),
    .O(__3809__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7972__ (
    .I1(RESET),
    .I0(__1635__),
    .O(__3810__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7973__ (
    .I1(RESET),
    .I0(__1361__),
    .O(__3811__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7974__ (
    .I2(RESET),
    .I1(__1694__),
    .I0(__1696__),
    .O(__3812__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7975__ (
    .I1(RESET),
    .I0(__966__),
    .O(__3813__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7976__ (
    .I1(RESET),
    .I0(__1236__),
    .O(__3814__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7977__ (
    .I1(RESET),
    .I0(__210__),
    .O(__3815__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7978__ (
    .I1(RESET),
    .I0(__691__),
    .O(__3816__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7979__ (
    .I1(RESET),
    .I0(__1002__),
    .O(__3817__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7980__ (
    .I1(RESET),
    .I0(__854__),
    .O(__3818__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7981__ (
    .I1(RESET),
    .I0(__839__),
    .O(__3819__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7982__ (
    .I1(RESET),
    .I0(__1393__),
    .O(__3820__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7983__ (
    .I2(RESET),
    .I1(__1687__),
    .I0(__1703__),
    .O(__3821__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7984__ (
    .I1(RESET),
    .I0(__1614__),
    .O(__3822__)
  );
  LUT5 #(
    .INIT(32'h14414114)
  ) __7985__ (
    .I4(__1652__),
    .I3(__1620__),
    .I2(__1588__),
    .I1(__1684__),
    .I0(TM0),
    .O(__3823__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __7986__ (
    .I5(TM0),
    .I4(__1460__),
    .I3(__1428__),
    .I2(__1396__),
    .I1(__1492__),
    .I0(__1364__),
    .O(__3824__)
  );
  LUT6 #(
    .INIT(64'h00fff8f800000000)
  ) __7987__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__3824__),
    .I2(__3823__),
    .I1(TM0),
    .I0(__1515__),
    .O(__3825__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7988__ (
    .I1(RESET),
    .I0(__46__),
    .O(__3826__)
  );
  LUT2 #(
    .INIT(4'h4)
  ) __7989__ (
    .I1(RESET),
    .I0(__1344__),
    .O(__3827__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7990__ (
    .I1(RESET),
    .I0(__11__),
    .O(__3828__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7991__ (
    .I1(RESET),
    .I0(__984__),
    .O(__3829__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7992__ (
    .I1(RESET),
    .I0(__1642__),
    .O(__3830__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7993__ (
    .I1(TM0),
    .I0(__1147__),
    .O(__3831__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7994__ (
    .I1(TM0),
    .I0(__964__),
    .O(__3832__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __7995__ (
    .I5(TM1),
    .I4(__1060__),
    .I3(__1028__),
    .I2(__996__),
    .I1(__1092__),
    .I0(TM0),
    .O(__3833__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __7996__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__3833__),
    .I2(__3832__),
    .I1(__1953__),
    .I0(__3831__),
    .O(__3834__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7997__ (
    .I1(RESET),
    .I0(__1045__),
    .O(__3835__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __7998__ (
    .I1(RESET),
    .I0(__1563__),
    .O(__3836__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __7999__ (
    .I2(RESET),
    .I1(__1144__),
    .I0(__1094__),
    .O(__3837__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __8000__ (
    .I2(RESET),
    .I1(__1513__),
    .I0(__1493__),
    .O(__3838__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8001__ (
    .I1(RESET),
    .I0(__256__),
    .O(__3839__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8002__ (
    .I1(RESET),
    .I0(__252__),
    .O(__3840__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8003__ (
    .I1(RESET),
    .I0(__94__),
    .O(__3841__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8004__ (
    .I1(RESET),
    .I0(__648__),
    .O(__3842__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __8005__ (
    .I2(RESET),
    .I1(__160__),
    .I0(__100__),
    .O(__3843__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __8006__ (
    .I5(TM0),
    .I4(__884__),
    .I3(__852__),
    .I2(__820__),
    .I1(__916__),
    .I0(__747__),
    .O(__3844__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __8007__ (
    .I5(TM0),
    .I4(__692__),
    .I3(__660__),
    .I2(__628__),
    .I1(__724__),
    .I0(__596__),
    .O(__3845__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __8008__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__3845__),
    .I0(__3844__),
    .O(__3846__)
  );
  LUT6 #(
    .INIT(64'h6996966996696996)
  ) __8009__ (
    .I5(TM1),
    .I4(__140__),
    .I3(__171__),
    .I2(__204__),
    .I1(__107__),
    .I0(__1863__),
    .O(__3847__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8010__ (
    .I1(RESET),
    .I0(__464__),
    .O(__3848__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8011__ (
    .I1(RESET),
    .I0(__1636__),
    .O(__3849__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8012__ (
    .I1(RESET),
    .I0(__828__),
    .O(__3850__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8013__ (
    .I1(RESET),
    .I0(__110__),
    .O(__3851__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8014__ (
    .I1(RESET),
    .I0(__395__),
    .O(__3852__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8015__ (
    .I1(RESET),
    .I0(__1570__),
    .O(__3853__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8016__ (
    .I1(RESET),
    .I0(__1469__),
    .O(__3854__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8017__ (
    .I1(RESET),
    .I0(__1348__),
    .O(__3855__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __8018__ (
    .I2(RESET),
    .I1(__526__),
    .I0(__560__),
    .O(__3856__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8019__ (
    .I1(RESET),
    .I0(__507__),
    .O(__3857__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8020__ (
    .I1(RESET),
    .I0(__56__),
    .O(__3858__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8021__ (
    .I1(RESET),
    .I0(__242__),
    .O(__3859__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8022__ (
    .I1(RESET),
    .I0(__270__),
    .O(__3860__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __8023__ (
    .I2(RESET),
    .I1(__1714__),
    .I0(__1676__),
    .O(__3861__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __8024__ (
    .I2(TM0),
    .I1(__1707__),
    .I0(DATA_0_11),
    .O(__3862__)
  );
  LUT6 #(
    .INIT(64'hff88f0f000000000)
  ) __8025__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__3823__),
    .I2(__3862__),
    .I1(TM0),
    .I0(__1556__),
    .O(__3863__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8026__ (
    .I1(RESET),
    .I0(__1351__),
    .O(__3864__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8027__ (
    .I1(RESET),
    .I0(__1073__),
    .O(__3865__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8028__ (
    .I1(RESET),
    .I0(__883__),
    .O(__3866__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8029__ (
    .I1(RESET),
    .I0(__1608__),
    .O(__3867__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8030__ (
    .I1(RESET),
    .I0(__873__),
    .O(__3868__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __8031__ (
    .I2(RESET),
    .I1(__1340__),
    .I0(__1282__),
    .O(__3869__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8032__ (
    .I1(RESET),
    .I0(__1653__),
    .O(__3870__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8033__ (
    .I1(RESET),
    .I0(__682__),
    .O(__3871__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8034__ (
    .I1(RESET),
    .I0(__468__),
    .O(__3872__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8035__ (
    .I1(RESET),
    .I0(__258__),
    .O(__3873__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8036__ (
    .I1(RESET),
    .I0(__289__),
    .O(__3874__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8037__ (
    .I1(RESET),
    .I0(__872__),
    .O(__3875__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8038__ (
    .I1(RESET),
    .I0(__240__),
    .O(__3876__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8039__ (
    .I1(RESET),
    .I0(__1062__),
    .O(__3877__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8040__ (
    .I1(RESET),
    .I0(__1538__),
    .O(__3878__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __8041__ (
    .I5(TM0),
    .I4(__1074__),
    .I3(__1042__),
    .I2(__1010__),
    .I1(__1106__),
    .I0(__941__),
    .O(__3879__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __8042__ (
    .I5(TM0),
    .I4(__882__),
    .I3(__850__),
    .I2(__818__),
    .I1(__914__),
    .I0(__786__),
    .O(__3880__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __8043__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__3880__),
    .I0(__3879__),
    .O(__3881__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8044__ (
    .I1(TM0),
    .I0(__237__),
    .O(__3882__)
  );
  LUT6 #(
    .INIT(64'h6996966996696996)
  ) __8045__ (
    .I5(TM1),
    .I4(__142__),
    .I3(__187__),
    .I2(__173__),
    .I1(__206__),
    .I0(__3882__),
    .O(__3883__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8046__ (
    .I1(RESET),
    .I0(__823__),
    .O(__3884__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8047__ (
    .I1(RESET),
    .I0(__1245__),
    .O(__3885__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __8048__ (
    .I2(TM0),
    .I1(__1697__),
    .I0(DATA_0_1),
    .O(__3886__)
  );
  LUT6 #(
    .INIT(64'hff88f0f000000000)
  ) __8049__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__3741__),
    .I2(__3886__),
    .I1(TM0),
    .I0(__1566__),
    .O(__3887__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8050__ (
    .I1(RESET),
    .I0(__1458__),
    .O(__3888__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8051__ (
    .I1(RESET),
    .I0(__463__),
    .O(__3889__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8052__ (
    .I1(RESET),
    .I0(__1398__),
    .O(__3890__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8053__ (
    .I1(RESET),
    .I0(__291__),
    .O(__3891__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __8054__ (
    .I2(RESET),
    .I1(__914__),
    .I0(__940__),
    .O(__3892__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8055__ (
    .I1(TM0),
    .I0(__71__),
    .O(__3893__)
  );
  LUT5 #(
    .INIT(32'h41141441)
  ) __8056__ (
    .I4(__142__),
    .I3(__187__),
    .I2(__173__),
    .I1(__206__),
    .I0(TM0),
    .O(__3894__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __8057__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__3894__),
    .I2(__3882__),
    .I1(__2191__),
    .I0(__3893__),
    .O(__3895__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __8058__ (
    .I2(RESET),
    .I1(__1721__),
    .I0(__1669__),
    .O(__3896__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8059__ (
    .I1(RESET),
    .I0(__875__),
    .O(__3897__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __8060__ (
    .I2(RESET),
    .I1(__1531__),
    .I0(__1475__),
    .O(__3898__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8061__ (
    .I1(RESET),
    .I0(__1402__),
    .O(__3899__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8062__ (
    .I1(RESET),
    .I0(__1433__),
    .O(__3900__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8063__ (
    .I1(TM0),
    .I0(__570__),
    .O(__3901__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8064__ (
    .I1(TM0),
    .I0(__389__),
    .O(__3902__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __8065__ (
    .I5(TM1),
    .I4(__485__),
    .I3(__453__),
    .I2(__421__),
    .I1(__517__),
    .I0(TM0),
    .O(__3903__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __8066__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__3903__),
    .I2(__3902__),
    .I1(__2178__),
    .I0(__3901__),
    .O(__3904__)
  );
  LUT6 #(
    .INIT(64'h6996966996696996)
  ) __8067__ (
    .I5(TM1),
    .I4(__211__),
    .I3(__243__),
    .I2(__276__),
    .I1(__177__),
    .I0(__2640__),
    .O(__3905__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8068__ (
    .I1(RESET),
    .I0(__694__),
    .O(__3906__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __8069__ (
    .I2(RESET),
    .I1(__1668__),
    .I0(__1722__),
    .O(__3907__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __8070__ (
    .I2(RESET),
    .I1(__1532__),
    .I0(__1474__),
    .O(__3908__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8071__ (
    .I1(RESET),
    .I0(__772__),
    .O(__3909__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8072__ (
    .I1(RESET),
    .I0(__260__),
    .O(__3910__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8073__ (
    .I1(RESET),
    .I0(__1432__),
    .O(__3911__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8074__ (
    .I1(RESET),
    .I0(__1026__),
    .O(__3912__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __8075__ (
    .I2(RESET),
    .I1(__70__),
    .I0(__175__),
    .O(__3913__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8076__ (
    .I1(RESET),
    .I0(__1270__),
    .O(__3914__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8077__ (
    .I1(RESET),
    .I0(__608__),
    .O(__3915__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __8078__ (
    .I5(TM0),
    .I4(__507__),
    .I3(__475__),
    .I2(__443__),
    .I1(__539__),
    .I0(__356__),
    .O(__3916__)
  );
  LUT6 #(
    .INIT(64'hff880f0f00000000)
  ) __8079__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__1741__),
    .I2(__3916__),
    .I1(TM0),
    .I0(__86__),
    .O(__3917__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8080__ (
    .I1(RESET),
    .I0(__789__),
    .O(__3918__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8081__ (
    .I1(RESET),
    .I0(__443__),
    .O(__3919__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8082__ (
    .I1(TM0),
    .I0(__1531__),
    .O(__3920__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8083__ (
    .I1(TM0),
    .I0(__1348__),
    .O(__3921__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __8084__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__3921__),
    .I2(__1951__),
    .I1(__2107__),
    .I0(__3920__),
    .O(__3922__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8085__ (
    .I1(RESET),
    .I0(__1345__),
    .O(__3923__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __8086__ (
    .I2(RESET),
    .I1(__374__),
    .I0(__328__),
    .O(__3924__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __8087__ (
    .I2(RESET),
    .I1(__1280__),
    .I0(__1342__),
    .O(__3925__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8088__ (
    .I1(RESET),
    .I0(__450__),
    .O(__3926__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __8089__ (
    .I2(RESET),
    .I1(__1520__),
    .I0(__1486__),
    .O(__3927__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __8090__ (
    .I5(TM0),
    .I4(__881__),
    .I3(__849__),
    .I2(__817__),
    .I1(__913__),
    .I0(__750__),
    .O(__3928__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __8091__ (
    .I5(TM0),
    .I4(__625__),
    .I3(__689__),
    .I2(__657__),
    .I1(__721__),
    .I0(__593__),
    .O(__3929__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __8092__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__3929__),
    .I0(__3928__),
    .O(__3930__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8093__ (
    .I1(RESET),
    .I0(__1269__),
    .O(__3931__)
  );
  LUT6 #(
    .INIT(64'h6996966996696996)
  ) __8094__ (
    .I5(TM1),
    .I4(__139__),
    .I3(__170__),
    .I2(__203__),
    .I1(__106__),
    .I0(__3204__),
    .O(__3932__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8095__ (
    .I1(RESET),
    .I0(__1__),
    .O(__3933__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8096__ (
    .I1(RESET),
    .I0(__421__),
    .O(__3934__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __8097__ (
    .I5(TM0),
    .I4(__882__),
    .I3(__850__),
    .I2(__818__),
    .I1(__914__),
    .I0(__749__),
    .O(__3935__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __8098__ (
    .I5(TM0),
    .I4(__690__),
    .I3(__658__),
    .I2(__626__),
    .I1(__722__),
    .I0(__594__),
    .O(__3936__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __8099__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__3936__),
    .I0(__3935__),
    .O(__3937__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __8100__ (
    .I2(RESET),
    .I1(__519__),
    .I0(__567__),
    .O(__3938__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8101__ (
    .I1(RESET),
    .I0(__140__),
    .O(__3939__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8102__ (
    .I1(RESET),
    .I0(__1461__),
    .O(__3940__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8103__ (
    .I1(RESET),
    .I0(__865__),
    .O(__3941__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8104__ (
    .I1(RESET),
    .I0(__678__),
    .O(__3942__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8105__ (
    .I1(TM0),
    .I0(__956__),
    .O(__3943__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8106__ (
    .I1(TM0),
    .I0(__771__),
    .O(__3944__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __8107__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__3944__),
    .I2(__2400__),
    .I1(__2028__),
    .I0(__3943__),
    .O(__3945__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8108__ (
    .I1(RESET),
    .I0(__67__),
    .O(__3946__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8109__ (
    .I1(RESET),
    .I0(__79__),
    .O(__3947__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8110__ (
    .I1(RESET),
    .I0(__415__),
    .O(__3948__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8111__ (
    .I1(RESET),
    .I0(__1659__),
    .O(__3949__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8112__ (
    .I1(RESET),
    .I0(__1040__),
    .O(__3950__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __8113__ (
    .I5(TM0),
    .I4(__1271__),
    .I3(__1239__),
    .I2(__1207__),
    .I1(__1303__),
    .I0(__1128__),
    .O(__3951__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __8114__ (
    .I5(TM0),
    .I4(__1079__),
    .I3(__1047__),
    .I2(__1015__),
    .I1(__1111__),
    .I0(__983__),
    .O(__3952__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __8115__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__3952__),
    .I0(__3951__),
    .O(__3953__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8116__ (
    .I1(RESET),
    .I0(__693__),
    .O(__3954__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8117__ (
    .I1(RESET),
    .I0(__637__),
    .O(__3955__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8118__ (
    .I1(RESET),
    .I0(__1198__),
    .O(__3956__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8119__ (
    .I1(RESET),
    .I0(__1249__),
    .O(__3957__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __8120__ (
    .I2(RESET),
    .I1(__334__),
    .I0(__368__),
    .O(__3958__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __8121__ (
    .I2(RESET),
    .I1(__957__),
    .I0(__897__),
    .O(__3959__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __8122__ (
    .I5(TM0),
    .I4(__1468__),
    .I3(__1436__),
    .I2(__1404__),
    .I1(__1500__),
    .I0(__1372__),
    .O(__3960__)
  );
  LUT6 #(
    .INIT(64'h00fff8f800000000)
  ) __8123__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__3960__),
    .I2(__3588__),
    .I1(TM0),
    .I0(__1507__),
    .O(__3961__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8124__ (
    .I1(RESET),
    .I0(__861__),
    .O(__3962__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8125__ (
    .I1(RESET),
    .I0(__491__),
    .O(__3963__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8126__ (
    .I1(RESET),
    .I0(__1586__),
    .O(__3964__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8127__ (
    .I1(RESET),
    .I0(__835__),
    .O(__3965__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8128__ (
    .I1(RESET),
    .I0(__811__),
    .O(__3966__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8129__ (
    .I1(RESET),
    .I0(__319__),
    .O(__3967__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8130__ (
    .I1(TM0),
    .I0(__957__),
    .O(__3968__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8131__ (
    .I1(TM0),
    .I0(__770__),
    .O(__3969__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __8132__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__3969__),
    .I2(__2854__),
    .I1(__3794__),
    .I0(__3968__),
    .O(__3970__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8133__ (
    .I1(RESET),
    .I0(__21__),
    .O(__3971__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8134__ (
    .I1(RESET),
    .I0(__84__),
    .O(__3972__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8135__ (
    .I1(RESET),
    .I0(__30__),
    .O(__3973__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8136__ (
    .I1(RESET),
    .I0(__1164__),
    .O(__3974__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __8137__ (
    .I5(TM0),
    .I4(__635__),
    .I3(__699__),
    .I2(__667__),
    .I1(__731__),
    .I0(__548__),
    .O(__3975__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __8138__ (
    .I5(TM0),
    .I4(__507__),
    .I3(__475__),
    .I2(__443__),
    .I1(__539__),
    .I0(__411__),
    .O(__3976__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __8139__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__3976__),
    .I0(__3975__),
    .O(__3977__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8140__ (
    .I1(RESET),
    .I0(__457__),
    .O(__3978__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8141__ (
    .I1(RESET),
    .I0(__198__),
    .O(__3979__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8142__ (
    .I1(RESET),
    .I0(__92__),
    .O(__3980__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __8143__ (
    .I2(RESET),
    .I1(__1128__),
    .I0(__1110__),
    .O(__3981__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8144__ (
    .I1(RESET),
    .I0(__8__),
    .O(__3982__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8145__ (
    .I1(RESET),
    .I0(__1548__),
    .O(__3983__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __8146__ (
    .I5(TM0),
    .I4(__198__),
    .I3(__230__),
    .I2(__264__),
    .I1(__164__),
    .I0(__290__),
    .O(__3984__)
  );
  LUT6 #(
    .INIT(64'h00fff8f800000000)
  ) __8147__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__3984__),
    .I2(__1924__),
    .I1(TM0),
    .I0(__162__),
    .O(__3985__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8148__ (
    .I1(RESET),
    .I0(__692__),
    .O(__3986__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8149__ (
    .I1(RESET),
    .I0(__890__),
    .O(__3987__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8150__ (
    .I1(RESET),
    .I0(__1413__),
    .O(__3988__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8151__ (
    .I1(RESET),
    .I0(__481__),
    .O(__3989__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8152__ (
    .I1(RESET),
    .I0(__1465__),
    .O(__3990__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8153__ (
    .I1(RESET),
    .I0(__972__),
    .O(__3991__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8154__ (
    .I1(RESET),
    .I0(__500__),
    .O(__3992__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8155__ (
    .I1(RESET),
    .I0(__1378__),
    .O(__3993__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8156__ (
    .I1(RESET),
    .I0(__1240__),
    .O(__3994__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8157__ (
    .I1(RESET),
    .I0(__1163__),
    .O(__3995__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8158__ (
    .I1(RESET),
    .I0(__403__),
    .O(__3996__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8159__ (
    .I1(RESET),
    .I0(__211__),
    .O(__3997__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8160__ (
    .I1(RESET),
    .I0(__1429__),
    .O(__3998__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __8161__ (
    .I2(RESET),
    .I1(__956__),
    .I0(__898__),
    .O(__3999__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __8162__ (
    .I5(TM0),
    .I4(__215__),
    .I3(__149__),
    .I2(__181__),
    .I1(__247__),
    .I0(__280__),
    .O(__4000__)
  );
  LUT6 #(
    .INIT(64'h00fff8f800000000)
  ) __8163__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__4000__),
    .I2(__2289__),
    .I1(TM0),
    .I0(__155__),
    .O(__4001__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8164__ (
    .I1(RESET),
    .I0(__1604__),
    .O(__4002__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8165__ (
    .I1(RESET),
    .I0(__392__),
    .O(__4003__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __8166__ (
    .I2(RESET),
    .I1(__144__),
    .I0(__149__),
    .O(__4004__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8167__ (
    .I1(RESET),
    .I0(__601__),
    .O(__4005__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8168__ (
    .I1(RESET),
    .I0(__1243__),
    .O(__4006__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8169__ (
    .I1(RESET),
    .I0(__208__),
    .O(__4007__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8170__ (
    .I1(RESET),
    .I0(__1039__),
    .O(__4008__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __8171__ (
    .I2(RESET),
    .I1(__754__),
    .I0(__716__),
    .O(__4009__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8172__ (
    .I1(RESET),
    .I0(__24__),
    .O(__4010__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8173__ (
    .I1(RESET),
    .I0(__593__),
    .O(__4011__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8174__ (
    .I1(RESET),
    .I0(__215__),
    .O(__4012__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8175__ (
    .I1(RESET),
    .I0(__1376__),
    .O(__4013__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8176__ (
    .I1(RESET),
    .I0(__1354__),
    .O(__4014__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __8177__ (
    .I2(RESET),
    .I1(__1321__),
    .I0(__1301__),
    .O(__4015__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8178__ (
    .I1(RESET),
    .I0(__426__),
    .O(__4016__)
  );
  LUT6 #(
    .INIT(64'h6996966996696996)
  ) __8179__ (
    .I5(TM1),
    .I4(__192__),
    .I3(__174__),
    .I2(__207__),
    .I1(__188__),
    .I0(__2917__),
    .O(__4017__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8180__ (
    .I1(RESET),
    .I0(__829__),
    .O(__4018__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8181__ (
    .I1(TM0),
    .I0(__381__),
    .O(__4019__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8182__ (
    .I1(TM0),
    .I0(__130__),
    .O(__4020__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __8183__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__4020__),
    .I2(__2258__),
    .I1(__2929__),
    .I0(__4019__),
    .O(__4021__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __8184__ (
    .I5(TM0),
    .I4(__1467__),
    .I3(__1435__),
    .I2(__1403__),
    .I1(__1499__),
    .I0(__1316__),
    .O(__4022__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __8185__ (
    .I5(TM0),
    .I4(__1275__),
    .I3(__1243__),
    .I2(__1211__),
    .I1(__1307__),
    .I0(__1179__),
    .O(__4023__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __8186__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__4023__),
    .I0(__4022__),
    .O(__4024__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8187__ (
    .I1(RESET),
    .I0(__1181__),
    .O(__4025__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8188__ (
    .I1(RESET),
    .I0(__1609__),
    .O(__4026__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8189__ (
    .I1(RESET),
    .I0(__814__),
    .O(__4027__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8190__ (
    .I1(RESET),
    .I0(__277__),
    .O(__4028__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8191__ (
    .I1(RESET),
    .I0(__172__),
    .O(__4029__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __8192__ (
    .I2(TM0),
    .I1(__1700__),
    .I0(DATA_0_4),
    .O(__4030__)
  );
  LUT6 #(
    .INIT(64'hff88f0f000000000)
  ) __8193__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__2829__),
    .I2(__4030__),
    .I1(TM0),
    .I0(__1563__),
    .O(__4031__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8194__ (
    .I1(RESET),
    .I0(__1587__),
    .O(__4032__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __8195__ (
    .I5(TM0),
    .I4(__1456__),
    .I3(__1424__),
    .I2(__1392__),
    .I1(__1488__),
    .I0(__1360__),
    .O(__4033__)
  );
  LUT6 #(
    .INIT(64'h00fff8f800000000)
  ) __8196__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__4033__),
    .I2(__2375__),
    .I1(TM0),
    .I0(__1519__),
    .O(__4034__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8197__ (
    .I1(RESET),
    .I0(__1360__),
    .O(__4035__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8198__ (
    .I1(RESET),
    .I0(__624__),
    .O(__4036__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8199__ (
    .I1(RESET),
    .I0(__977__),
    .O(__4037__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8200__ (
    .I1(TM0),
    .I0(__1525__),
    .O(__4038__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8201__ (
    .I1(TM0),
    .I0(__1354__),
    .O(__4039__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __8202__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__4039__),
    .I2(__2452__),
    .I1(__2728__),
    .I0(__4038__),
    .O(__4040__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8203__ (
    .I1(RESET),
    .I0(__1414__),
    .O(__4041__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8204__ (
    .I1(RESET),
    .I0(__1216__),
    .O(__4042__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8205__ (
    .I1(RESET),
    .I0(__782__),
    .O(__4043__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8206__ (
    .I1(RESET),
    .I0(__824__),
    .O(__4044__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8207__ (
    .I1(RESET),
    .I0(__218__),
    .O(__4045__)
  );
  LUT6 #(
    .INIT(64'h6996966996696996)
  ) __8208__ (
    .I5(TM1),
    .I4(__222__),
    .I3(__256__),
    .I2(__287__),
    .I1(__190__),
    .I0(__3269__),
    .O(__4046__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8209__ (
    .I1(RESET),
    .I0(__1230__),
    .O(__4047__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8210__ (
    .I1(RESET),
    .I0(__311__),
    .O(__4048__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8211__ (
    .I1(RESET),
    .I0(__29__),
    .O(__4049__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8212__ (
    .I1(RESET),
    .I0(__53__),
    .O(__4050__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8213__ (
    .I1(RESET),
    .I0(__282__),
    .O(__4051__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8214__ (
    .I1(TM0),
    .I0(__369__),
    .O(__4052__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8215__ (
    .I1(TM0),
    .I0(__121__),
    .O(__4053__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __8216__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__4053__),
    .I2(__1861__),
    .I1(__3660__),
    .I0(__4052__),
    .O(__4054__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __8217__ (
    .I2(RESET),
    .I1(__1314__),
    .I0(__1308__),
    .O(__4055__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __8218__ (
    .I2(RESET),
    .I1(__955__),
    .I0(__899__),
    .O(__4056__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8219__ (
    .I1(RESET),
    .I0(__401__),
    .O(__4057__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8220__ (
    .I1(RESET),
    .I0(__1583__),
    .O(__4058__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8221__ (
    .I1(RESET),
    .I0(__179__),
    .O(__4059__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __8222__ (
    .I2(RESET),
    .I1(__357__),
    .I0(__345__),
    .O(__4060__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8223__ (
    .I1(RESET),
    .I0(__1209__),
    .O(__4061__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8224__ (
    .I1(RESET),
    .I0(__470__),
    .O(__4062__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8225__ (
    .I1(RESET),
    .I0(__857__),
    .O(__4063__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8226__ (
    .I1(RESET),
    .I0(__1254__),
    .O(__4064__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __8227__ (
    .I2(RESET),
    .I1(__937__),
    .I0(__917__),
    .O(__4065__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8228__ (
    .I1(RESET),
    .I0(__168__),
    .O(__4066__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8229__ (
    .I1(RESET),
    .I0(__27__),
    .O(__4067__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8230__ (
    .I1(RESET),
    .I0(__489__),
    .O(__4068__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8231__ (
    .I1(RESET),
    .I0(__309__),
    .O(__4069__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8232__ (
    .I1(RESET),
    .I0(__659__),
    .O(__4070__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8233__ (
    .I1(RESET),
    .I0(__635__),
    .O(__4071__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __8234__ (
    .I2(RESET),
    .I1(__1330__),
    .I0(__1292__),
    .O(__4072__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8235__ (
    .I1(RESET),
    .I0(__446__),
    .O(__4073__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8236__ (
    .I1(RESET),
    .I0(__286__),
    .O(__4074__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8237__ (
    .I1(RESET),
    .I0(__642__),
    .O(__4075__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8238__ (
    .I1(RESET),
    .I0(__479__),
    .O(__4076__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8239__ (
    .I1(RESET),
    .I0(__1082__),
    .O(__4077__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __8240__ (
    .I5(TM0),
    .I4(__702__),
    .I3(__670__),
    .I2(__638__),
    .I1(__734__),
    .I0(__545__),
    .O(__4078__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __8241__ (
    .I5(TM0),
    .I4(__510__),
    .I3(__478__),
    .I2(__446__),
    .I1(__542__),
    .I0(__414__),
    .O(__4079__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __8242__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__4079__),
    .I0(__4078__),
    .O(__4080__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8243__ (
    .I1(RESET),
    .I0(__400__),
    .O(__4081__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8244__ (
    .I1(TM0),
    .I0(__1522__),
    .O(__4082__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8245__ (
    .I1(TM0),
    .I0(__1357__),
    .O(__4083__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __8246__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__4083__),
    .I2(__2981__),
    .I1(__3311__),
    .I0(__4082__),
    .O(__4084__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8247__ (
    .I1(RESET),
    .I0(__1165__),
    .O(__4085__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8248__ (
    .I1(RESET),
    .I0(__31__),
    .O(__4086__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __8249__ (
    .I2(RESET),
    .I1(__72__),
    .I0(__187__),
    .O(__4087__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8250__ (
    .I1(RESET),
    .I0(__95__),
    .O(__4088__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8251__ (
    .I1(RESET),
    .I0(__142__),
    .O(__4089__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8252__ (
    .I1(RESET),
    .I0(__1382__),
    .O(__4090__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8253__ (
    .I1(TM0),
    .I0(__562__),
    .O(__4091__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8254__ (
    .I1(TM0),
    .I0(__397__),
    .O(__4092__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __8255__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__4092__),
    .I2(__2275__),
    .I1(__2648__),
    .I0(__4091__),
    .O(__4093__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8256__ (
    .I1(RESET),
    .I0(__1407__),
    .O(__4094__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8257__ (
    .I1(RESET),
    .I0(__1395__),
    .O(__4095__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8258__ (
    .I1(RESET),
    .I0(__787__),
    .O(__4096__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8259__ (
    .I1(TM0),
    .I0(__372__),
    .O(__4097__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8260__ (
    .I1(TM0),
    .I0(__122__),
    .O(__4098__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __8261__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__4098__),
    .I2(__2915__),
    .I1(__2716__),
    .I0(__4097__),
    .O(__4099__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8262__ (
    .I1(RESET),
    .I0(__1375__),
    .O(__4100__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8263__ (
    .I1(RESET),
    .I0(__1043__),
    .O(__4101__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8264__ (
    .I1(RESET),
    .I0(__645__),
    .O(__4102__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8265__ (
    .I1(RESET),
    .I0(__202__),
    .O(__4103__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8266__ (
    .I1(RESET),
    .I0(__679__),
    .O(__4104__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8267__ (
    .I1(RESET),
    .I0(__894__),
    .O(__4105__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8268__ (
    .I1(RESET),
    .I0(__639__),
    .O(__4106__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8269__ (
    .I1(RESET),
    .I0(__1415__),
    .O(__4107__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8270__ (
    .I1(RESET),
    .I0(__235__),
    .O(__4108__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8271__ (
    .I1(RESET),
    .I0(__983__),
    .O(__4109__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __8272__ (
    .I2(RESET),
    .I1(__553__),
    .I0(__533__),
    .O(__4110__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __8273__ (
    .I2(RESET),
    .I1(__929__),
    .I0(__925__),
    .O(__4111__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8274__ (
    .I1(TM0),
    .I0(__378__),
    .O(__4112__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8275__ (
    .I1(TM0),
    .I0(__124__),
    .O(__4113__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __8276__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__4113__),
    .I2(__3267__),
    .I1(__3903__),
    .I0(__4112__),
    .O(__4114__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8277__ (
    .I1(RESET),
    .I0(__295__),
    .O(__4115__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8278__ (
    .I1(TM0),
    .I0(__955__),
    .O(__4116__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8279__ (
    .I1(TM0),
    .I0(__772__),
    .O(__4117__)
  );
  LUT6 #(
    .INIT(64'h4114144114414114)
  ) __8280__ (
    .I5(TM1),
    .I4(__868__),
    .I3(__836__),
    .I2(__804__),
    .I1(__900__),
    .I0(TM0),
    .O(__4118__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __8281__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__4118__),
    .I2(__4117__),
    .I1(__3833__),
    .I0(__4116__),
    .O(__4119__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8282__ (
    .I1(RESET),
    .I0(__1237__),
    .O(__4120__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8283__ (
    .I1(RESET),
    .I0(__404__),
    .O(__4121__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8284__ (
    .I1(TM0),
    .I0(__376__),
    .O(__4122__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8285__ (
    .I1(TM0),
    .I0(__110__),
    .O(__4123__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __8286__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__4123__),
    .I2(__2763__),
    .I1(__2616__),
    .I0(__4122__),
    .O(__4124__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8287__ (
    .I1(RESET),
    .I0(__1203__),
    .O(__4125__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8288__ (
    .I1(TM0),
    .I0(__949__),
    .O(__4126__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8289__ (
    .I1(TM0),
    .I0(__778__),
    .O(__4127__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __8290__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__4127__),
    .I2(__1866__),
    .I1(__1819__),
    .I0(__4126__),
    .O(__4128__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8291__ (
    .I1(RESET),
    .I0(__448__),
    .O(__4129__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8292__ (
    .I1(RESET),
    .I0(__625__),
    .O(__4130__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __8293__ (
    .I5(TM0),
    .I4(__506__),
    .I3(__474__),
    .I2(__442__),
    .I1(__538__),
    .I0(__357__),
    .O(__4131__)
  );
  LUT6 #(
    .INIT(64'hff880f0f00000000)
  ) __8294__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__2889__),
    .I2(__4131__),
    .I1(TM0),
    .I0(__82__),
    .O(__4132__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8295__ (
    .I1(RESET),
    .I0(__1598__),
    .O(__4133__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8296__ (
    .I1(RESET),
    .I0(__1201__),
    .O(__4134__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8297__ (
    .I1(TM0),
    .I0(__1151__),
    .O(__4135__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8298__ (
    .I1(TM0),
    .I0(__960__),
    .O(__4136__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __8299__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__4136__),
    .I2(__3041__),
    .I1(__2838__),
    .I0(__4135__),
    .O(__4137__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __8300__ (
    .I2(RESET),
    .I1(__358__),
    .I0(__344__),
    .O(__4138__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8301__ (
    .I1(RESET),
    .I0(__1008__),
    .O(__4139__)
  );
  LUT3 #(
    .INIT(8'h90)
  ) __8302__ (
    .I2(RESET),
    .I1(__1120__),
    .I0(__1118__),
    .O(__4140__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8303__ (
    .I1(RESET),
    .I0(__1276__),
    .O(__4141__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __8304__ (
    .I5(TM0),
    .I4(__1463__),
    .I3(__1431__),
    .I2(__1399__),
    .I1(__1495__),
    .I0(__1367__),
    .O(__4142__)
  );
  LUT6 #(
    .INIT(64'h00fff8f800000000)
  ) __8305__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__4142__),
    .I2(__3369__),
    .I1(TM0),
    .I0(__1512__),
    .O(__4143__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8306__ (
    .I1(RESET),
    .I0(__804__),
    .O(__4144__)
  );
  LUT3 #(
    .INIT(8'hca)
  ) __8307__ (
    .I2(TM0),
    .I1(__1727__),
    .I0(DATA_0_31),
    .O(__4145__)
  );
  LUT6 #(
    .INIT(64'hff88f0f000000000)
  ) __8308__ (
    .I5(RESET),
    .I4(TM1),
    .I3(__3305__),
    .I2(__4145__),
    .I1(TM0),
    .I0(__1536__),
    .O(__4146__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __8309__ (
    .I5(TM0),
    .I4(__695__),
    .I3(__663__),
    .I2(__631__),
    .I1(__727__),
    .I0(__552__),
    .O(__4147__)
  );
  LUT6 #(
    .INIT(64'h55555555c33c3cc3)
  ) __8310__ (
    .I5(TM0),
    .I4(__503__),
    .I3(__471__),
    .I2(__439__),
    .I1(__535__),
    .I0(__407__),
    .O(__4148__)
  );
  LUT4 #(
    .INIT(16'h3500)
  ) __8311__ (
    .I3(RESET),
    .I2(TM1),
    .I1(__4148__),
    .I0(__4147__),
    .O(__4149__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8312__ (
    .I1(RESET),
    .I0(__1447__),
    .O(__4150__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8313__ (
    .I1(RESET),
    .I0(__301__),
    .O(__4151__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8314__ (
    .I1(RESET),
    .I0(__136__),
    .O(__4152__)
  );
  LUT6 #(
    .INIT(64'h4bb4b44bb44b4bb4)
  ) __8315__ (
    .I5(__180__),
    .I4(__214__),
    .I3(__246__),
    .I2(__148__),
    .I1(TM0),
    .I0(__279__),
    .O(__4153__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8316__ (
    .I1(RESET),
    .I0(__1275__),
    .O(__4154__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8317__ (
    .I1(TM0),
    .I0(__763__),
    .O(__4155__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8318__ (
    .I1(TM0),
    .I0(__580__),
    .O(__4156__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __8319__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__4156__),
    .I2(__2485__),
    .I1(__4118__),
    .I0(__4155__),
    .O(__4157__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8320__ (
    .I1(TM0),
    .I0(__1138__),
    .O(__4158__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8321__ (
    .I1(__973__),
    .I0(TM0),
    .O(__4159__)
  );
  LUT6 #(
    .INIT(64'hfff00000eeee0000)
  ) __8322__ (
    .I5(TM1),
    .I4(RESET),
    .I3(__4159__),
    .I2(__3598__),
    .I1(__2983__),
    .I0(__4158__),
    .O(__4160__)
  );
  LUT2 #(
    .INIT(4'h8)
  ) __8323__ (
    .I1(__408__),
    .I0(RESET),
    .O(__4161__)
  );
  assign CRC_OUT_9_24 = __119__;
  assign CRC_OUT_5_23 = __951__;
  assign CRC_OUT_2_14 = __1518__;
  assign CRC_OUT_7_5 = __549__;
  assign CRC_OUT_4_23 = __1143__;
  assign CRC_OUT_1_28 = __1724__;
  assign CRC_OUT_6_13 = __749__;
  assign CRC_OUT_1_19 = __1715__;
  assign CRC_OUT_9_31 = __131__;
  assign CRC_OUT_4_14 = __1134__;
  assign CRC_OUT_5_3 = __931__;
  assign CRC_OUT_2_15 = __1519__;
  assign CRC_OUT_7_15 = __559__;
  assign CRC_OUT_2_3 = __1507__;
  assign CRC_OUT_3_12 = __1324__;
  assign CRC_OUT_1_6 = __1702__;
  assign CRC_OUT_6_21 = __757__;
  assign CRC_OUT_9_25 = __133__;
  assign CRC_OUT_2_25 = __1529__;
  assign DATA_9_15 = __2129__;
  assign CRC_OUT_6_26 = __762__;
  assign DATA_9_4 = __2731__;
  assign CRC_OUT_6_3 = __739__;
  assign CRC_OUT_2_29 = __1533__;
  assign CRC_OUT_3_10 = __1322__;
  assign CRC_OUT_5_6 = __934__;
  assign CRC_OUT_2_20 = __1524__;
  assign CRC_OUT_3_27 = __1339__;
  assign CRC_OUT_6_30 = __766__;
  assign CRC_OUT_2_5 = __1509__;
  assign CRC_OUT_1_20 = __1716__;
  assign CRC_OUT_6_11 = __747__;
  assign CRC_OUT_7_29 = __573__;
  assign CRC_OUT_9_19 = __71__;
  assign CRC_OUT_1_16 = __1712__;
  assign CRC_OUT_5_1 = __929__;
  assign CRC_OUT_3_8 = __1320__;
  assign CRC_OUT_7_3 = __547__;
  assign CRC_OUT_2_8 = __1512__;
  assign DATA_9_20 = __4017__;
  assign CRC_OUT_9_11 = __154__;
  assign CRC_OUT_7_26 = __570__;
  assign CRC_OUT_1_7 = __1703__;
  assign CRC_OUT_2_17 = __1521__;
  assign CRC_OUT_2_6 = __1510__;
  assign CRC_OUT_4_11 = __1131__;
  assign CRC_OUT_9_4 = __145__;
  assign CRC_OUT_9_6 = __161__;
  assign CRC_OUT_8_3 = __355__;
  assign DATA_9_21 = __2119__;
  assign CRC_OUT_7_19 = __563__;
  assign CRC_OUT_7_22 = __566__;
  assign DATA_9_17 = __3847__;
  assign CRC_OUT_9_22 = __68__;
  assign CRC_OUT_4_31 = __1151__;
  assign CRC_OUT_2_12 = __1516__;
  assign CRC_OUT_9_21 = __69__;
  assign CRC_OUT_8_29 = __381__;
  assign CRC_OUT_9_7 = __144__;
  assign CRC_OUT_9_5 = __156__;
  assign CRC_OUT_6_7 = __743__;
  assign DATA_9_11 = __1805__;
  assign CRC_OUT_3_9 = __1321__;
  assign CRC_OUT_4_18 = __1138__;
  assign CRC_OUT_7_20 = __564__;
  assign CRC_OUT_1_11 = __1707__;
  assign CRC_OUT_3_15 = __1327__;
  assign CRC_OUT_8_31 = __383__;
  assign CRC_OUT_5_13 = __941__;
  assign CRC_OUT_1_31 = __1727__;
  assign CRC_OUT_6_28 = __764__;
  assign CRC_OUT_5_19 = __947__;
  assign CRC_OUT_3_3 = __1315__;
  assign CRC_OUT_6_0 = __736__;
  assign DATA_9_8 = __2750__;
  assign CRC_OUT_9_29 = __113__;
  assign CRC_OUT_8_21 = __373__;
  assign DATA_9_0 = __3068__;
  assign CRC_OUT_9_26 = __114__;
  assign CRC_OUT_1_4 = __1700__;
  assign CRC_OUT_1_22 = __1718__;
  assign CRC_OUT_4_24 = __1144__;
  assign CRC_OUT_6_6 = __742__;
  assign CRC_OUT_4_13 = __1133__;
  assign CRC_OUT_3_16 = __1328__;
  assign CRC_OUT_4_10 = __1130__;
  assign CRC_OUT_5_25 = __953__;
  assign CRC_OUT_7_2 = __546__;
  assign CRC_OUT_5_12 = __940__;
  assign CRC_OUT_8_10 = __362__;
  assign CRC_OUT_4_0 = __1120__;
  assign CRC_OUT_6_16 = __752__;
  assign CRC_OUT_7_4 = __548__;
  assign CRC_OUT_5_14 = __942__;
  assign CRC_OUT_3_24 = __1336__;
  assign CRC_OUT_6_18 = __754__;
  assign CRC_OUT_9_14 = __125__;
  assign CRC_OUT_3_7 = __1319__;
  assign CRC_OUT_6_24 = __760__;
  assign CRC_OUT_5_5 = __933__;
  assign CRC_OUT_6_19 = __755__;
  assign CRC_OUT_3_11 = __1323__;
  assign CRC_OUT_8_11 = __363__;
  assign CRC_OUT_6_20 = __756__;
  assign CRC_OUT_5_24 = __952__;
  assign CRC_OUT_4_2 = __1122__;
  assign CRC_OUT_3_6 = __1318__;
  assign CRC_OUT_4_27 = __1147__;
  assign CRC_OUT_6_9 = __745__;
  assign CRC_OUT_2_2 = __1506__;
  assign CRC_OUT_5_4 = __932__;
  assign CRC_OUT_7_27 = __571__;
  assign CRC_OUT_2_26 = __1530__;
  assign CRC_OUT_5_7 = __935__;
  assign CRC_OUT_2_27 = __1531__;
  assign CRC_OUT_5_20 = __948__;
  assign CRC_OUT_4_17 = __1137__;
  assign CRC_OUT_8_6 = __358__;
  assign CRC_OUT_2_11 = __1515__;
  assign CRC_OUT_4_3 = __1123__;
  assign CRC_OUT_8_26 = __378__;
  assign CRC_OUT_1_5 = __1701__;
  assign CRC_OUT_4_4 = __1124__;
  assign CRC_OUT_5_0 = __928__;
  assign CRC_OUT_4_22 = __1142__;
  assign CRC_OUT_9_27 = __118__;
  assign CRC_OUT_9_8 = __155__;
  assign DATA_9_13 = __2385__;
  assign DATA_9_7 = __3809__;
  assign CRC_OUT_3_14 = __1326__;
  assign CRC_OUT_3_2 = __1314__;
  assign CRC_OUT_3_5 = __1317__;
  assign CRC_OUT_3_20 = __1332__;
  assign CRC_OUT_8_2 = __354__;
  assign CRC_OUT_7_17 = __561__;
  assign CRC_OUT_2_24 = __1528__;
  assign CRC_OUT_8_25 = __377__;
  assign DATA_9_1 = __2604__;
  assign CRC_OUT_2_16 = __1520__;
  assign CRC_OUT_5_29 = __957__;
  assign DATA_9_29 = __2526__;
  assign CRC_OUT_2_22 = __1526__;
  assign CRC_OUT_4_19 = __1139__;
  assign DATA_9_27 = __3905__;
  assign CRC_OUT_1_15 = __1711__;
  assign CRC_OUT_2_4 = __1508__;
  assign CRC_OUT_9_28 = __132__;
  assign CRC_OUT_4_5 = __1125__;
  assign CRC_OUT_2_7 = __1511__;
  assign DATA_9_30 = __2520__;
  assign CRC_OUT_5_30 = __958__;
  assign CRC_OUT_2_23 = __1527__;
  assign CRC_OUT_6_31 = __767__;
  assign CRC_OUT_1_17 = __1713__;
  assign CRC_OUT_4_7 = __1127__;
  assign CRC_OUT_4_25 = __1145__;
  assign CRC_OUT_6_14 = __750__;
  assign CRC_OUT_3_18 = __1330__;
  assign CRC_OUT_5_26 = __954__;
  assign CRC_OUT_5_28 = __956__;
  assign CRC_OUT_1_27 = __1723__;
  assign CRC_OUT_7_12 = __556__;
  assign CRC_OUT_3_28 = __1340__;
  assign CRC_OUT_9_16 = __74__;
  assign CRC_OUT_4_12 = __1132__;
  assign CRC_OUT_7_7 = __551__;
  assign CRC_OUT_4_15 = __1135__;
  assign CRC_OUT_6_10 = __746__;
  assign DATA_9_25 = __1893__;
  assign CRC_OUT_7_8 = __552__;
  assign CRC_OUT_9_30 = __117__;
  assign CRC_OUT_8_1 = __353__;
  assign CRC_OUT_8_16 = __368__;
  assign CRC_OUT_3_31 = __1343__;
  assign CRC_OUT_1_3 = __1699__;
  assign CRC_OUT_2_30 = __1534__;
  assign CRC_OUT_4_8 = __1128__;
  assign CRC_OUT_1_23 = __1719__;
  assign CRC_OUT_8_30 = __382__;
  assign CRC_OUT_6_1 = __737__;
  assign CRC_OUT_8_7 = __359__;
  assign CRC_OUT_8_8 = __360__;
  assign CRC_OUT_9_13 = __158__;
  assign CRC_OUT_5_11 = __939__;
  assign CRC_OUT_1_0 = __1696__;
  assign CRC_OUT_3_29 = __1341__;
  assign CRC_OUT_7_9 = __553__;
  assign CRC_OUT_5_8 = __936__;
  assign CRC_OUT_5_21 = __949__;
  assign CRC_OUT_9_2 = __157__;
  assign CRC_OUT_2_0 = __1504__;
  assign DATA_9_26 = __4046__;
  assign CRC_OUT_3_17 = __1329__;
  assign CRC_OUT_8_15 = __367__;
  assign DATA_9_2 = __3322__;
  assign CRC_OUT_2_28 = __1532__;
  assign DATA_9_14 = __3221__;
  assign CRC_OUT_9_17 = __73__;
  assign CRC_OUT_9_3 = __162__;
  assign DATA_9_9 = __3716__;
  assign CRC_OUT_8_17 = __369__;
  assign DATA_9_19 = __3883__;
  assign DATA_9_10 = __2111__;
  assign CRC_OUT_7_13 = __557__;
  assign CRC_OUT_7_23 = __567__;
  assign CRC_OUT_2_1 = __1505__;
  assign CRC_OUT_1_26 = __1722__;
  assign CRC_OUT_9_9 = __160__;
  assign CRC_OUT_8_14 = __366__;
  assign CRC_OUT_1_14 = __1710__;
  assign CRC_OUT_7_16 = __560__;
  assign CRC_OUT_3_23 = __1335__;
  assign CRC_OUT_8_13 = __365__;
  assign CRC_OUT_9_23 = __115__;
  assign CRC_OUT_8_19 = __371__;
  assign DATA_9_23 = __2577__;
  assign CRC_OUT_8_28 = __380__;
  assign CRC_OUT_9_18 = __72__;
  assign CRC_OUT_1_21 = __1717__;
  assign CRC_OUT_4_1 = __1121__;
  assign CRC_OUT_1_24 = __1720__;
  assign CRC_OUT_2_21 = __1525__;
  assign CRC_OUT_4_26 = __1146__;
  assign CRC_OUT_6_2 = __738__;
  assign CRC_OUT_7_25 = __569__;
  assign CRC_OUT_3_25 = __1337__;
  assign CRC_OUT_9_12 = __159__;
  assign CRC_OUT_9_15 = __75__;
  assign DATA_9_22 = __2305__;
  assign CRC_OUT_1_1 = __1697__;
  assign DATA_9_5 = __4153__;
  assign CRC_OUT_8_0 = __352__;
  assign DATA_9_31 = __3237__;
  assign CRC_OUT_7_21 = __565__;
  assign DATA_9_16 = __3932__;
  assign CRC_OUT_2_13 = __1517__;
  assign CRC_OUT_9_10 = __143__;
  assign DATA_9_28 = __3634__;
  assign CRC_OUT_8_4 = __356__;
  assign CRC_OUT_4_29 = __1149__;
  assign CRC_OUT_6_8 = __744__;
  assign CRC_OUT_3_13 = __1325__;
  assign CRC_OUT_3_30 = __1342__;
  assign CRC_OUT_1_30 = __1726__;
  assign CRC_OUT_8_5 = __357__;
  assign CRC_OUT_6_15 = __751__;
  assign CRC_OUT_6_5 = __741__;
  assign CRC_OUT_1_10 = __1706__;
  assign CRC_OUT_7_18 = __562__;
  assign CRC_OUT_4_9 = __1129__;
  assign CRC_OUT_1_13 = __1709__;
  assign CRC_OUT_8_27 = __379__;
  assign CRC_OUT_5_2 = __930__;
  assign CRC_OUT_8_12 = __364__;
  assign CRC_OUT_8_22 = __374__;
  assign CRC_OUT_7_11 = __555__;
  assign CRC_OUT_7_10 = __554__;
  assign CRC_OUT_6_25 = __761__;
  assign CRC_OUT_6_23 = __759__;
  assign CRC_OUT_1_9 = __1705__;
  assign CRC_OUT_7_0 = __544__;
  assign CRC_OUT_7_1 = __545__;
  assign CRC_OUT_4_21 = __1141__;
  assign CRC_OUT_9_0 = __146__;
  assign CRC_OUT_1_2 = __1698__;
  assign CRC_OUT_6_17 = __753__;
  assign CRC_OUT_5_10 = __938__;
  assign CRC_OUT_8_9 = __361__;
  assign CRC_OUT_7_24 = __568__;
  assign CRC_OUT_5_22 = __950__;
  assign CRC_OUT_7_14 = __558__;
  assign DATA_9_18 = __3610__;
  assign CRC_OUT_7_28 = __572__;
  assign CRC_OUT_3_22 = __1334__;
  assign CRC_OUT_6_29 = __765__;
  assign CRC_OUT_8_20 = __372__;
  assign CRC_OUT_6_22 = __758__;
  assign CRC_OUT_5_17 = __945__;
  assign CRC_OUT_3_1 = __1313__;
  assign CRC_OUT_3_19 = __1331__;
  assign CRC_OUT_5_9 = __937__;
  assign CRC_OUT_3_4 = __1316__;
  assign CRC_OUT_1_18 = __1714__;
  assign CRC_OUT_5_16 = __944__;
  assign CRC_OUT_6_4 = __740__;
  assign CRC_OUT_8_24 = __376__;
  assign CRC_OUT_2_10 = __1514__;
  assign DATA_9_24 = __2105__;
  assign CRC_OUT_8_23 = __375__;
  assign CRC_OUT_8_18 = __370__;
  assign CRC_OUT_1_8 = __1704__;
  assign CRC_OUT_2_31 = __1535__;
  assign CRC_OUT_2_19 = __1523__;
  assign CRC_OUT_4_16 = __1136__;
  assign CRC_OUT_7_31 = __575__;
  assign CRC_OUT_2_18 = __1522__;
  assign CRC_OUT_4_6 = __1126__;
  assign CRC_OUT_2_9 = __1513__;
  assign CRC_OUT_5_31 = __959__;
  assign CRC_OUT_5_18 = __946__;
  assign CRC_OUT_6_27 = __763__;
  assign CRC_OUT_3_21 = __1333__;
  assign CRC_OUT_1_25 = __1721__;
  assign CRC_OUT_4_30 = __1150__;
  assign DATA_9_3 = __2346__;
  assign CRC_OUT_1_12 = __1708__;
  assign CRC_OUT_7_6 = __550__;
  assign CRC_OUT_9_1 = __150__;
  assign CRC_OUT_5_15 = __943__;
  assign CRC_OUT_5_27 = __955__;
  assign CRC_OUT_7_30 = __574__;
  assign CRC_OUT_3_26 = __1338__;
  assign CRC_OUT_3_0 = __1312__;
  assign CRC_OUT_1_29 = __1725__;
  assign CRC_OUT_9_20 = __70__;
  assign DATA_9_12 = __3224__;
  assign CRC_OUT_6_12 = __748__;
  assign DATA_9_6 = __3518__;
  assign CRC_OUT_4_20 = __1140__;
  assign CRC_OUT_4_28 = __1148__;
endmodule
