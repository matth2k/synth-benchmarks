// IWLS benchmark module "CM85" printed on Wed May 29 16:31:28 2002
module CM85(a, b, c, d, e, f, g, h, i, j, k, l, m, n);
input
  a,
  b,
  c,
  d,
  e,
  f,
  g,
  h,
  i,
  j,
  k;
output
  l,
  m,
  n;
wire
  d0,
  e0,
  q0,
  f0,
  g0,
  h0,
  \[0] ,
  t0,
  i0,
  \[1] ,
  u0,
  j0,
  \[2] ,
  u,
  v,
  w,
  \xx ,
  v0,
  k0,
  w0,
  l0,
  a0,
  m0,
  n0;
assign
  d0 = f | ~g,
  e0 = ~f | g,
  q0 = (~i & ~h) | (i & h),
  f0 = ~a0 | ~b,
  g0 = (~g & f) | (g & ~f),
  h0 = ~g0 & ~f0,
  \[0]  = (~t0 & ~v0) | ~n0,
  t0 = j | ~k,
  i0 = (~f0 & ~e0) | ~v,
  \[1]  = ~w0 & ~v0,
  l = \[0] ,
  m = \[1] ,
  n = \[2] ,
  u0 = ~j | k,
  j0 = (~d0 & ~f0) | ~\xx ,
  \[2]  = (~u0 & ~v0) | ~l0,
  u = d & ~e,
  v = (~c & ~u) | (~c & ~b),
  w = ~d & e,
  \xx  = (~a & ~w) | (~a & ~b),
  v0 = ~q0 | ~h0,
  k0 = h & ~i,
  w0 = (~k & j) | (k & ~j),
  l0 = (~i0 & ~k0) | (~i0 & ~h0),
  a0 = (~e & ~d) | (e & d),
  m0 = ~h & i,
  n0 = (~j0 & ~m0) | (~j0 & ~h0);
endmodule

