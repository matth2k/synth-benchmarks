// IWLS benchmark module "C880.iscas" printed on Wed May 29 16:31:25 2002
module C880 (\1GAT(0) , \8GAT(1) , \13GAT(2) , \17GAT(3) , \26GAT(4) , \29GAT(5) , \36GAT(6) , \42GAT(7) , \51GAT(8) , \55GAT(9) , \59GAT(10) , \68GAT(11) , \72GAT(12) , \73GAT(13) , \74GAT(14) , \75GAT(15) , \80GAT(16) , \85GAT(17) , \86GAT(18) , \87GAT(19) , \88GAT(20) , \89GAT(21) , \90GAT(22) , \91GAT(23) , \96GAT(24) , \101GAT(25) , \106GAT(26) , \111GAT(27) , \116GAT(28) , \121GAT(29) , \126GAT(30) , \130GAT(31) , \135GAT(32) , \138GAT(33) , \143GAT(34) , \146GAT(35) , \149GAT(36) , \152GAT(37) , \153GAT(38) , \156GAT(39) , \159GAT(40) , \165GAT(41) , \171GAT(42) , \177GAT(43) , \183GAT(44) , \189GAT(45) , \195GAT(46) , \201GAT(47) , \207GAT(48) , \210GAT(49) , \219GAT(50) , \228GAT(51) , \237GAT(52) , \246GAT(53) , \255GAT(54) , \259GAT(55) , \260GAT(56) , \261GAT(57) , \267GAT(58) , \268GAT(59) , \388GAT(133) , \389GAT(132) , \390GAT(131) , \391GAT(124) , \418GAT(168) , \419GAT(164) , \420GAT(158) , \421GAT(162) , \422GAT(161) , \423GAT(155) , \446GAT(183) , \447GAT(182) , \448GAT(179) , \449GAT(176) , \450GAT(173) , \767GAT(349) , \768GAT(334) , \850GAT(404) , \863GAT(424) , \864GAT(423) , \865GAT(422) , \866GAT(426) , \874GAT(433) , \878GAT(442) , \879GAT(441) , \880GAT(440) );
input
  \87GAT(19) ,
  \86GAT(18) ,
  \85GAT(17) ,
  \195GAT(46) ,
  \126GAT(30) ,
  \210GAT(49) ,
  \207GAT(48) ,
  \80GAT(16) ,
  \51GAT(8) ,
  \183GAT(44) ,
  \201GAT(47) ,
  \26GAT(4) ,
  \219GAT(50) ,
  \90GAT(22) ,
  \91GAT(23) ,
  \189GAT(45) ,
  \36GAT(6) ,
  \171GAT(42) ,
  \96GAT(24) ,
  \228GAT(51) ,
  \17GAT(3) ,
  \177GAT(43) ,
  \101GAT(25) ,
  \106GAT(26) ,
  \156GAT(39) ,
  \42GAT(7) ,
  \237GAT(52) ,
  \165GAT(41) ,
  \1GAT(0) ,
  \153GAT(38) ,
  \152GAT(37) ,
  \13GAT(2) ,
  \246GAT(53) ,
  \259GAT(55) ,
  \159GAT(40) ,
  \130GAT(31) ,
  \255GAT(54) ,
  \138GAT(33) ,
  \267GAT(58) ,
  \135GAT(32) ,
  \121GAT(29) ,
  \59GAT(10) ,
  \116GAT(28) ,
  \268GAT(59) ,
  \143GAT(34) ,
  \149GAT(36) ,
  \261GAT(57) ,
  \260GAT(56) ,
  \29GAT(5) ,
  \111GAT(27) ,
  \146GAT(35) ,
  \68GAT(11) ,
  \73GAT(13) ,
  \72GAT(12) ,
  \8GAT(1) ,
  \55GAT(9) ,
  \75GAT(15) ,
  \74GAT(14) ,
  \88GAT(20) ,
  \89GAT(21) ;
output
  \865GAT(422) ,
  \420GAT(158) ,
  \419GAT(164) ,
  \418GAT(168) ,
  \864GAT(423) ,
  \421GAT(162) ,
  \874GAT(433) ,
  \866GAT(426) ,
  \448GAT(179) ,
  \850GAT(404) ,
  \388GAT(133) ,
  \422GAT(161) ,
  \423GAT(155) ,
  \449GAT(176) ,
  \389GAT(132) ,
  \768GAT(334) ,
  \879GAT(441) ,
  \880GAT(440) ,
  \863GAT(424) ,
  \447GAT(182) ,
  \767GAT(349) ,
  \391GAT(124) ,
  \878GAT(442) ,
  \446GAT(183) ,
  \450GAT(173) ,
  \390GAT(131) ;
wire
  \569GAT(247) ,
  \425GAT(172) ,
  \792GAT(363) ,
  \815GAT(388) ,
  \526GAT(212) ,
  \734GAT(287) ,
  \269GAT(112) ,
  \503GAT(203) ,
  \782GAT(353) ,
  \499GAT(225) ,
  \350GAT(126) ,
  \696GAT(305) ,
  \765GAT(346) ,
  \322GAT(105) ,
  \405GAT(152) ,
  \506GAT(232) ,
  \773GAT(351) ,
  \844GAT(408) ,
  \478GAT(189) ,
  \327GAT(68) ,
  \326GAT(69) ,
  \632GAT(275) ,
  \628GAT(276) ,
  \687GAT(304) ,
  \631GAT(264) ,
  \353GAT(130) ,
  \336GAT(77) ,
  \489GAT(185) ,
  \527GAT(211) ,
  \796GAT(373) ,
  \855GAT(418) ,
  \477GAT(196) ,
  \498GAT(226) ,
  \338GAT(76) ,
  \347GAT(138) ,
  \329GAT(66) ,
  \328GAT(67) ,
  \686GAT(308) ,
  \417GAT(142) ,
  \736GAT(333) ,
  \747GAT(341) ,
  \757GAT(317) ,
  \360GAT(120) ,
  \460GAT(199) ,
  \660GAT(315) ,
  \867GAT(432) ,
  \825GAT(385) ,
  \843GAT(409) ,
  \661GAT(293) ,
  \640GAT(263) ,
  \346GAT(140) ,
  \733GAT(288) ,
  \379GAT(116) ,
  \586GAT(255) ,
  \834GAT(397) ,
  \406GAT(153) ,
  \751GAT(328) ,
  \410GAT(160) ,
  \528GAT(210) ,
  \332GAT(85) ,
  \333GAT(84) ,
  \340GAT(73) ,
  \593GAT(284) ,
  \369GAT(113) ,
  \399GAT(166) ,
  \542GAT(237) ,
  \443GAT(180) ,
  \408GAT(149) ,
  \488GAT(184) ,
  \587GAT(256) ,
  \794GAT(362) ,
  \856GAT(417) ,
  \509GAT(206) ,
  \416GAT(144) ,
  \759GAT(326) ,
  \758GAT(316) ,
  \762GAT(339) ,
  \804GAT(370) ,
  \875GAT(439) ,
  \310GAT(60) ,
  \619GAT(278) ,
  \760GAT(318) ,
  \442GAT(175) ,
  \344GAT(136) ,
  \544GAT(242) ,
  \814GAT(383) ,
  \704GAT(302) ,
  \492GAT(193) ,
  \285GAT(102) ,
  \407GAT(151) ,
  \764GAT(343) ,
  \735GAT(348) ,
  \557GAT(252) ,
  \654GAT(270) ,
  \334GAT(81) ,
  \335GAT(80) ,
  \833GAT(400) ,
  \732GAT(289) ,
  \466GAT(201) ,
  \352GAT(127) ,
  \432GAT(181) ,
  \519GAT(223) ,
  \835GAT(398) ,
  \476GAT(188) ,
  \669GAT(314) ,
  \504GAT(233) ,
  \753GAT(338) ,
  \533GAT(241) ,
  \480GAT(190) ,
  \363GAT(119) ,
  \317GAT(106) ,
  \589GAT(269) ,
  \616GAT(279) ,
  \345GAT(139) ,
  \510GAT(220) ,
  \785GAT(355) ,
  \543GAT(236) ,
  \737GAT(325) ,
  \615GAT(266) ,
  \857GAT(416) ,
  \415GAT(143) ,
  \341GAT(61) ,
  \400GAT(157) ,
  \763GAT(337) ,
  \861GAT(427) ,
  \522GAT(216) ,
  \318GAT(72) ,
  \382GAT(115) ,
  \805GAT(374) ,
  \479GAT(195) ,
  \577GAT(249) ,
  \512GAT(219) ,
  \513GAT(229) ,
  \872GAT(435) ,
  \673GAT(309) ,
  \813GAT(382) ,
  \518GAT(224) ,
  \705GAT(299) ,
  \662GAT(313) ,
  \641GAT(273) ,
  \273GAT(103) ,
  \609GAT(280) ,
  \845GAT(412) ,
  \717GAT(296) ,
  \870GAT(429) ,
  \309GAT(107) ,
  \551GAT(257) ,
  \786GAT(350) ,
  \540GAT(239) ,
  \401GAT(163) ,
  \727GAT(294) ,
  \290GAT(100) ,
  \331GAT(64) ,
  \330GAT(65) ,
  \501GAT(221) ,
  \413GAT(147) ,
  \297GAT(89) ,
  \414GAT(145) ,
  \777GAT(357) ,
  \481GAT(194) ,
  \812GAT(381) ,
  \561GAT(253) ,
  \822GAT(386) ,
  \860GAT(428) ,
  \550GAT(260) ,
  \859GAT(421) ,
  \624GAT(265) ,
  \502GAT(234) ,
  \745GAT(330) ,
  \339GAT(62) ,
  \298GAT(88) ,
  \659GAT(261) ,
  \409GAT(150) ,
  \507GAT(205) ,
  \841GAT(403) ,
  \325GAT(70) ,
  \324GAT(71) ,
  \819GAT(387) ,
  \355GAT(123) ,
  \463GAT(198) ,
  \836GAT(392) ,
  \791GAT(366) ,
  \873GAT(434) ,
  \692GAT(303) ,
  \354GAT(129) ,
  \581GAT(250) ,
  \337GAT(63) ,
  \744GAT(342) ,
  \746GAT(322) ,
  \802GAT(372) ,
  \303GAT(83) ,
  \552GAT(258) ,
  \482GAT(191) ,
  \837GAT(396) ,
  \426GAT(171) ,
  \393GAT(165) ,
  \295GAT(97) ,
  \590GAT(285) ,
  \742GAT(331) ,
  \523GAT(215) ,
  \286GAT(92) ,
  \348GAT(128) ,
  \831GAT(402) ,
  \296GAT(96) ,
  \284GAT(95) ,
  \541GAT(238) ,
  \279GAT(109) ,
  \605GAT(267) ,
  \749GAT(321) ,
  \293GAT(91) ,
  \539GAT(240) ,
  \412GAT(146) ,
  \402GAT(159) ,
  \511GAT(230) ,
  \445GAT(169) ,
  \682GAT(306) ,
  \342GAT(141) ,
  \787GAT(354) ,
  \392GAT(167) ,
  \495GAT(192) ,
  \600GAT(282) ,
  \803GAT(371) ,
  \826GAT(391) ,
  \750GAT(340) ,
  \752GAT(320) ,
  \851GAT(415) ,
  \858GAT(420) ,
  \761GAT(336) ,
  \810GAT(375) ,
  \427GAT(178) ,
  \301GAT(87) ,
  \304GAT(82) ,
  \343GAT(135) ,
  \789GAT(368) ,
  \500GAT(222) ,
  \830GAT(401) ,
  \302GAT(86) ,
  \848GAT(405) ,
  \316GAT(93) ,
  \319GAT(90) ,
  \748GAT(329) ,
  \292GAT(98) ,
  \276GAT(110) ,
  \597GAT(283) ,
  \491GAT(187) ,
  \829GAT(384) ,
  \306GAT(78) ,
  \811GAT(378) ,
  \721GAT(291) ,
  \625GAT(277) ,
  \291GAT(99) ,
  \294GAT(94) ,
  \808GAT(377) ,
  \700GAT(300) ,
  \305GAT(79) ,
  \514GAT(218) ,
  \515GAT(228) ,
  \847GAT(406) ,
  \828GAT(389) ,
  \437GAT(177) ,
  \868GAT(431) ,
  \778GAT(352) ,
  \411GAT(148) ,
  \871GAT(436) ,
  \650GAT(262) ,
  \588GAT(286) ,
  \790GAT(365) ,
  \366GAT(118) ,
  \524GAT(214) ,
  \357GAT(121) ,
  \838GAT(395) ,
  \771GAT(359) ,
  \740GAT(324) ,
  \530GAT(243) ,
  \553GAT(251) ,
  \508GAT(231) ,
  \308GAT(74) ,
  \538GAT(245) ,
  \403GAT(156) ,
  \280GAT(108) ,
  \644GAT(272) ,
  \827GAT(390) ,
  \307GAT(75) ,
  \852GAT(414) ,
  \708GAT(298) ,
  \606GAT(281) ,
  \788GAT(367) ,
  \505GAT(204) ,
  \376GAT(117) ,
  \483GAT(202) ,
  \769GAT(361) ,
  \385GAT(114) ,
  \490GAT(186) ,
  \756GAT(335) ,
  \770GAT(360) ,
  \846GAT(407) ,
  \781GAT(356) ,
  \809GAT(376) ,
  \475GAT(197) ,
  \678GAT(307) ,
  \665GAT(312) ,
  \840GAT(393) ,
  \722GAT(295) ,
  \862GAT(425) ,
  \731GAT(290) ,
  \869GAT(430) ,
  \755GAT(319) ,
  \876GAT(438) ,
  \754GAT(327) ,
  \849GAT(411) ,
  \424GAT(174) ,
  \270GAT(111) ,
  \741GAT(345) ,
  \573GAT(248) ,
  \793GAT(364) ,
  \525GAT(213) ,
  \839GAT(394) ,
  \772GAT(358) ,
  \677GAT(311) ,
  \697GAT(301) ,
  \743GAT(323) ,
  \521GAT(207) ,
  \738GAT(347) ,
  \529GAT(209) ,
  \537GAT(244) ,
  \806GAT(379) ,
  \853GAT(413) ,
  \404GAT(154) ,
  \712GAT(292) ,
  \635GAT(274) ,
  \375GAT(137) ,
  \356GAT(122) ,
  \832GAT(399) ,
  \651GAT(271) ,
  \444GAT(170) ,
  \349GAT(134) ,
  \323GAT(104) ,
  \713GAT(297) ,
  \585GAT(259) ,
  \536GAT(246) ,
  \565GAT(254) ,
  \287GAT(101) ,
  \596GAT(268) ,
  \854GAT(419) ,
  \451GAT(200) ,
  \516GAT(217) ,
  \517GAT(227) ,
  \547GAT(235) ,
  \670GAT(310) ,
  \807GAT(380) ,
  \795GAT(369) ,
  \842GAT(410) ,
  \351GAT(125) ,
  \877GAT(437) ,
  \739GAT(332) ,
  \766GAT(344) ,
  \520GAT(208) ;
assign
  \569GAT(247)  = ~\540GAT(239)  | ~\488GAT(184) ,
  \425GAT(172)  = \405GAT(152)  & \404GAT(154) ,
  \792GAT(363)  = ~\782GAT(353)  & ~\717GAT(296) ,
  \815GAT(388)  = ~\814GAT(383)  | (~\766GAT(344)  | (~\765GAT(346)  | ~\738GAT(347) )),
  \526GAT(212)  = \183GAT(44)  & \451GAT(200) ,
  \734GAT(287)  = ~\261GAT(57)  | (~\654GAT(270)  | (~\644GAT(272)  | ~\635GAT(274) )),
  \865GAT(422)  = \857GAT(416) ,
  \269GAT(112)  = ~\17GAT(3)  | (~\13GAT(2)  | (~\8GAT(1)  | ~\1GAT(0) )),
  \503GAT(203)  = ~\476GAT(188)  & ~\475GAT(197) ,
  \782GAT(353)  = ~\732GAT(289)  | ~\756GAT(335) ,
  \499GAT(225)  = \460GAT(199)  | \130GAT(31) ,
  \350GAT(126)  = \286GAT(92)  | \280GAT(108) ,
  \696GAT(305)  = ~\525GAT(213)  & ~\624GAT(265) ,
  \765GAT(346)  = ~\678GAT(307)  | ~\600GAT(282) ,
  \420GAT(158)  = \351GAT(125) ,
  \322GAT(105)  = ~\42GAT(7)  & ~\17GAT(3) ,
  \405GAT(152)  = ~\360GAT(120) ,
  \506GAT(232)  = \466GAT(201)  & \101GAT(25) ,
  \773GAT(351)  = ~\734GAT(287)  | (~\763GAT(337)  | (~\762GAT(339)  | ~\750GAT(340) )),
  \844GAT(408)  = ~\835GAT(398)  & ~\834GAT(397) ,
  \478GAT(189)  = \432GAT(181)  & \310GAT(60) ,
  \327GAT(68)  = \177GAT(43)  | \171GAT(42) ,
  \326GAT(69)  = ~\177GAT(43)  | ~\171GAT(42) ,
  \632GAT(275)  = ~\189GAT(45)  | ~\573GAT(248) ,
  \419GAT(164)  = \344GAT(136) ,
  \628GAT(276)  = \183GAT(44)  | \569GAT(247) ,
  \687GAT(304)  = ~\616GAT(279) ,
  \631GAT(264)  = \569GAT(247)  & \246GAT(53) ,
  \353GAT(130)  = ~\295GAT(97) ,
  \336GAT(77)  = \111GAT(27)  & \210GAT(49) ,
  \489GAT(185)  = \437GAT(177)  | \369GAT(113) ,
  \527GAT(211)  = ~\189GAT(45)  | ~\451GAT(200) ,
  \796GAT(373)  = ~\747GAT(341)  | ~\795GAT(369) ,
  \855GAT(418)  = ~\846GAT(407) ,
  \477GAT(196)  = \427GAT(178)  & \146GAT(35) ,
  \498GAT(226)  = ~\460GAT(199)  | ~\130GAT(31) ,
  \338GAT(76)  = \116GAT(28)  & \210GAT(49) ,
  \347GAT(138)  = ~\279GAT(109) ,
  \329GAT(66)  = \189GAT(45)  | \183GAT(44) ,
  \328GAT(67)  = ~\189GAT(45)  | ~\183GAT(44) ,
  \418GAT(168)  = \342GAT(141) ,
  \686GAT(308)  = ~\524GAT(214)  & ~\615GAT(266) ,
  \417GAT(142)  = \369GAT(113)  & \210GAT(49) ,
  \736GAT(333)  = \665GAT(312)  & \228GAT(51) ,
  \747GAT(341)  = ~\697GAT(301) ,
  \757GAT(317)  = ~\261GAT(57)  & ~\727GAT(294) ,
  \360GAT(120)  = ~\304GAT(82)  | ~\303GAT(83) ,
  \864GAT(423)  = \856GAT(417) ,
  \460GAT(199)  = ~\425GAT(172)  & ~\406GAT(153) ,
  \660GAT(315)  = ~\588GAT(286)  & ~\552GAT(258) ,
  \867GAT(432)  = ~\669GAT(314)  | (~\769GAT(361)  | ~\859GAT(421) ),
  \825GAT(385)  = ~\807GAT(380)  & ~\806GAT(379) ,
  \843GAT(409)  = ~\833GAT(400)  & ~\832GAT(399) ,
  \661GAT(293)  = ~\589GAT(269)  & ~\587GAT(256) ,
  \640GAT(263)  = \573GAT(248)  & \246GAT(53) ,
  \346GAT(140)  = ~\276GAT(110) ,
  \421GAT(162)  = \353GAT(130) ,
  \733GAT(288)  = ~\261GAT(57)  | (~\654GAT(270)  | ~\644GAT(272) ),
  \379GAT(116)  = ~\327GAT(68)  | ~\326GAT(69) ,
  \586GAT(255)  = ~\547GAT(235) ,
  \834GAT(397)  = ~\822GAT(386)  & ~\682GAT(306) ,
  \406GAT(153)  = \360GAT(120)  & \357GAT(121) ,
  \751GAT(328)  = \708GAT(298)  & \228GAT(51) ,
  \410GAT(160)  = ~\352GAT(127)  | ~\347GAT(138) ,
  \528GAT(210)  = ~\195GAT(46)  | ~\451GAT(200) ,
  \332GAT(85)  = \91GAT(23)  & \210GAT(49) ,
  \333GAT(84)  = \96GAT(24)  & \210GAT(49) ,
  \340GAT(73)  = \121GAT(29)  & \210GAT(49) ,
  \593GAT(284)  = \159GAT(40)  | \553GAT(251) ,
  \369GAT(113)  = ~\310GAT(60) ,
  \399GAT(166)  = ~\346GAT(140) ,
  \542GAT(237)  = ~\515GAT(228)  & ~\514GAT(218) ,
  \443GAT(180)  = ~\17GAT(3)  | (~\319GAT(90)  | ~\393GAT(165) ),
  \874GAT(433)  = \870GAT(429) ,
  \408GAT(149)  = ~\366GAT(118) ,
  \488GAT(184)  = \437GAT(177)  | \369GAT(113) ,
  \587GAT(256)  = \547GAT(235)  & \544GAT(242) ,
  \794GAT(362)  = \786GAT(350)  & \219GAT(50) ,
  \856GAT(417)  = ~\847GAT(406) ,
  \509GAT(206)  = ~\482GAT(191)  & ~\481GAT(194) ,
  \416GAT(144)  = \385GAT(114)  & \382GAT(115) ,
  \759GAT(326)  = \727GAT(294)  & \228GAT(51) ,
  \758GAT(316)  = \261GAT(57)  & \727GAT(294) ,
  \762GAT(339)  = ~\713GAT(297)  | ~\635GAT(274) ,
  \804GAT(370)  = ~\793GAT(364)  & ~\792GAT(363) ,
  \875GAT(439)  = ~\871GAT(436) ,
  \310GAT(60)  = ~\268GAT(59) ,
  \619GAT(278)  = \177GAT(43)  | \565GAT(254) ,
  \760GAT(318)  = \722GAT(295)  & \237GAT(52) ,
  \442GAT(175)  = ~\393GAT(165)  | (~\156GAT(39)  | (~\59GAT(10)  | ~\375GAT(137) )),
  \344GAT(136)  = \273GAT(103)  | \270GAT(111) ,
  \544GAT(242)  = ~\519GAT(223)  | ~\518GAT(224) ,
  \814GAT(383)  = ~\796GAT(373)  | (~\619GAT(278)  | (~\609GAT(280)  | ~\600GAT(282) )),
  \704GAT(302)  = ~\526GAT(212)  & ~\631GAT(264) ,
  \492GAT(193)  = ~\444GAT(170)  & ~\413GAT(147) ,
  \285GAT(102)  = ~\68GAT(11)  | ~\29GAT(5) ,
  \407GAT(151)  = ~\363GAT(119) ,
  \764GAT(343)  = ~\687GAT(304)  | ~\609GAT(280) ,
  \735GAT(348)  = ~\662GAT(313) ,
  \557GAT(252)  = ~\505GAT(204)  | ~\537GAT(244) ,
  \654GAT(270)  = \201GAT(47)  | \581GAT(250) ,
  \334GAT(81)  = \101GAT(25)  & \210GAT(49) ,
  \335GAT(80)  = \106GAT(26)  & \210GAT(49) ,
  \833GAT(400)  = \819GAT(387)  & \673GAT(309) ,
  \732GAT(289)  = ~\261GAT(57)  | ~\654GAT(270) ,
  \466GAT(201)  = ~\410GAT(160)  | ~\442GAT(175) ,
  \352GAT(127)  = ~\294GAT(94) ,
  \432GAT(181)  = \287GAT(101)  & (\17GAT(3)  & \393GAT(165) ),
  \519GAT(223)  = \492GAT(193)  | \130GAT(31) ,
  \835GAT(398)  = \822GAT(386)  & \682GAT(306) ,
  \476GAT(188)  = \432GAT(181)  & \310GAT(60) ,
  \669GAT(314)  = ~\522GAT(216)  & ~\596GAT(268) ,
  \866GAT(426)  = \858GAT(420) ,
  \504GAT(233)  = \466GAT(201)  & \96GAT(24) ,
  \753GAT(338)  = ~\713GAT(297) ,
  \533GAT(241)  = ~\501GAT(221)  | ~\500GAT(222) ,
  \480GAT(190)  = \432GAT(181)  & \310GAT(60) ,
  \363GAT(119)  = ~\306GAT(78)  | ~\305GAT(79) ,
  \317GAT(106)  = \138GAT(33)  & \17GAT(3) ,
  \589GAT(269)  = \586GAT(255)  & \585GAT(259) ,
  \616GAT(279)  = ~\177GAT(43)  | ~\565GAT(254) ,
  \345GAT(139)  = ~\276GAT(110) ,
  \510GAT(220)  = \483GAT(202)  & \143GAT(34) ,
  \785GAT(355)  = ~\755GAT(319)  & ~\754GAT(327) ,
  \543GAT(236)  = ~\517GAT(227)  & ~\516GAT(217) ,
  \737GAT(325)  = \662GAT(313)  & \237GAT(52) ,
  \615GAT(266)  = \561GAT(253)  & \246GAT(53) ,
  \857GAT(416)  = ~\848GAT(405) ,
  \415GAT(143)  = ~\385GAT(114) ,
  \341GAT(61)  = \267GAT(58)  & \255GAT(54) ,
  \400GAT(157)  = \73GAT(13)  & \348GAT(128) ,
  \763GAT(337)  = ~\722GAT(295)  | (~\644GAT(272)  | ~\635GAT(274) ),
  \448GAT(179)  = \401GAT(163) ,
  \861GAT(427)  = ~\853GAT(413)  & ~\333GAT(84) ,
  \522GAT(216)  = \159GAT(40)  & \451GAT(200) ,
  \318GAT(72)  = \138GAT(33)  & \152GAT(37) ,
  \382GAT(115)  = ~\329GAT(66)  | ~\328GAT(67) ,
  \805GAT(374)  = ~\794GAT(362)  & ~\340GAT(73) ,
  \479GAT(195)  = \427GAT(178)  & \149GAT(36) ,
  \577GAT(249)  = ~\542GAT(237)  | ~\490GAT(186) ,
  \512GAT(219)  = \483GAT(202)  & \146GAT(35) ,
  \513GAT(229)  = \466GAT(201)  & \116GAT(28) ,
  \872GAT(435)  = ~\868GAT(431) ,
  \673GAT(309)  = \597GAT(283)  & \600GAT(282) ,
  \813GAT(382)  = ~\796GAT(373)  | (~\619GAT(278)  | ~\609GAT(280) ),
  \518GAT(224)  = ~\492GAT(193)  | ~\130GAT(31) ,
  \705GAT(299)  = ~\632GAT(275) ,
  \850GAT(404)  = \840GAT(393) ,
  \662GAT(313)  = ~\590GAT(285) ,
  \641GAT(273)  = ~\195GAT(46)  | ~\577GAT(249) ,
  \273GAT(103)  = \42GAT(7)  & (\36GAT(6)  & \29GAT(5) ),
  \609GAT(280)  = \171GAT(42)  | \561GAT(253) ,
  \388GAT(133)  = \290GAT(100) ,
  \845GAT(412)  = ~\836GAT(392)  & ~\334GAT(81) ,
  \717GAT(296)  = \641GAT(273)  & \644GAT(272) ,
  \870GAT(429)  = ~\862GAT(425) ,
  \309GAT(107)  = \138GAT(33)  & \8GAT(1) ,
  \551GAT(257)  = ~\533GAT(241) ,
  \786GAT(350)  = ~\758GAT(316)  & ~\757GAT(317) ,
  \540GAT(239)  = ~\511GAT(230)  & ~\510GAT(220) ,
  \401GAT(163)  = ~\349GAT(134) ,
  \727GAT(294)  = \651GAT(271)  & \654GAT(270) ,
  \290GAT(100)  = \42GAT(7)  & (\75GAT(15)  & \29GAT(5) ),
  \331GAT(64)  = \201GAT(47)  | \195GAT(46) ,
  \330GAT(65)  = ~\201GAT(47)  | ~\195GAT(46) ,
  \501GAT(221)  = \135GAT(32)  | \463GAT(198) ,
  \413GAT(147)  = \379GAT(116)  & \376GAT(117) ,
  \297GAT(89)  = \86GAT(18)  & \85GAT(17) ,
  \414GAT(145)  = ~\382GAT(115) ,
  \777GAT(357)  = ~\749GAT(321)  & ~\748GAT(329) ,
  \481GAT(194)  = \427GAT(178)  & \153GAT(38) ,
  \812GAT(381)  = ~\796GAT(373)  | ~\619GAT(278) ,
  \561GAT(253)  = ~\507GAT(205)  | ~\538GAT(245) ,
  \822GAT(386)  = ~\812GAT(381)  | ~\744GAT(342) ,
  \422GAT(161)  = \354GAT(129) ,
  \860GAT(428)  = ~\852GAT(414)  & ~\332GAT(85) ,
  \550GAT(260)  = ~\530GAT(243) ,
  \859GAT(421)  = ~\851GAT(415)  & ~\417GAT(142) ,
  \624GAT(265)  = \565GAT(254)  & \246GAT(53) ,
  \502GAT(234)  = \466GAT(201)  & \91GAT(23) ,
  \745GAT(330)  = \692GAT(303)  & \228GAT(51) ,
  \339GAT(62)  = \260GAT(56)  & \255GAT(54) ,
  \298GAT(88)  = \88GAT(20)  | \87GAT(19) ,
  \659GAT(261)  = \581GAT(250)  & \246GAT(53) ,
  \423GAT(155)  = \356GAT(122) ,
  \409GAT(150)  = \366GAT(118)  & \363GAT(119) ,
  \507GAT(205)  = ~\480GAT(190)  & ~\479GAT(195) ,
  \841GAT(403)  = ~\593GAT(284)  | ~\815GAT(388) ,
  \449GAT(176)  = \402GAT(159) ,
  \325GAT(70)  = \165GAT(41)  | \159GAT(40) ,
  \324GAT(71)  = ~\165GAT(41)  | ~\159GAT(40) ,
  \819GAT(387)  = ~\813GAT(382)  | (~\764GAT(343)  | ~\741GAT(345) ),
  \355GAT(123)  = ~\298GAT(88)  | ~\89GAT(21) ,
  \463GAT(198)  = ~\426GAT(171)  & ~\409GAT(150) ,
  \836GAT(392)  = \825GAT(385)  & \219GAT(50) ,
  \791GAT(366)  = \778GAT(352)  & \708GAT(298) ,
  \873GAT(434)  = ~\869GAT(430) ,
  \692GAT(303)  = \616GAT(279)  & \619GAT(278) ,
  \354GAT(129)  = ~\296GAT(96) ,
  \581GAT(250)  = ~\543GAT(236)  | ~\491GAT(187) ,
  \337GAT(63)  = \259GAT(55)  & \255GAT(54) ,
  \744GAT(342)  = ~\687GAT(304) ,
  \746GAT(322)  = \687GAT(304)  & \237GAT(52) ,
  \802GAT(372)  = ~\789GAT(368)  & ~\788GAT(367) ,
  \303GAT(83)  = ~\106GAT(26)  | ~\101GAT(25) ,
  \552GAT(258)  = \533GAT(241)  & \530GAT(243) ,
  \482GAT(191)  = \432GAT(181)  & \310GAT(60) ,
  \389GAT(132)  = \291GAT(99) ,
  \837GAT(396)  = ~\704GAT(302)  | (~\777GAT(357)  | ~\826GAT(391) ),
  \426GAT(171)  = \408GAT(149)  & \407GAT(151) ,
  \393GAT(165)  = ~\345GAT(139) ,
  \295GAT(97)  = \80GAT(16)  & (\36GAT(6)  & \59GAT(10) ),
  \590GAT(285)  = ~\159GAT(40)  | ~\553GAT(251) ,
  \742GAT(331)  = \682GAT(306)  & \228GAT(51) ,
  \523GAT(215)  = \165GAT(41)  & \451GAT(200) ,
  \286GAT(92)  = ~\74GAT(14)  | (~\68GAT(11)  | ~\59GAT(10) ),
  \348GAT(128)  = ~\284GAT(95)  & ~\280GAT(108) ,
  \831GAT(402)  = \815GAT(388)  & \665GAT(312) ,
  \296GAT(96)  = \42GAT(7)  & (\36GAT(6)  & \59GAT(10) ),
  \284GAT(95)  = ~\72GAT(12)  | (~\68GAT(11)  | (~\42GAT(7)  | ~\59GAT(10) )),
  \541GAT(238)  = ~\513GAT(229)  & ~\512GAT(219) ,
  \279GAT(109)  = ~\17GAT(3)  | (~\51GAT(8)  | (~\8GAT(1)  | ~\1GAT(0) )),
  \605GAT(267)  = \557GAT(252)  & \246GAT(53) ,
  \749GAT(321)  = \697GAT(301)  & \237GAT(52) ,
  \293GAT(91)  = \80GAT(16)  & (\75GAT(15)  & \59GAT(10) ),
  \539GAT(240)  = ~\508GAT(231)  & ~\318GAT(72) ,
  \412GAT(146)  = ~\379GAT(116) ,
  \402GAT(159)  = ~\350GAT(126) ,
  \511GAT(230)  = \466GAT(201)  & \111GAT(27) ,
  \445GAT(169)  = \415GAT(143)  & \414GAT(145) ,
  \682GAT(306)  = \606GAT(281)  & \609GAT(280) ,
  \768GAT(334)  = \661GAT(293) ,
  \342GAT(141)  = ~\269GAT(112) ,
  \787GAT(354)  = ~\760GAT(318)  & ~\759GAT(326) ,
  \392GAT(167)  = \343GAT(135)  | \270GAT(111) ,
  \495GAT(192)  = ~\445GAT(169)  & ~\416GAT(144) ,
  \600GAT(282)  = \165GAT(41)  | \557GAT(252) ,
  \803GAT(371)  = ~\791GAT(366)  & ~\790GAT(365) ,
  \826GAT(391)  = ~\808GAT(377)  & ~\335GAT(80) ,
  \750GAT(340)  = ~\705GAT(299) ,
  \752GAT(320)  = \705GAT(299)  & \237GAT(52) ,
  \851GAT(415)  = \842GAT(410)  & \219GAT(50) ,
  \858GAT(420)  = ~\849GAT(411) ,
  \761GAT(336)  = ~\722GAT(295)  | ~\644GAT(272) ,
  \810GAT(375)  = \804GAT(370)  & \219GAT(50) ,
  \427GAT(178)  = \55GAT(9)  & (\393GAT(165)  & \319GAT(90) ),
  \301GAT(87)  = ~\96GAT(24)  | ~\91GAT(23) ,
  \304GAT(82)  = \106GAT(26)  | \101GAT(25) ,
  \343GAT(135)  = ~\273GAT(103) ,
  \789GAT(368)  = \773GAT(351)  & \700GAT(300) ,
  \500GAT(222)  = ~\135GAT(32)  | ~\463GAT(198) ,
  \879GAT(441)  = \876GAT(438) ,
  \830GAT(401)  = ~\815GAT(388)  & ~\665GAT(312) ,
  \302GAT(86)  = \96GAT(24)  | \91GAT(23) ,
  \848GAT(405)  = ~\839GAT(394) ,
  \316GAT(93)  = \138GAT(33)  & \51GAT(8) ,
  \319GAT(90)  = ~\156GAT(39)  | ~\59GAT(10) ,
  \748GAT(329)  = \700GAT(300)  & \228GAT(51) ,
  \292GAT(98)  = \42GAT(7)  & (\36GAT(6)  & \29GAT(5) ),
  \276GAT(110)  = \51GAT(8)  & (\26GAT(4)  & \1GAT(0) ),
  \597GAT(283)  = ~\165GAT(41)  | ~\557GAT(252) ,
  \491GAT(187)  = \437GAT(177)  | \369GAT(113) ,
  \829GAT(384)  = ~\811GAT(378) ,
  \306GAT(78)  = \116GAT(28)  | \111GAT(27) ,
  \811GAT(378)  = ~\529GAT(209)  | (~\731GAT(290)  | (~\787GAT(354)  | ~\805GAT(374) )),
  \721GAT(291)  = ~\650GAT(262)  & ~\339GAT(62) ,
  \625GAT(277)  = ~\183GAT(44)  | ~\569GAT(247) ,
  \291GAT(99)  = \80GAT(16)  & (\36GAT(6)  & \29GAT(5) ),
  \294GAT(94)  = \42GAT(7)  & (\75GAT(15)  & \59GAT(10) ),
  \808GAT(377)  = \802GAT(372)  & \219GAT(50) ,
  \700GAT(300)  = \625GAT(277)  & \628GAT(276) ,
  \305GAT(79)  = ~\116GAT(28)  | ~\111GAT(27) ,
  \514GAT(218)  = \483GAT(202)  & \149GAT(36) ,
  \515GAT(228)  = \466GAT(201)  & \121GAT(29) ,
  \847GAT(406)  = ~\838GAT(395) ,
  \828GAT(389)  = ~\810GAT(375)  & ~\338GAT(76) ,
  \437GAT(177)  = ~\55GAT(9)  | (~\287GAT(101)  | ~\393GAT(165) ),
  \868GAT(431)  = ~\677GAT(311)  | (~\770GAT(360)  | ~\860GAT(428) ),
  \778GAT(352)  = ~\733GAT(288)  | (~\761GAT(336)  | ~\753GAT(338) ),
  \880GAT(440)  = \877GAT(437) ,
  \411GAT(148)  = ~\376GAT(117) ,
  \871GAT(436)  = ~\867GAT(432) ,
  \863GAT(424)  = \855GAT(418) ,
  \447GAT(182)  = \399GAT(166) ,
  \650GAT(262)  = \577GAT(249)  & \246GAT(53) ,
  \588GAT(286)  = \551GAT(257)  & \550GAT(260) ,
  \790GAT(365)  = ~\778GAT(352)  & ~\708GAT(298) ,
  \366GAT(118)  = ~\308GAT(74)  | ~\307GAT(75) ,
  \524GAT(214)  = \171GAT(42)  & \451GAT(200) ,
  \357GAT(121)  = ~\302GAT(86)  | ~\301GAT(87) ,
  \838GAT(395)  = ~\527GAT(211)  | (~\712GAT(292)  | (~\781GAT(356)  | ~\827GAT(390) )),
  \771GAT(359)  = ~\743GAT(323)  & ~\742GAT(331) ,
  \740GAT(324)  = \670GAT(310)  & \237GAT(52) ,
  \530GAT(243)  = ~\499GAT(225)  | ~\498GAT(226) ,
  \553GAT(251)  = ~\503GAT(203)  | ~\536GAT(246) ,
  \508GAT(231)  = \466GAT(201)  & \106GAT(26) ,
  \308GAT(74)  = \126GAT(30)  | \121GAT(29) ,
  \538GAT(245)  = ~\506GAT(232)  & ~\317GAT(106) ,
  \403GAT(156)  = ~\355GAT(123) ,
  \280GAT(108)  = ~\55GAT(9)  | (~\13GAT(2)  | (~\8GAT(1)  | ~\1GAT(0) )),
  \644GAT(272)  = \195GAT(46)  | \577GAT(249) ,
  \767GAT(349)  = \660GAT(315) ,
  \827GAT(390)  = ~\809GAT(376)  & ~\336GAT(77) ,
  \307GAT(75)  = ~\126GAT(30)  | ~\121GAT(29) ,
  \852GAT(414)  = \843GAT(409)  & \219GAT(50) ,
  \708GAT(298)  = \632GAT(275)  & \635GAT(274) ,
  \606GAT(281)  = ~\171GAT(42)  | ~\561GAT(253) ,
  \391GAT(124)  = \297GAT(89) ,
  \788GAT(367)  = ~\773GAT(351)  & ~\700GAT(300) ,
  \505GAT(204)  = ~\478GAT(189)  & ~\477GAT(196) ,
  \376GAT(117)  = ~\325GAT(70)  | ~\324GAT(71) ,
  \483GAT(202)  = ~\1GAT(0)  | ~\443GAT(180) ,
  \769GAT(361)  = ~\737GAT(325)  & ~\736GAT(333) ,
  \385GAT(114)  = ~\331GAT(64)  | ~\330GAT(65) ,
  \490GAT(186)  = \437GAT(177)  | \369GAT(113) ,
  \756GAT(335)  = ~\722GAT(295) ,
  \770GAT(360)  = ~\740GAT(324)  & ~\739GAT(332) ,
  \846GAT(407)  = ~\837GAT(396) ,
  \781GAT(356)  = ~\752GAT(320)  & ~\751GAT(328) ,
  \809GAT(376)  = \803GAT(371)  & \219GAT(50) ,
  \475GAT(197)  = \427GAT(178)  & \143GAT(34) ,
  \678GAT(307)  = ~\606GAT(281) ,
  \665GAT(312)  = \590GAT(285)  & \593GAT(284) ,
  \840GAT(393)  = ~\829GAT(384) ,
  \878GAT(442)  = \875GAT(439) ,
  \722GAT(295)  = ~\651GAT(271) ,
  \862GAT(425)  = ~\854GAT(419) ,
  \731GAT(290)  = ~\659GAT(261)  & ~\341GAT(61) ,
  \869GAT(430)  = ~\686GAT(308)  | (~\771GAT(359)  | ~\861GAT(427) ),
  \755GAT(319)  = \713GAT(297)  & \237GAT(52) ,
  \446GAT(183)  = \392GAT(167) ,
  \876GAT(438)  = ~\872GAT(435) ,
  \754GAT(327)  = \717GAT(296)  & \228GAT(51) ,
  \849GAT(411)  = \841GAT(403)  & \735GAT(348) ,
  \424GAT(174)  = ~\400GAT(157) ,
  \270GAT(111)  = ~\17GAT(3)  | (~\13GAT(2)  | (~\26GAT(4)  | ~\1GAT(0) )),
  \741GAT(345)  = ~\678GAT(307) ,
  \573GAT(248)  = ~\541GAT(238)  | ~\489GAT(185) ,
  \793GAT(364)  = \782GAT(353)  & \717GAT(296) ,
  \525GAT(213)  = \177GAT(43)  & \451GAT(200) ,
  \839GAT(394)  = ~\528GAT(210)  | (~\721GAT(291)  | (~\785GAT(355)  | ~\828GAT(389) )),
  \772GAT(358)  = ~\746GAT(322)  & ~\745GAT(330) ,
  \677GAT(311)  = ~\523GAT(215)  & ~\605GAT(267) ,
  \697GAT(301)  = ~\625GAT(277) ,
  \743GAT(323)  = \678GAT(307)  & \237GAT(52) ,
  \521GAT(207)  = \207GAT(48)  | \495GAT(192) ,
  \738GAT(347)  = ~\670GAT(310) ,
  \529GAT(209)  = ~\201GAT(47)  | ~\451GAT(200) ,
  \537GAT(244)  = ~\504GAT(233)  & ~\316GAT(93) ,
  \806GAT(379)  = ~\796GAT(373)  & ~\692GAT(303) ,
  \853GAT(413)  = \844GAT(408)  & \219GAT(50) ,
  \404GAT(154)  = ~\357GAT(121) ,
  \712GAT(292)  = ~\640GAT(263)  & ~\337GAT(63) ,
  \635GAT(274)  = \189GAT(45)  | \573GAT(248) ,
  \375GAT(137)  = ~\323GAT(104)  & ~\322GAT(105) ,
  \356GAT(122)  = \298GAT(88)  & \90GAT(22) ,
  \832GAT(399)  = ~\819GAT(387)  & ~\673GAT(309) ,
  \651GAT(271)  = ~\201GAT(47)  | ~\581GAT(250) ,
  \444GAT(170)  = \412GAT(146)  & \411GAT(148) ,
  \349GAT(134)  = \285GAT(102)  | \280GAT(108) ,
  \323GAT(104)  = \42GAT(7)  & \17GAT(3) ,
  \713GAT(297)  = ~\641GAT(273) ,
  \585GAT(259)  = ~\544GAT(242) ,
  \536GAT(246)  = ~\502GAT(234)  & ~\309GAT(107) ,
  \565GAT(254)  = ~\509GAT(206)  | ~\539GAT(240) ,
  \287GAT(101)  = \80GAT(16)  & (\75GAT(15)  & \29GAT(5) ),
  \596GAT(268)  = \553GAT(251)  & \246GAT(53) ,
  \854GAT(419)  = ~\696GAT(305)  | (~\772GAT(358)  | ~\845GAT(412) ),
  \451GAT(200)  = ~\424GAT(174) ,
  \516GAT(217)  = \483GAT(202)  & \153GAT(38) ,
  \517GAT(227)  = \466GAT(201)  & \126GAT(30) ,
  \547GAT(235)  = ~\521GAT(207)  | ~\520GAT(208) ,
  \670GAT(310)  = ~\597GAT(283) ,
  \450GAT(173)  = \403GAT(156) ,
  \807GAT(380)  = \796GAT(373)  & \692GAT(303) ,
  \795GAT(369)  = ~\773GAT(351)  | ~\628GAT(276) ,
  \842GAT(410)  = ~\831GAT(402)  & ~\830GAT(401) ,
  \351GAT(125)  = ~\293GAT(91) ,
  \877GAT(437)  = ~\873GAT(434) ,
  \739GAT(332)  = \673GAT(309)  & \228GAT(51) ,
  \390GAT(131)  = \292GAT(98) ,
  \766GAT(344)  = ~\687GAT(304)  | (~\609GAT(280)  | ~\600GAT(282) ),
  \520GAT(208)  = ~\207GAT(48)  | ~\495GAT(192) ;
endmodule

