// IWLS benchmark module "C499.iscas" printed on Wed May 29 16:29:38 2002
module C499 (\ID0(0) , \ID1(1) , \ID2(2) , \ID3(3) , \ID4(4) , \ID5(5) , \ID6(6) , \ID7(7) , \ID8(8) , \ID9(9) , \ID10(10) , \ID11(11) , \ID12(12) , \ID13(13) , \ID14(14) , \ID15(15) , \ID16(16) , \ID17(17) , \ID18(18) , \ID19(19) , \ID20(20) , \ID21(21) , \ID22(22) , \ID23(23) , \ID24(24) , \ID25(25) , \ID26(26) , \ID27(27) , \ID28(28) , \ID29(29) , \ID30(30) , \ID31(31) , \IC0(32) , \IC1(33) , \IC2(34) , \IC3(35) , \IC4(36) , \IC5(37) , \IC6(38) , \IC7(39) , \R(40) , \OD0(242) , \OD1(241) , \OD2(240) , \OD3(239) , \OD4(238) , \OD5(237) , \OD6(236) , \OD7(235) , \OD8(234) , \OD9(233) , \OD10(232) , \OD11(231) , \OD12(230) , \OD13(229) , \OD14(228) , \OD15(227) , \OD16(226) , \OD17(225) , \OD18(224) , \OD19(223) , \OD20(222) , \OD21(221) , \OD22(220) , \OD23(219) , \OD24(218) , \OD25(217) , \OD26(216) , \OD27(215) , \OD28(214) , \OD29(213) , \OD30(212) , \OD31(211) );
input
  \ID0(0) ,
  \ID10(10) ,
  \ID21(21) ,
  \ID26(26) ,
  \R(40) ,
  \ID1(1) ,
  \ID15(15) ,
  \IC0(32) ,
  \IC6(38) ,
  \ID2(2) ,
  \ID3(3) ,
  \ID20(20) ,
  \ID31(31) ,
  \ID4(4) ,
  \ID14(14) ,
  \IC5(37) ,
  \ID25(25) ,
  \ID5(5) ,
  \ID19(19) ,
  \ID6(6) ,
  \ID13(13) ,
  \ID7(7) ,
  \ID30(30) ,
  \IC4(36) ,
  \ID24(24) ,
  \ID8(8) ,
  \ID18(18) ,
  \ID29(29) ,
  \ID9(9) ,
  \IC3(35) ,
  \ID12(12) ,
  \ID23(23) ,
  \ID17(17) ,
  \ID28(28) ,
  \IC2(34) ,
  \ID22(22) ,
  \ID11(11) ,
  \ID16(16) ,
  \ID27(27) ,
  \IC1(33) ,
  \IC7(39) ;
output
  \OD21(221) ,
  \OD13(229) ,
  \OD22(220) ,
  \OD14(228) ,
  \OD0(242) ,
  \OD1(241) ,
  \OD15(227) ,
  \OD17(225) ,
  \OD2(240) ,
  \OD30(212) ,
  \OD16(226) ,
  \OD18(224) ,
  \OD31(211) ,
  \OD23(219) ,
  \OD19(223) ,
  \OD24(218) ,
  \OD3(239) ,
  \OD25(217) ,
  \OD27(215) ,
  \OD4(238) ,
  \OD10(232) ,
  \OD26(216) ,
  \OD28(214) ,
  \OD5(237) ,
  \OD11(231) ,
  \OD29(213) ,
  \OD6(236) ,
  \OD7(235) ,
  \OD12(230) ,
  \OD8(234) ,
  \OD9(233) ,
  \OD20(222) ;
wire
  \XD5(107) ,
  \XD0(112) ,
  \WA(173) ,
  \Y7D(123) ,
  \Y0B(157) ,
  \XA10(58) ,
  \G3(102) ,
  \XD6(106) ,
  \XC2(68) ,
  \F6(84) ,
  \H4(44) ,
  \[0] ,
  \[1] ,
  \XE4(86) ,
  \XC6(52) ,
  \[2] ,
  \XB2(76) ,
  \[3] ,
  \[4] ,
  \Y0C(158) ,
  \Y2C(147) ,
  \F1(95) ,
  \G7(98) ,
  \[5] ,
  \WB(171) ,
  \E28(194) ,
  \XD1(111) ,
  \[6] ,
  \T1(166) ,
  \[7] ,
  \[8] ,
  \E9(205) ,
  \[9] ,
  \XA6(66) ,
  \G4(100) ,
  \E29(190) ,
  \E8(209) ,
  \WC(174) ,
  \E7(196) ,
  \XD7(105) ,
  \XD2(110) ,
  \XB6(60) ,
  \Y2D(148) ,
  \XA1(77) ,
  \T2(167) ,
  \E10(201) ,
  \WD(172) ,
  \Y6J(129) ,
  \Y1A(151) ,
  \H3(45) ,
  \Y1B(152) ,
  \F5(87) ,
  \Y2L(150) ,
  \E11(197) ,
  \Y4K(139) ,
  \Y4L(140) ,
  \S0(120) ,
  \XC5(54) ,
  \S1(119) ,
  \XB1(78) ,
  \T3(168) ,
  \T4(161) ,
  \F0(96) ,
  \G6(99) ,
  \XC1(70) ,
  \XB5(62) ,
  \Y3B(141) ,
  \T5(162) ,
  \[10] ,
  \E13(206) ,
  \Y3C(142) ,
  \U0(170) ,
  \[11] ,
  \U1(169) ,
  \XE3(90) ,
  \XA5(69) ,
  \[12] ,
  \Y5I(134) ,
  \[13] ,
  \XA14(50) ,
  \[14] ,
  \S2(118) ,
  \[15] ,
  \[16] ,
  \WF(175) ,
  \E21(188) ,
  \WE(177) ,
  \[17] ,
  \Y7I(124) ,
  \[18] ,
  \T6(163) ,
  \[19] ,
  \Y1D(153) ,
  \S3(117) ,
  \Y3D(143) ,
  \XE7(82) ,
  \Y5J(135) ,
  \H2(46) ,
  \E12(210) ,
  \F4(88) ,
  \XC4(55) ,
  \XA0(80) ,
  \[20] ,
  \XB0(79) ,
  \G5(97) ,
  \[21] ,
  \XC0(71) ,
  \[22] ,
  \[23] ,
  \H7(41) ,
  \S5(115) ,
  \XB4(63) ,
  \E20(192) ,
  \Y4A(136) ,
  \[24] ,
  \T7(164) ,
  \S4(116) ,
  \[25] ,
  \E30(186) ,
  \XA13(53) ,
  \E14(202) ,
  \[26] ,
  \XE2(91) ,
  \[27] ,
  \E1(203) ,
  \[28] ,
  \Y6A(126) ,
  \[29] ,
  \E0(207) ,
  \Y7K(125) ,
  \XA9(61) ,
  \XA4(72) ,
  \E22(184) ,
  \WG(178) ,
  \S6(114) ,
  \Y4B(137) ,
  \E15(198) ,
  \[30] ,
  \[31] ,
  \E23(180) ,
  \XE6(83) ,
  \WH(176) ,
  \E17(187) ,
  \S7(113) ,
  \H1(47) ,
  \F3(89) ,
  \XA12(56) ,
  \Y2J(149) ,
  \XE1(93) ,
  \Y4C(138) ,
  \E19(179) ,
  \E31(182) ,
  \H6(42) ,
  \Y6C(127) ,
  \E25(189) ,
  \XA8(64) ,
  \XA15(49) ,
  \Y0K(159) ,
  \Y0L(160) ,
  \XA3(73) ,
  \E16(191) ,
  \Y6D(128) ,
  \E3(195) ,
  \Y5A(131) ,
  \E18(183) ,
  \Y1I(154) ,
  \E24(193) ,
  \Y3I(144) ,
  \XE5(85) ,
  \E2(199) ,
  \Y5B(132) ,
  \XB3(75) ,
  \G0(104) ,
  \H0(48) ,
  \Y6L(130) ,
  \E5(204) ,
  \XA11(57) ,
  \XD3(109) ,
  \XC3(67) ,
  \F7(81) ,
  \E4(208) ,
  \XE0(94) ,
  \H5(43) ,
  \E26(185) ,
  \Y1J(155) ,
  \XA7(65) ,
  \F2(92) ,
  \Y7B(121) ,
  \XD4(108) ,
  \E27(181) ,
  \Y7C(122) ,
  \XB7(59) ,
  \XA2(74) ,
  \Y0A(156) ,
  \G1(101) ,
  \E6(200) ,
  \XC7(51) ,
  \Y2A(146) ,
  \T0(165) ,
  \G2(103) ,
  \Y3K(145) ,
  \Y5D(133) ;
assign
  \XD5(107)  = (~\G1(101)  & \H5(43) ) | (\G1(101)  & ~\H5(43) ),
  \XD0(112)  = (~\G4(100)  & \H0(48) ) | (\G4(100)  & ~\H0(48) ),
  \WA(173)  = \U0(170)  & (\Y7I(124)  & (\S6(114)  & (\Y5I(134)  & \S4(116) ))),
  \Y7D(123)  = ~\S7(113) ,
  \Y0B(157)  = ~\S0(120) ,
  \XA10(58)  = (~\ID21(21)  & \ID20(20) ) | (\ID21(21)  & ~\ID20(20) ),
  \G3(102)  = (~\F3(89)  & \F1(95) ) | (\F3(89)  & ~\F1(95) ),
  \OD21(221)  = \[21] ,
  \XD6(106)  = (~\G2(103)  & \H6(42) ) | (\G2(103)  & ~\H6(42) ),
  \OD13(229)  = \[13] ,
  \XC2(68)  = (~\ID14(14)  & \ID10(10) ) | (\ID14(14)  & ~\ID10(10) ),
  \F6(84)  = (~\XA13(53)  & \XA12(56) ) | (\XA13(53)  & ~\XA12(56) ),
  \H4(44)  = \R(40)  & \IC4(36) ,
  \[0]  = (~\E0(207)  & \ID0(0) ) | (\E0(207)  & ~\ID0(0) ),
  \[1]  = (~\E1(203)  & \ID1(1) ) | (\E1(203)  & ~\ID1(1) ),
  \XE4(86)  = (~\XC4(55)  & \XB4(63) ) | (\XC4(55)  & ~\XB4(63) ),
  \XC6(52)  = (~\ID30(30)  & \ID26(26) ) | (\ID30(30)  & ~\ID26(26) ),
  \[2]  = (~\E2(199)  & \ID2(2) ) | (\E2(199)  & ~\ID2(2) ),
  \XB2(76)  = (~\ID6(6)  & \ID2(2) ) | (\ID6(6)  & ~\ID2(2) ),
  \[3]  = (~\E3(195)  & \ID3(3) ) | (\E3(195)  & ~\ID3(3) ),
  \[4]  = (~\E4(208)  & \ID4(4) ) | (\E4(208)  & ~\ID4(4) ),
  \Y0C(158)  = ~\S0(120) ,
  \Y2C(147)  = ~\S2(118) ,
  \F1(95)  = (~\XA3(73)  & \XA2(74) ) | (\XA3(73)  & ~\XA2(74) ),
  \G7(98)  = (~\F7(81)  & \F5(87) ) | (\F7(81)  & ~\F5(87) ),
  \[5]  = (~\E5(204)  & \ID5(5) ) | (\E5(204)  & ~\ID5(5) ),
  \WB(171)  = \U0(170)  & (\S7(113)  & (\Y6J(129)  & (\Y5J(135)  & \S4(116) ))),
  \E28(194)  = \WH(176)  & \S4(116) ,
  \XD1(111)  = (~\G5(97)  & \H1(47) ) | (\G5(97)  & ~\H1(47) ),
  \[6]  = (~\E6(200)  & \ID6(6) ) | (\E6(200)  & ~\ID6(6) ),
  \T1(166)  = \Y3B(141)  & (\S2(118)  & (\Y1B(152)  & \Y0B(157) )),
  \[7]  = (~\E7(196)  & \ID7(7) ) | (\E7(196)  & ~\ID7(7) ),
  \OD22(220)  = \[22] ,
  \OD14(228)  = \[14] ,
  \[8]  = (~\E8(209)  & \ID8(8) ) | (\E8(209)  & ~\ID8(8) ),
  \E9(205)  = \WC(174)  & \S1(119) ,
  \[9]  = (~\E9(205)  & \ID9(9) ) | (\E9(205)  & ~\ID9(9) ),
  \OD0(242)  = \[0] ,
  \XA6(66)  = (~\ID13(13)  & \ID12(12) ) | (\ID13(13)  & ~\ID12(12) ),
  \G4(100)  = (~\F5(87)  & \F4(88) ) | (\F5(87)  & ~\F4(88) ),
  \E29(190)  = \WH(176)  & \S5(115) ,
  \E8(209)  = \WC(174)  & \S0(120) ,
  \WC(174)  = \U0(170)  & (\Y7K(125)  & (\S6(114)  & (\S5(115)  & \Y4K(139) ))),
  \E7(196)  = \WB(171)  & \S3(117) ,
  \OD1(241)  = \[1] ,
  \XD7(105)  = (~\G3(102)  & \H7(41) ) | (\G3(102)  & ~\H7(41) ),
  \XD2(110)  = (~\G6(99)  & \H2(46) ) | (\G6(99)  & ~\H2(46) ),
  \XB6(60)  = (~\ID22(22)  & \ID18(18) ) | (\ID22(22)  & ~\ID18(18) ),
  \Y2D(148)  = ~\S2(118) ,
  \XA1(77)  = (~\ID3(3)  & \ID2(2) ) | (\ID3(3)  & ~\ID2(2) ),
  \T2(167)  = \Y3C(142)  & (\Y2C(147)  & (\S1(119)  & \Y0C(158) )),
  \E10(201)  = \WC(174)  & \S2(118) ,
  \OD15(227)  = \[15] ,
  \WD(172)  = \U0(170)  & (\S7(113)  & (\Y6L(130)  & (\S5(115)  & \Y4L(140) ))),
  \Y6J(129)  = ~\S6(114) ,
  \Y1A(151)  = ~\S1(119) ,
  \H3(45)  = \R(40)  & \IC3(35) ,
  \Y1B(152)  = ~\S1(119) ,
  \OD17(225)  = \[17] ,
  \OD2(240)  = \[2] ,
  \F5(87)  = (~\XA11(57)  & \XA10(58) ) | (\XA11(57)  & ~\XA10(58) ),
  \Y2L(150)  = ~\S2(118) ,
  \E11(197)  = \WC(174)  & \S3(117) ,
  \Y4K(139)  = ~\S4(116) ,
  \Y4L(140)  = ~\S4(116) ,
  \S0(120)  = (~\XD0(112)  & \XE0(94) ) | (\XD0(112)  & ~\XE0(94) ),
  \XC5(54)  = (~\ID29(29)  & \ID25(25) ) | (\ID29(29)  & ~\ID25(25) ),
  \S1(119)  = (~\XD1(111)  & \XE1(93) ) | (\XD1(111)  & ~\XE1(93) ),
  \XB1(78)  = (~\ID5(5)  & \ID1(1) ) | (\ID5(5)  & ~\ID1(1) ),
  \T3(168)  = \Y3D(143)  & (\Y2D(148)  & (\Y1D(153)  & \S0(120) )),
  \T4(161)  = \S7(113)  & (\Y6A(126)  & (\Y5A(131)  & \Y4A(136) )),
  \F0(96)  = (~\XA1(77)  & \XA0(80) ) | (\XA1(77)  & ~\XA0(80) ),
  \OD30(212)  = \[30] ,
  \G6(99)  = (~\F6(84)  & \F4(88) ) | (\F6(84)  & ~\F4(88) ),
  \OD16(226)  = \[16] ,
  \XC1(70)  = (~\ID13(13)  & \ID9(9) ) | (\ID13(13)  & ~\ID9(9) ),
  \XB5(62)  = (~\ID21(21)  & \ID17(17) ) | (\ID21(21)  & ~\ID17(17) ),
  \Y3B(141)  = ~\S3(117) ,
  \T5(162)  = \Y7B(121)  & (\S6(114)  & (\Y5B(132)  & \Y4B(137) )),
  \[10]  = (~\E10(201)  & \ID10(10) ) | (\E10(201)  & ~\ID10(10) ),
  \E13(206)  = \WD(172)  & \S1(119) ,
  \Y3C(142)  = ~\S3(117) ,
  \U0(170)  = \T3(168)  | (\T2(167)  | (\T1(166)  | \T0(165) )),
  \OD18(224)  = \[18] ,
  \[11]  = (~\E11(197)  & \ID11(11) ) | (\E11(197)  & ~\ID11(11) ),
  \U1(169)  = \T7(164)  | (\T6(163)  | (\T5(162)  | \T4(161) )),
  \XE3(90)  = (~\XC3(67)  & \XB3(75) ) | (\XC3(67)  & ~\XB3(75) ),
  \XA5(69)  = (~\ID11(11)  & \ID10(10) ) | (\ID11(11)  & ~\ID10(10) ),
  \[12]  = (~\E12(210)  & \ID12(12) ) | (\E12(210)  & ~\ID12(12) ),
  \Y5I(134)  = ~\S5(115) ,
  \[13]  = (~\E13(206)  & \ID13(13) ) | (\E13(206)  & ~\ID13(13) ),
  \XA14(50)  = (~\ID29(29)  & \ID28(28) ) | (\ID29(29)  & ~\ID28(28) ),
  \[14]  = (~\E14(202)  & \ID14(14) ) | (\E14(202)  & ~\ID14(14) ),
  \S2(118)  = (~\XD2(110)  & \XE2(91) ) | (\XD2(110)  & ~\XE2(91) ),
  \[15]  = (~\E15(198)  & \ID15(15) ) | (\E15(198)  & ~\ID15(15) ),
  \[16]  = (~\E16(191)  & \ID16(16) ) | (\E16(191)  & ~\ID16(16) ),
  \OD31(211)  = \[31] ,
  \WF(175)  = \U1(169)  & (\S3(117)  & (\Y2J(149)  & (\Y1J(155)  & \S0(120) ))),
  \E21(188)  = \WF(175)  & \S5(115) ,
  \WE(177)  = \U1(169)  & (\Y3I(144)  & (\S2(118)  & (\Y1I(154)  & \S0(120) ))),
  \OD23(219)  = \[23] ,
  \[17]  = (~\E17(187)  & \ID17(17) ) | (\E17(187)  & ~\ID17(17) ),
  \Y7I(124)  = ~\S7(113) ,
  \[18]  = (~\E18(183)  & \ID18(18) ) | (\E18(183)  & ~\ID18(18) ),
  \T6(163)  = \Y7C(122)  & (\Y6C(127)  & (\S5(115)  & \Y4C(138) )),
  \[19]  = (~\E19(179)  & \ID19(19) ) | (\E19(179)  & ~\ID19(19) ),
  \Y1D(153)  = ~\S1(119) ,
  \S3(117)  = (~\XD3(109)  & \XE3(90) ) | (\XD3(109)  & ~\XE3(90) ),
  \Y3D(143)  = ~\S3(117) ,
  \OD19(223)  = \[19] ,
  \XE7(82)  = (~\XC7(51)  & \XB7(59) ) | (\XC7(51)  & ~\XB7(59) ),
  \Y5J(135)  = ~\S5(115) ,
  \H2(46)  = \R(40)  & \IC2(34) ,
  \E12(210)  = \WD(172)  & \S0(120) ,
  \F4(88)  = (~\XA9(61)  & \XA8(64) ) | (\XA9(61)  & ~\XA8(64) ),
  \XC4(55)  = (~\ID28(28)  & \ID24(24) ) | (\ID28(28)  & ~\ID24(24) ),
  \XA0(80)  = (~\ID1(1)  & \ID0(0) ) | (\ID1(1)  & ~\ID0(0) ),
  \[20]  = (~\E20(192)  & \ID20(20) ) | (\E20(192)  & ~\ID20(20) ),
  \XB0(79)  = (~\ID4(4)  & \ID0(0) ) | (\ID4(4)  & ~\ID0(0) ),
  \G5(97)  = (~\F7(81)  & \F6(84) ) | (\F7(81)  & ~\F6(84) ),
  \[21]  = (~\E21(188)  & \ID21(21) ) | (\E21(188)  & ~\ID21(21) ),
  \OD24(218)  = \[24] ,
  \XC0(71)  = (~\ID12(12)  & \ID8(8) ) | (\ID12(12)  & ~\ID8(8) ),
  \[22]  = (~\E22(184)  & \ID22(22) ) | (\E22(184)  & ~\ID22(22) ),
  \[23]  = (~\E23(180)  & \ID23(23) ) | (\E23(180)  & ~\ID23(23) ),
  \H7(41)  = \R(40)  & \IC7(39) ,
  \S5(115)  = (~\XD5(107)  & \XE5(85) ) | (\XD5(107)  & ~\XE5(85) ),
  \XB4(63)  = (~\ID20(20)  & \ID16(16) ) | (\ID20(20)  & ~\ID16(16) ),
  \E20(192)  = \WF(175)  & \S4(116) ,
  \Y4A(136)  = ~\S4(116) ,
  \[24]  = (~\E24(193)  & \ID24(24) ) | (\E24(193)  & ~\ID24(24) ),
  \T7(164)  = \Y7D(123)  & (\Y6D(128)  & (\Y5D(133)  & \S4(116) )),
  \S4(116)  = (~\XD4(108)  & \XE4(86) ) | (\XD4(108)  & ~\XE4(86) ),
  \[25]  = (~\E25(189)  & \ID25(25) ) | (\E25(189)  & ~\ID25(25) ),
  \E30(186)  = \WH(176)  & \S6(114) ,
  \XA13(53)  = (~\ID27(27)  & \ID26(26) ) | (\ID27(27)  & ~\ID26(26) ),
  \E14(202)  = \WD(172)  & \S2(118) ,
  \[26]  = (~\E26(185)  & \ID26(26) ) | (\E26(185)  & ~\ID26(26) ),
  \XE2(91)  = (~\XC2(68)  & \XB2(76) ) | (\XC2(68)  & ~\XB2(76) ),
  \[27]  = (~\E27(181)  & \ID27(27) ) | (\E27(181)  & ~\ID27(27) ),
  \OD3(239)  = \[3] ,
  \E1(203)  = \WA(173)  & \S1(119) ,
  \[28]  = (~\E28(194)  & \ID28(28) ) | (\E28(194)  & ~\ID28(28) ),
  \Y6A(126)  = ~\S6(114) ,
  \[29]  = (~\E29(190)  & \ID29(29) ) | (\E29(190)  & ~\ID29(29) ),
  \E0(207)  = \WA(173)  & \S0(120) ,
  \Y7K(125)  = ~\S7(113) ,
  \XA9(61)  = (~\ID19(19)  & \ID18(18) ) | (\ID19(19)  & ~\ID18(18) ),
  \XA4(72)  = (~\ID9(9)  & \ID8(8) ) | (\ID9(9)  & ~\ID8(8) ),
  \OD25(217)  = \[25] ,
  \E22(184)  = \WF(175)  & \S6(114) ,
  \WG(178)  = \U1(169)  & (\Y3K(145)  & (\S2(118)  & (\S1(119)  & \Y0K(159) ))),
  \S6(114)  = (~\XD6(106)  & \XE6(83) ) | (\XD6(106)  & ~\XE6(83) ),
  \Y4B(137)  = ~\S4(116) ,
  \E15(198)  = \WD(172)  & \S3(117) ,
  \[30]  = (~\E30(186)  & \ID30(30) ) | (\E30(186)  & ~\ID30(30) ),
  \OD27(215)  = \[27] ,
  \[31]  = (~\E31(182)  & \ID31(31) ) | (\E31(182)  & ~\ID31(31) ),
  \E23(180)  = \WF(175)  & \S7(113) ,
  \OD4(238)  = \[4] ,
  \XE6(83)  = (~\XC6(52)  & \XB6(60) ) | (\XC6(52)  & ~\XB6(60) ),
  \WH(176)  = \U1(169)  & (\S3(117)  & (\Y2L(150)  & (\S1(119)  & \Y0L(160) ))),
  \E17(187)  = \WE(177)  & \S5(115) ,
  \OD10(232)  = \[10] ,
  \S7(113)  = (~\XD7(105)  & \XE7(82) ) | (\XD7(105)  & ~\XE7(82) ),
  \H1(47)  = \R(40)  & \IC1(33) ,
  \OD26(216)  = \[26] ,
  \F3(89)  = (~\XA7(65)  & \XA6(66) ) | (\XA7(65)  & ~\XA6(66) ),
  \XA12(56)  = (~\ID25(25)  & \ID24(24) ) | (\ID25(25)  & ~\ID24(24) ),
  \Y2J(149)  = ~\S2(118) ,
  \XE1(93)  = (~\XC1(70)  & \XB1(78) ) | (\XC1(70)  & ~\XB1(78) ),
  \Y4C(138)  = ~\S4(116) ,
  \E19(179)  = \WE(177)  & \S7(113) ,
  \E31(182)  = \WH(176)  & \S7(113) ,
  \H6(42)  = \R(40)  & \IC6(38) ,
  \OD28(214)  = \[28] ,
  \OD5(237)  = \[5] ,
  \Y6C(127)  = ~\S6(114) ,
  \E25(189)  = \WG(178)  & \S5(115) ,
  \OD11(231)  = \[11] ,
  \XA8(64)  = (~\ID17(17)  & \ID16(16) ) | (\ID17(17)  & ~\ID16(16) ),
  \XA15(49)  = (~\ID31(31)  & \ID30(30) ) | (\ID31(31)  & ~\ID30(30) ),
  \Y0K(159)  = ~\S0(120) ,
  \Y0L(160)  = ~\S0(120) ,
  \XA3(73)  = (~\ID7(7)  & \ID6(6) ) | (\ID7(7)  & ~\ID6(6) ),
  \E16(191)  = \WE(177)  & \S4(116) ,
  \OD29(213)  = \[29] ,
  \OD6(236)  = \[6] ,
  \Y6D(128)  = ~\S6(114) ,
  \OD7(235)  = \[7] ,
  \OD12(230)  = \[12] ,
  \E3(195)  = \WA(173)  & \S3(117) ,
  \Y5A(131)  = ~\S5(115) ,
  \E18(183)  = \WE(177)  & \S6(114) ,
  \Y1I(154)  = ~\S1(119) ,
  \E24(193)  = \WG(178)  & \S4(116) ,
  \Y3I(144)  = ~\S3(117) ,
  \XE5(85)  = (~\XC5(54)  & \XB5(62) ) | (\XC5(54)  & ~\XB5(62) ),
  \E2(199)  = \WA(173)  & \S2(118) ,
  \Y5B(132)  = ~\S5(115) ,
  \XB3(75)  = (~\ID7(7)  & \ID3(3) ) | (\ID7(7)  & ~\ID3(3) ),
  \G0(104)  = (~\F1(95)  & \F0(96) ) | (\F1(95)  & ~\F0(96) ),
  \H0(48)  = \R(40)  & \IC0(32) ,
  \Y6L(130)  = ~\S6(114) ,
  \E5(204)  = \WB(171)  & \S1(119) ,
  \XA11(57)  = (~\ID23(23)  & \ID22(22) ) | (\ID23(23)  & ~\ID22(22) ),
  \XD3(109)  = (~\G7(98)  & \H3(45) ) | (\G7(98)  & ~\H3(45) ),
  \XC3(67)  = (~\ID15(15)  & \ID11(11) ) | (\ID15(15)  & ~\ID11(11) ),
  \F7(81)  = (~\XA15(49)  & \XA14(50) ) | (\XA15(49)  & ~\XA14(50) ),
  \E4(208)  = \WB(171)  & \S0(120) ,
  \XE0(94)  = (~\XC0(71)  & \XB0(79) ) | (\XC0(71)  & ~\XB0(79) ),
  \H5(43)  = \R(40)  & \IC5(37) ,
  \E26(185)  = \WG(178)  & \S6(114) ,
  \OD8(234)  = \[8] ,
  \Y1J(155)  = ~\S1(119) ,
  \XA7(65)  = (~\ID15(15)  & \ID14(14) ) | (\ID15(15)  & ~\ID14(14) ),
  \F2(92)  = (~\XA5(69)  & \XA4(72) ) | (\XA5(69)  & ~\XA4(72) ),
  \Y7B(121)  = ~\S7(113) ,
  \XD4(108)  = (~\G0(104)  & \H4(44) ) | (\G0(104)  & ~\H4(44) ),
  \E27(181)  = \WG(178)  & \S7(113) ,
  \Y7C(122)  = ~\S7(113) ,
  \XB7(59)  = (~\ID23(23)  & \ID19(19) ) | (\ID23(23)  & ~\ID19(19) ),
  \XA2(74)  = (~\ID5(5)  & \ID4(4) ) | (\ID5(5)  & ~\ID4(4) ),
  \Y0A(156)  = ~\S0(120) ,
  \G1(101)  = (~\F3(89)  & \F2(92) ) | (\F3(89)  & ~\F2(92) ),
  \E6(200)  = \WB(171)  & \S2(118) ,
  \XC7(51)  = (~\ID31(31)  & \ID27(27) ) | (\ID31(31)  & ~\ID27(27) ),
  \Y2A(146)  = ~\S2(118) ,
  \OD9(233)  = \[9] ,
  \OD20(222)  = \[20] ,
  \T0(165)  = \S3(117)  & (\Y2A(146)  & (\Y1A(151)  & \Y0A(156) )),
  \G2(103)  = (~\F2(92)  & \F0(96) ) | (\F2(92)  & ~\F0(96) ),
  \Y3K(145)  = ~\S3(117) ,
  \Y5D(133)  = ~\S5(115) ;
endmodule

