// IWLS benchmark module "C1908.iscas" printed on Wed May 29 16:27:48 2002
module C1908 (\101(0) , \104(1) , \107(2) , \110(3) , \113(4) , \116(5) , \119(6) , \122(7) , \125(8) , \128(9) , \131(10) , \134(11) , \137(12) , \140(13) , \143(14) , \146(15) , \210(16) , \214(17) , \217(18) , \221(19) , \224(20) , \227(21) , \234(22) , \237(23) , \469(24) , \472(25) , \475(26) , \478(27) , \898(28) , \900(29) , \902(30) , \952(31) , \953(32) , \3(865) , \6(864) , \9(863) , \12(862) , \30(856) , \45(851) , \48(850) , \15(861) , \18(860) , \21(859) , \24(858) , \27(857) , \33(855) , \36(854) , \39(853) , \42(852) , \75(866) , \51(899) , \54(900) , \60(901) , \63(902) , \66(903) , \69(908) , \72(909) , \57(912) );
input
  \472(25) ,
  \143(14) ,
  \134(11) ,
  \125(8) ,
  \217(18) ,
  \902(30) ,
  \110(3) ,
  \128(9) ,
  \113(4) ,
  \475(26) ,
  \146(15) ,
  \137(12) ,
  \953(32) ,
  \234(22) ,
  \116(5) ,
  \221(19) ,
  \101(0) ,
  \478(27) ,
  \469(24) ,
  \119(6) ,
  \237(23) ,
  \104(1) ,
  \898(28) ,
  \952(31) ,
  \900(29) ,
  \224(20) ,
  \107(2) ,
  \227(21) ,
  \140(13) ,
  \131(10) ,
  \214(17) ,
  \122(7) ,
  \210(16) ;
output
  \66(903) ,
  \21(859) ,
  \69(908) ,
  \42(852) ,
  \3(865) ,
  \24(858) ,
  \45(851) ,
  \6(864) ,
  \27(857) ,
  \48(850) ,
  \9(863) ,
  \72(909) ,
  \54(900) ,
  \30(856) ,
  \57(912) ,
  \33(855) ,
  \12(862) ,
  \15(861) ,
  \36(854) ,
  \60(901) ,
  \18(860) ,
  \39(853) ,
  \75(866) ,
  \51(899) ,
  \63(902) ;
wire
  \175(75) ,
  \457(205) ,
  \1485(596) ,
  \529(51) ,
  \521(712) ,
  \728(666) ,
  \355(126) ,
  \1244(138) ,
  \400(563) ,
  \828(771) ,
  \710(728) ,
  \202(61) ,
  \1266(395) ,
  \949(33) ,
  \1394(846) ,
  \428(886) ,
  \1325(481) ,
  \1355(533) ,
  \74(843) ,
  \1039(412) ,
  \1189(550) ,
  \796(755) ,
  \1758(514) ,
  \546(656) ,
  \1304(311) ,
  \832(772) ,
  \1529(787) ,
  \1418(280) ,
  \349(883) ,
  \1030(248) ,
  \449(560) ,
  \361(297) ,
  \1748(305) ,
  \330(134) ,
  \241(54) ,
  \1421(692) ,
  \548(637) ,
  \1589(776) ,
  \273(436) ,
  \1352(499) ,
  \1868(447) ,
  \13(814) ,
  \1362(627) ,
  \1610(64) ,
  \564(654) ,
  \1116(303) ,
  \865(793) ,
  \1215(887) ,
  \1170(295) ,
  \369(117) ,
  \994(330) ,
  \34(807) ,
  \1068(231) ,
  \258(442) ,
  \482(202) ,
  \1253(362) ,
  \1833(123) ,
  \1089(561) ,
  \1629(781) ,
  \1668(332) ,
  \1255(407) ,
  \347(607) ,
  \1357(552) ,
  \281(588) ,
  \62(95) ,
  \1608(133) ,
  \566(277) ,
  \274(453) ,
  \1050(163) ,
  \1504(186) ,
  \1171(369) ,
  \1018(435) ,
  \1417(699) ,
  \1466(108) ,
  \1120(308) ,
  \1822(431) ,
  \756(677) ,
  \1718(213) ,
  \1429(615) ,
  \410(470) ,
  \1557(764) ,
  \1586(70) ,
  \61(896) ,
  \1496(185) ,
  \1278(170) ,
  \524(711) ,
  \1029(682) ,
  \348(625) ,
  \1193(566) ,
  \171(77) ,
  \373(283) ,
  \1782(216) ,
  \1166(194) ,
  \343(492) ,
  \1908(513) ,
  \1225(317) ,
  \873(743) ,
  \1326(523) ,
  \1242(457) ,
  \277(570) ,
  \1220(391) ,
  \1440(337) ,
  \1144(849) ,
  \1164(388) ,
  \1282(324) ,
  \862(38) ,
  \1780(645) ,
  \1577(795) ,
  \1115(346) ,
  \1681(503) ,
  \1530(84) ,
  \573(738) ,
  \1344(534) ,
  \533(704) ,
  \1056(251) ,
  \1785(164) ,
  \1525(760) ,
  \1894(490) ,
  \1686(626) ,
  \16(813) ,
  \1676(496) ,
  \1626(60) ,
  \1892(475) ,
  \1902(491) ,
  \248(55) ,
  \1448(191) ,
  \1643(889) ,
  \663(684) ,
  \911(46) ,
  \37(806) ,
  \1207(177) ,
  \1477(595) ,
  \1814(161) ,
  \1264(287) ,
  \1361(568) ,
  \1393(612) ,
  \1493(579) ,
  \1560(156) ,
  \[0] ,
  \1401(584) ,
  \1385(425) ,
  \1000(410) ,
  \1757(222) ,
  \800(756) ,
  \1111(429) ,
  \[1] ,
  \1489(614) ,
  \[2] ,
  \569(730) ,
  \1232(387) ,
  \1194(206) ,
  \[3] ,
  \1125(558) ,
  \1028(869) ,
  \1130(530) ,
  \1377(460) ,
  \549(655) ,
  \294(415) ,
  \[4] ,
  \1445(693) ,
  \1061(341) ,
  \55(911) ,
  \[5] ,
  \1083(538) ,
  \[6] ,
  \1817(150) ,
  \[7] ,
  \362(315) ,
  \863(783) ,
  \1639(881) ,
  \1049(413) ,
  \1099(554) ,
  \[8] ,
  \1647(840) ,
  \1777(461) ,
  \445(578) ,
  \[9] ,
  \1501(580) ,
  \1117(374) ,
  \1040(249) ,
  \1464(189) ,
  \1701(242) ,
  \1732(313) ,
  \558(636) ,
  \1057(239) ,
  \1025(670) ,
  \1528(171) ,
  \1609(799) ,
  \1433(633) ,
  \510(673) ,
  \413(574) ,
  \1174(268) ,
  \824(770) ,
  \310(451) ,
  \1450(110) ,
  \792(754) ,
  \1035(381) ,
  \536(703) ,
  \1265(400) ,
  \421(657) ,
  \731(676) ,
  \153(87) ,
  \244(53) ,
  \492(204) ,
  \1546(80) ,
  \1221(907) ,
  \1689(581) ,
  \1126(543) ,
  \1386(847) ,
  \67(891) ,
  \390(446) ,
  \1901(510) ,
  \883(748) ,
  \932(40) ,
  \19(812) ,
  \918(45) ,
  \1321(377) ,
  \770(679) ,
  \666(685) ,
  \41(825) ,
  \1461(689) ,
  \969(266) ,
  \788(753) ,
  \1131(593) ,
  \291(157) ,
  \1063(365) ,
  \73(741) ,
  \1413(691) ,
  \1267(426) ,
  \1295(483) ,
  \1200(281) ,
  \1517(759) ,
  \879(746) ,
  \1825(445) ,
  \1861(241) ,
  \20(832) ,
  \259(459) ,
  \1227(351) ,
  \1846(220) ,
  \534(710) ,
  \1158(293) ,
  \1182(236) ,
  \887(819) ,
  \1288(386) ,
  \269(378) ,
  \1750(225) ,
  \297(316) ,
  \1400(871) ,
  \427(880) ,
  \1139(577) ,
  \1772(537) ,
  \1392(872) ,
  \56(93) ,
  \516(686) ,
  \1330(390) ,
  \53(893) ,
  \282(608) ,
  \1844(299) ,
  \508(643) ,
  \49(894) ,
  \909(47) ,
  \1549(763) ,
  \1159(368) ,
  \1458(107) ,
  \513(672) ,
  \1310(375) ,
  \1108(307) ,
  \1350(573) ,
  \2(838) ,
  \1781(480) ,
  \414(591) ,
  \532(698) ,
  \1644(100) ,
  \358(389) ,
  \669(715) ,
  \388(396) ,
  \1238(487) ,
  \1187(507) ,
  \1638(867) ,
  \397(416) ,
  \1869(456) ,
  \979(179) ,
  \1700(322) ,
  \23(831) ,
  \1569(792) ,
  \1773(501) ,
  \1335(114) ,
  \1203(282) ,
  \1134(509) ,
  \1432(336) ,
  \544(620) ,
  \375(906) ,
  \1010(411) ,
  \1632(121) ,
  \44(824) ,
  \552(667) ,
  \231(58) ,
  \165(81) ,
  \1469(690) ,
  \1673(502) ,
  \1368(648) ,
  \1272(300) ,
  \1149(669) ,
  \497(721) ,
  \52(92) ,
  \251(175) ,
  \1082(517) ,
  \299(140) ,
  \1721(119) ,
  \980(261) ,
  \1488(188) ,
  \261(441) ,
  \1749(221) ,
  \431(877) ,
  \893(111) ,
  \1918(632) ,
  \565(276) ,
  \453(599) ,
  \393(548) ,
  \1100(227) ,
  \462(820) ,
  \1256(210) ,
  \1885(233) ,
  \1332(132) ,
  \1473(696) ,
  \509(662) ,
  \1184(370) ,
  \1098(270) ,
  \1838(219) ,
  \1853(238) ,
  \1490(103) ,
  \1649(882) ,
  \1670(472) ,
  \419(683) ,
  \1071(342) ,
  \1405(604) ,
  \1552(159) ,
  \156(85) ,
  \958(265) ,
  \1410(279) ,
  \441(675) ,
  \1320(254) ,
  \437(688) ,
  \1349(567) ,
  \318(113) ,
  \5(837) ,
  \1309(367) ,
  \1281(318) ,
  \382(120) ,
  \1249(338) ,
  \535(697) ,
  \1169(356) ,
  \1669(256) ,
  \1247(291) ,
  \1243(527) ,
  \68(904) ,
  \40(805) ,
  \459(200) ,
  \1093(495) ,
  \1231(379) ,
  \1038(325) ,
  \1271(349) ,
  \1594(68) ,
  \572(737) ,
  \588B(740) ,
  \1210(284) ,
  \272(414) ,
  \326(582) ,
  \191(67) ,
  \1521(786) ,
  \1045(382) ,
  \26(830) ,
  \1378(630) ,
  \1600(136) ,
  \1300(135) ,
  \1820(250) ,
  \1294(465) ,
  \1924(651) ,
  \416(660) ,
  \1343(532) ,
  \1801(493) ,
  \1153(681) ,
  \47(823) ,
  \365(585) ,
  \1769(478) ,
  \1642(183) ,
  \1202(359) ,
  \1737(469) ,
  \1237(462) ,
  \784(752) ,
  \1132(586) ,
  \254(172) ,
  \820(769) ,
  \1877(215) ,
  \1340(498) ,
  \376(910) ,
  \287(876) ,
  \1925(841) ,
  \420(668) ,
  \1073(366) ,
  \1660(331) ,
  \1592(139) ,
  \1104(302) ,
  \1338(223) ,
  \1753(131) ,
  \816(768) ,
  \547(619) ,
  \1509(758) ,
  \1621(780) ,
  \1004(540) ,
  \1365(603) ,
  \389(427) ,
  \321(144) ,
  \1(818) ,
  \1273(372) ,
  \1742(224) ,
  \379(575) ,
  \257(422) ,
  \1090(196) ,
  \29(829) ,
  \1710(212) ,
  \926(42) ,
  \1633(802) ,
  \59(898) ,
  \280(569) ,
  \1764(536) ,
  \8(836) ,
  \1311(404) ,
  \1472(190) ,
  \1345(551) ,
  \1836(203) ,
  \22(811) ,
  \1434(275) ,
  \875(744) ,
  \1581(775) ,
  \989(417) ,
  \1505(598) ,
  \168(79) ,
  \423(663) ,
  \1849(147) ,
  \1103(345) ,
  \990(262) ,
  \1900(512) ,
  \43(804) ,
  \1648(868) ,
  \265(479) ,
  \1154(193) ,
  \615(272) ,
  \1662(259) ,
  \1053(149) ,
  \556(601) ,
  \983(357) ,
  \1921(821) ,
  \487(197) ,
  \198(63) ,
  \1283(352) ,
  \1465(695) ,
  \64(96) ,
  \1317(347) ,
  \385(128) ,
  \1860(247) ,
  \415(611) ,
  \1685(525) ,
  \859(39) ,
  \1248(278) ,
  \1175(398) ,
  \340(484) ,
  \430(885) ,
  \1821(240) ,
  \1765(500) ,
  \947(34) ,
  \1287(380) ,
  \860(794) ,
  \853(97) ,
  \541(50) ,
  \70(892) ,
  \1204(207) ,
  \672(716) ,
  \262(458) ,
  \561(635) ,
  \922(43) ,
  \1554(78) ,
  \1741(489) ,
  \1152(874) ,
  \1798(448) ,
  \1725(209) ,
  \622(733) ,
  \639B(735) ,
  \1497(597) ,
  \401(583) ,
  \4(817) ,
  \1713(118) ,
  \1034(319) ,
  \399(547) ,
  \1624(125) ,
  \[10] ,
  \1133(606) ,
  \1424(340) ,
  \511(642) ,
  \372(360) ,
  \[11] ,
  \1481(613) ,
  \[12] ,
  \955(102) ,
  \[13] ,
  \1613(779) ,
  \978(180) ,
  \[14] ,
  \1545(789) ,
  \1796(296) ,
  \[15] ,
  \194(65) ,
  \404(273) ,
  \396(383) ,
  \25(810) ,
  \[16] ,
  \938(36) ,
  \495(708) ,
  \1774(624) ,
  \[17] ,
  \1845(237) ,
  \433(687) ,
  \[18] ,
  \1797(253) ,
  \1716(289) ,
  \426(888) ,
  \1003(519) ,
  \[19] ,
  \46(803) ,
  \943(35) ,
  \540(717) ,
  \1351(590) ,
  \559(600) ,
  \1105(373) ,
  \1087(553) ,
  \588A(739) ,
  \1601(798) ,
  \1705(154) ,
  \1886(455) ,
  \1048(326) ,
  \1520(174) ,
  \885(749) ,
  \780(751) ,
  \1162(267) ,
  \1593(797) ,
  \1212(363) ,
  \719(652) ,
  \1360(522) ,
  \1652(184) ,
  \1188(529) ,
  \675(725) ,
  \776(750) ,
  \360(444) ,
  \[20] ,
  \1697(153) ,
  \1917(842) ,
  \696(726) ,
  \[21] ,
  \988(333) ,
  \335(449) ,
  \557(618) ,
  \505(199) ,
  \286(884) ,
  \1692(647) ,
  \1916(650) ,
  \[22] ,
  \618(722) ,
  \1457(702) ,
  \1905(486) ,
  \1033(353) ,
  \886(782) ,
  \1014(541) ,
  \1259(348) ,
  \[23] ,
  \1482(106) ,
  \[24] ,
  \1729(468) ,
  \28(809) ,
  \1693(602) ,
  \522(719) ,
  \391(504) ,
  \1076(310) ,
  \1316(321) ,
  \512(661) ,
  \366(605) ,
  \7(816) ,
  \268(350) ,
  \1230(260) ,
  \1252(229) ,
  \934(37) ,
  \812(767) ,
  \1745(130) ,
  \553(49) ,
  \1121(403) ,
  \1009(571) ,
  \1078(195) ,
  \967(182) ,
  \1216(879) ,
  \999(418) ,
  \363(344) ,
  \422(680) ,
  \808(766) ,
  \1881(142) ,
  \1625(801) ,
  \1127(576) ,
  \71(905) ,
  \1339(198) ,
  \1897(485) ,
  \498(707) ,
  \1514(88) ,
  \1541(762) ,
  \1513(785) ,
  \1862(428) ,
  \1356(535) ,
  \1023(659) ,
  \496(714) ,
  \1544(162) ,
  \993(358) ,
  \160(83) ,
  \1829(463) ,
  \871(742) ,
  \639(724) ,
  \1573(774) ,
  \1913(822) ,
  \1286(257) ,
  \1234(440) ,
  \1425(700) ,
  \1088(545) ,
  \1426(274) ,
  \1067(393) ,
  \1373(443) ,
  \1062(285) ,
  \1665(169) ,
  \1561(791) ,
  \1806(848) ,
  \1884(244) ,
  \1837(214) ,
  \1376(664) ,
  \417(641) ,
  \1389(592) ,
  \856(98) ,
  \1634(99) ,
  \1654(258) ,
  \1616(129) ,
  \336(467) ,
  \867(736) ,
  \1276(288) ,
  \985(384) ,
  \405(304) ,
  \58(94) ,
  \1122(508) ,
  \525(718) ,
  \1137(559) ,
  \1142(531) ,
  \1095(539) ,
  \1677(524) ,
  \1416(339) ,
  \1809(610) ,
  \418(671) ,
  \377(542) ,
  \1756(306) ,
  \367(623) ,
  \1086(269) ,
  \11(835) ,
  \429(878) ,
  \1734(235) ,
  \406(335) ,
  \1873(124) ,
  \930(41) ,
  \1197(176) ,
  \278(589) ,
  \1005(555) ,
  \1239(505) ,
  \1480(187) ,
  \285(628) ,
  \1813(629) ,
  \1733(488) ,
  \1717(208) ,
  \1854(158) ,
  \407(474) ,
  \32(828) ,
  \1584(143) ,
  \1312(166) ,
  \1870(141) ,
  \295(437) ,
  \1024(640) ,
  \1044(320) ,
  \1562(76) ,
  \1889(464) ,
  \1277(401) ,
  \1157(355) ,
  \260(421) ,
  \520(706) ,
  \1709(243) ,
  \1512(178) ,
  \327(137) ,
  \1201(263) ,
  \1568(152) ,
  \1409(622) ,
  \857(784) ,
  \1165(423) ,
  \1766(515) ,
  \1910(631) ,
  \1192(399) ,
  \1537(788) ,
  \499(713) ,
  \424(644) ,
  \1605(778) ,
  \1474(105) ,
  \392(526) ,
  \1110(405) ,
  \614(271) ,
  \233(57) ,
  \836(773) ,
  \1138(544) ,
  \324(546) ,
  \1804(466) ,
  \1597(777) ,
  \1789(252) ,
  \1013(520) ,
  \1043(354) ,
  \1578(72) ,
  \1143(594) ,
  \306(433) ,
  \998(334) ,
  \528(723) ,
  \1909(511) ,
  \907(48) ,
  \1322(361) ,
  \425(674) ,
  \956(181) ,
  \188(69) ,
  \346(587) ,
  \296(454) ,
  \1397(564) ,
  \1081(494) ,
  \881(747) ,
  \1602(66) ,
  \305(409) ,
  \1293(476) ,
  \1183(218) ,
  \1585(796) ,
  \1327(528) ,
  \1830(116) ,
  \1702(246) ,
  \1788(294) ,
  \65(895) ,
  \688(727) ,
  \325(562) ,
  \1865(439) ,
  \1761(477) ,
  \517(52) ,
  \500(720) ,
  \14(834) ,
  \639A(734) ,
  \1408(870) ,
  \588(729) ,
  \1254(376) ,
  \1449(701) ,
  \1661(255) ,
  \288(160) ,
  \1226(327) ,
  \621(732) ,
  \1565(765) ,
  \364(565) ,
  \1381(392) ,
  \1348(521) ,
  \1058(230) ,
  \537(709) ,
  \359(424) ,
  \1303(292) ,
  \1618(62) ,
  \314(471) ,
  \35(827) ,
  \398(438) ,
  \1536(167) ,
  \1790(217) ,
  \1147(658) ,
  \1315(312) ,
  \50(91) ,
  \1369(621) ,
  \746(678) ,
  \1506(90) ,
  \1233(420) ,
  \1019(572) ,
  \1812(873) ,
  \1876(232) ,
  \877(745) ,
  \1299(506) ,
  \1077(394) ,
  \206(59) ,
  \1008(434) ,
  \503(731) ,
  \149(89) ,
  \1857(151) ,
  \1109(402) ,
  \1653(890) ,
  \984(329) ,
  \1305(343) ,
  \1637(839) ,
  \298(328) ,
  \307(452) ,
  \1260(298) ,
  \1793(165) ,
  \954(101) ,
  \1617(800) ,
  \1684(497) ,
  \1893(482) ,
  \1384(649) ,
  \1020(844) ,
  \1533(761) ,
  \1694(245) ,
  \309(432) ,
  \1442(109) ,
  \1708(323) ,
  \352(112) ,
  \1261(371) ,
  \1841(146) ,
  \1456(192) ,
  \1290(115) ,
  \722(653) ,
  \1437(616) ,
  \179(73) ,
  \1522(86) ,
  \560(617) ,
  \1828(450) ,
  \1094(518) ,
  \995(385) ,
  \1072(286) ,
  \308(408) ,
  \1148(639) ,
  \1402(845) ,
  \545(638) ,
  \10(815) ,
  \1298(201) ,
  \1268(211) ,
  \1289(419) ,
  \184(71) ,
  \1370(646) ,
  \1553(790) ,
  \725(665) ,
  \1657(168) ,
  \1112(228) ,
  \31(808) ,
  \523(705) ,
  \1576(148) ,
  \804(757) ,
  \1453(694) ,
  \302(122) ,
  \1163(397) ,
  \1176(145) ,
  \374(364) ,
  \1724(290) ,
  \1308(226) ,
  \1179(127) ,
  \1538(82) ,
  \17(833) ,
  \1331(549) ,
  \1066(309) ,
  \1498(104) ,
  \1222(173) ,
  \350(875) ,
  \378(557) ,
  \1678(473) ,
  \1740(314) ,
  \334(430) ,
  \919(44) ,
  \245(56) ,
  \1878(155) ,
  \38(826) ,
  \1015(556) ,
  \1726(234) ,
  \1570(74) ,
  \1805(516) ,
  \1217(897) ,
  \1441(634) ,
  \333(406) ,
  \1211(264) ,
  \1852(301) ,
  \279(609) ;
assign
  \175(75)  = ~\122(7) ,
  \457(205)  = \955(102)  & \210(16) ,
  \1485(596)  = \445(578) ,
  \529(51)  = ~\472(25) ,
  \521(712)  = ~\1457(702)  | ~\1450(110) ,
  \728(666)  = \549(655) ,
  \355(126)  = \198(63) ,
  \1244(138)  = \188(69) ,
  \400(563)  = ~\1331(549)  | ~\1322(361) ,
  \828(771)  = ~\969(266)  | (~\756(677)  | (~\688(727)  | (~\639B(735)  | ~\573(738) ))),
  \710(728)  = \672(716)  & \666(685) ,
  \202(61)  = ~\143(14) ,
  \1266(395)  = ~\1264(287)  | ~\1261(371) ,
  \949(33)  = ~\953(32) ,
  \1394(846)  = \462(820)  & (\911(46)  & \478(27) ),
  \428(886)  = ~\1400(871)  | ~\1397(564) ,
  \1325(481)  = ~\1892(475)  | ~\1889(464) ,
  \1355(533)  = ~\1908(513)  | ~\1905(486) ,
  \74(843)  = \887(819)  & (\952(31)  & (\867(736)  & \949(33) )),
  \1039(412)  = ~\1035(381) ,
  \1189(550)  = ~\1188(529)  | ~\1187(507) ,
  \66(903)  = \[21] ,
  \796(755)  = ~\958(265)  | (~\746(678)  | (~\696(726)  | (~\622(733)  | ~\588B(740) ))),
  \1758(514)  = \343(492) ,
  \546(656)  = ~\545(638)  | ~\544(620) ,
  \1304(311)  = ~\1877(215)  | ~\1870(141) ,
  \832(772)  = ~\969(266)  | (~\770(679)  | (~\696(726)  | (~\639B(735)  | ~\588B(740) ))),
  \1529(787)  = ~\1525(760) ,
  \1418(280)  = \492(204) ,
  \349(883)  = ~\1152(874)  | ~\1149(669) ,
  \1030(248)  = \288(160) ,
  \449(560)  = ~\918(45)  | ~\393(548) ,
  \361(297)  = ~\1182(236)  | ~\1179(127) ,
  \1748(305)  = ~\1742(224) ,
  \330(134)  = \191(67) ,
  \241(54)  = ~\237(23) ,
  \1421(692)  = \433(687) ,
  \548(637)  = ~\1481(613)  | ~\1474(105) ,
  \1589(776)  = \969(266)  & (\756(677)  & (\696(726)  & (\639B(735)  & \573(738) ))),
  \273(436)  = ~\1039(412)  | ~\1030(248) ,
  \1352(499)  = \407(474) ,
  \1868(447)  = ~\1862(428) ,
  \13(814)  = ~\1544(162)  | ~\1541(762) ,
  \1362(627)  = \282(608) ,
  \1610(64)  = \140(13) ,
  \564(654)  = ~\558(636) ,
  \1116(303)  = ~\1757(222)  | ~\1750(225) ,
  \865(793)  = \836(773)  & (\832(772)  & (\828(771)  & (\824(770)  & (\820(769)  & (\816(768)  & (\812(767)  & \808(766) )))))),
  \1215(887)  = ~\1812(873)  | ~\1809(610) ,
  \1170(295)  = ~\1797(253)  | ~\1790(217) ,
  \369(117)  = \938(36)  & (\241(54)  & \210(16) ),
  \994(330)  = ~\1669(256)  | ~\1662(259) ,
  \34(807)  = ~\1600(136)  | ~\1597(777) ,
  \1068(231)  = \299(140) ,
  \258(442)  = ~\999(418)  | ~\990(262) ,
  \482(202)  = ~\955(102)  | ~\214(17) ,
  \1253(362)  = ~\1249(338) ,
  \1833(123)  = \202(61) ,
  \1089(561)  = ~\1087(553)  | ~\1078(195) ,
  \1629(781)  = \969(266)  & (\756(677)  & (\710(728)  & (\639B(735)  & \588B(740) ))),
  \1668(332)  = ~\1662(259) ,
  \1255(407)  = ~\1253(362)  | ~\1244(138) ,
  \347(607)  = ~\1143(594)  | ~\1134(509) ,
  \1357(552)  = ~\1356(535)  | ~\1355(533) ,
  \281(588)  = ~\1009(571)  | ~\1000(410) ,
  \62(95)  = ~\947(34)  | ~\930(41) ,
  \1608(133)  = ~\1602(66) ,
  \566(277)  = \482(202) ,
  \274(453)  = ~\273(436)  | ~\272(414) ,
  \1050(163)  = \160(83) ,
  \1504(186)  = ~\1498(104) ,
  \1171(369)  = ~\1170(295)  | ~\1169(356) ,
  \1018(435)  = ~\1010(411) ,
  \1417(699)  = ~\1413(691) ,
  \1466(108)  = \529(51) ,
  \1120(308)  = ~\1112(228) ,
  \1822(431)  = ~\1255(407)  | ~\1254(376) ,
  \756(677)  = \728(666)  & \719(652) ,
  \1718(213)  = \302(122) ,
  \1429(615)  = \453(599) ,
  \410(470)  = \310(451) ,
  \1557(764)  = \958(265)  & (\731(676)  & (\710(728)  & (\622(733)  & \588B(740) ))),
  \1586(70)  = \131(10) ,
  \61(896)  = ~\429(878)  | ~\428(886) ,
  \1496(185)  = ~\1490(103) ,
  \1278(170)  = \156(85) ,
  \524(711)  = ~\1449(701)  | ~\1442(109) ,
  \1029(682)  = ~\1025(670) ,
  \21(859)  = \[9] ,
  \348(625)  = ~\347(607)  | ~\346(587) ,
  \1193(566)  = ~\1189(550) ,
  \171(77)  = ~\119(6) ,
  \373(283)  = ~\1211(264)  | ~\1204(207) ,
  \1782(216)  = \355(126) ,
  \1166(194)  = \352(112) ,
  \343(492)  = \314(471) ,
  \1908(513)  = ~\1902(491) ,
  \1225(317)  = ~\1820(250)  | ~\1817(150) ,
  \873(743)  = ~\979(179)  | (~\731(676)  | (~\675(725)  | (~\639B(735)  | ~\573(738) ))),
  \1326(523)  = ~\1893(482)  | ~\1886(455) ,
  \1242(457)  = ~\1234(440) ,
  \277(570)  = ~\1018(435)  | ~\1015(556) ,
  \1220(391)  = ~\1212(363) ,
  \1440(337)  = ~\1434(275) ,
  \1144(849)  = \462(820)  & (\911(46)  & \469(24) ),
  \1164(388)  = ~\1162(267)  | ~\1159(368) ,
  \1282(324)  = ~\1861(241)  | ~\1854(158) ,
  \862(38)  = ~\953(32) ,
  \1780(645)  = ~\1774(624) ,
  \1577(795)  = ~\1573(774) ,
  \1115(346)  = ~\1756(306)  | ~\1753(131) ,
  \1681(503)  = \265(479) ,
  \1530(84)  = \110(3) ,
  \573(738)  = \569(730)  & \566(277) ,
  \1344(534)  = ~\1901(510)  | ~\1894(490) ,
  \69(908)  = \[22] ,
  \533(704)  = ~\1473(696)  | ~\1466(108) ,
  \1056(251)  = ~\1050(163) ,
  \1785(164)  = \160(83) ,
  \1525(760)  = \958(265)  & (\746(678)  & (\675(725)  & (\639A(734)  & \588A(739) ))),
  \1894(490)  = \410(470) ,
  \1686(626)  = \282(608) ,
  \16(813)  = ~\1552(159)  | ~\1549(763) ,
  \1676(496)  = ~\1670(472) ,
  \1626(60)  = \146(15) ,
  \1892(475)  = ~\1886(455) ,
  \1902(491)  = \410(470) ,
  \248(55)  = \234(22) ,
  \1448(191)  = ~\1442(109) ,
  \1643(889)  = ~\1639(881) ,
  \42(852)  = \[15] ,
  \663(684)  = ~\513(672) ,
  \911(46)  = \902(30) ,
  \37(806)  = ~\1608(133)  | ~\1605(778) ,
  \1207(177)  = \149(89) ,
  \1477(595)  = \445(578) ,
  \1814(161)  = \165(81) ,
  \1264(287)  = ~\1256(210) ,
  \1361(568)  = ~\1357(552) ,
  \1393(612)  = ~\1389(592) ,
  \1493(579)  = \449(560) ,
  \1560(156)  = ~\1554(78) ,
  \[0]  = ~\2(838)  | ~\1(818) ,
  \1401(584)  = ~\1397(564) ,
  \1385(425)  = ~\1381(392) ,
  \1000(410)  = \269(378) ,
  \1757(222)  = ~\1753(131) ,
  \800(756)  = ~\958(265)  | (~\731(676)  | (~\710(728)  | (~\622(733)  | ~\588B(740) ))),
  \1111(429)  = ~\1109(402)  | ~\1100(227) ,
  \[1]  = ~\5(837)  | ~\4(817) ,
  \1489(614)  = ~\1485(596) ,
  \[2]  = ~\8(836)  | ~\7(816) ,
  \569(730)  = ~\500(720) ,
  \1232(387)  = ~\1230(260)  | ~\1227(351) ,
  \1194(206)  = \369(117) ,
  \[3]  = ~\11(835)  | ~\10(815) ,
  \1125(558)  = ~\1764(536)  | ~\1761(477) ,
  \1028(869)  = ~\1020(844) ,
  \1130(530)  = ~\1122(508) ,
  \1377(460)  = ~\1373(443) ,
  \549(655)  = ~\548(637)  | ~\547(619) ,
  \294(415)  = ~\1048(326)  | ~\1045(382) ,
  \[4]  = ~\29(829)  | ~\28(809) ,
  \1445(693)  = \437(688) ,
  \1061(341)  = ~\1716(289)  | ~\1713(118) ,
  \55(911)  = ~\376(910)  | ~\375(906) ,
  \[5]  = ~\44(824)  | ~\43(804) ,
  \1083(538)  = ~\1082(517)  | ~\1081(494) ,
  \[6]  = ~\47(823)  | ~\46(803) ,
  \1817(150)  = \175(75) ,
  \[7]  = ~\14(834)  | ~\13(814) ,
  \362(315)  = ~\1183(218)  | ~\1176(145) ,
  \863(783)  = \804(757)  & (\800(756)  & (\796(755)  & (\792(754)  & (\788(753)  & (\784(752)  & (\780(751)  & \776(750) )))))),
  \1639(881)  = ~\1638(867)  | ~\1637(839) ,
  \3(865)  = \[0] ,
  \1049(413)  = ~\1045(382) ,
  \1099(554)  = ~\1095(539) ,
  \[8]  = ~\17(833)  | ~\16(813) ,
  \24(858)  = \[10] ,
  \1647(840)  = ~\1924(651)  | ~\1921(821) ,
  \1777(461)  = ~\360(444) ,
  \445(578)  = ~\918(45)  | ~\379(575) ,
  \[9]  = ~\20(832)  | ~\19(812) ,
  \1501(580)  = \449(560) ,
  \1117(374)  = ~\1116(303)  | ~\1115(346) ,
  \1040(249)  = \288(160) ,
  \1464(189)  = ~\1458(107) ,
  \1701(242)  = ~\1697(153) ,
  \1732(313)  = ~\1726(234) ,
  \558(636)  = ~\557(618)  | ~\556(601) ,
  \1057(239)  = ~\1053(149) ,
  \1025(670)  = ~\1024(640)  | ~\1023(659) ,
  \1528(171)  = ~\1522(86) ,
  \1609(799)  = ~\1605(778) ,
  \1433(633)  = ~\1429(615) ,
  \510(673)  = ~\509(662)  | ~\508(643) ,
  \413(574)  = ~\1360(522)  | ~\1357(552) ,
  \1174(268)  = ~\1166(194) ,
  \824(770)  = ~\969(266)  | (~\731(676)  | (~\710(728)  | (~\639B(735)  | ~\573(738) ))),
  \310(451)  = ~\309(432)  | ~\308(408) ,
  \45(851)  = \[5] ,
  \1450(110)  = \517(52) ,
  \792(754)  = ~\958(265)  | (~\756(677)  | (~\696(726)  | (~\622(733)  | ~\588A(739) ))),
  \1035(381)  = ~\1034(319)  | ~\1033(353) ,
  \536(703)  = ~\1465(695)  | ~\1458(107) ,
  \1265(400)  = ~\1261(371) ,
  \421(657)  = ~\1377(460)  | ~\1370(646) ,
  \731(676)  = \725(665)  & \719(652) ,
  \153(87)  = ~\104(1) ,
  \244(53)  = ~\237(23) ,
  \492(204)  = ~\955(102)  | ~\210(16) ,
  \1546(80)  = \116(5) ,
  \1221(907)  = ~\1217(897) ,
  \1689(581)  = ~\1089(561)  | ~\1088(545) ,
  \1126(543)  = ~\1765(500)  | ~\1758(514) ,
  \1386(847)  = \462(820)  & (\911(46)  & \475(26) ),
  \67(891)  = ~\1642(183)  | ~\1639(881) ,
  \390(446)  = ~\389(427)  | ~\388(396) ,
  \1901(510)  = ~\1897(485) ,
  \883(748)  = ~\979(179)  | (~\731(676)  | (~\675(725)  | (~\621(732)  | ~\573(738) ))),
  \932(40)  = ~\952(31) ,
  \19(812)  = ~\1560(156)  | ~\1557(764) ,
  \918(45)  = ~\902(30) ,
  \1321(377)  = ~\1317(347) ,
  \770(679)  = \728(666)  & \722(653) ,
  \666(685)  = \513(672) ,
  \41(825)  = ~\1617(800)  | ~\1610(64) ,
  \1461(689)  = \441(675) ,
  \969(266)  = ~\978(180)  | ~\967(182) ,
  \788(753)  = ~\958(265)  | (~\731(676)  | (~\688(727)  | (~\639A(734)  | ~\588A(739) ))),
  \1131(593)  = ~\1127(576) ,
  \291(157)  = \168(79) ,
  \1063(365)  = ~\1062(285)  | ~\1061(341) ,
  \73(741)  = \867(736)  & (\932(40)  & \949(33) ),
  \1413(691)  = \433(687) ,
  \1267(426)  = ~\1265(400)  | ~\1256(210) ,
  \1295(483)  = ~\1294(465)  | ~\1293(476) ,
  \1200(281)  = ~\1194(206) ,
  \1517(759)  = \958(265)  & (\756(677)  & (\675(725)  & (\639A(734)  & \588A(739) ))),
  \879(746)  = ~\979(179)  | (~\746(678)  | (~\675(725)  | (~\622(733)  | ~\573(738) ))),
  \1825(445)  = ~\1267(426)  | ~\1266(395) ,
  \1861(241)  = ~\1857(151) ,
  \20(832)  = ~\1561(791)  | ~\1554(78) ,
  \259(459)  = ~\258(442)  | ~\257(422) ,
  \1227(351)  = ~\1226(327)  | ~\1225(317) ,
  \1846(220)  = \385(128) ,
  \534(710)  = ~\533(704)  | ~\532(698) ,
  \1158(293)  = ~\1789(252)  | ~\1782(216) ,
  \1182(236)  = ~\1176(145) ,
  \887(819)  = \886(782)  & (\865(793)  & \863(783) ),
  \1288(386)  = ~\1286(257)  | ~\1283(352) ,
  \269(378)  = ~\268(350) ,
  \1750(225)  = \330(134) ,
  \297(316)  = ~\1056(251)  | ~\1053(149) ,
  \1400(871)  = ~\1394(846) ,
  \427(880)  = ~\1393(612)  | ~\1386(847) ,
  \1139(577)  = ~\1138(544)  | ~\1137(559) ,
  \1772(537)  = ~\1766(515) ,
  \1392(872)  = ~\1386(847) ,
  \56(93)  = ~\947(34)  | ~\930(41) ,
  \516(686)  = ~\510(673) ,
  \1330(390)  = ~\1322(361) ,
  \53(893)  = ~\350(875)  | ~\349(883) ,
  \6(864)  = \[1] ,
  \282(608)  = ~\281(588)  | ~\280(569) ,
  \1844(299)  = ~\1838(219) ,
  \508(643)  = ~\1440(337)  | ~\1437(616) ,
  \49(894)  = ~\287(876)  | ~\286(884) ,
  \27(857)  = \[11] ,
  \909(47)  = ~\900(29) ,
  \1549(763)  = \958(265)  & (\746(678)  & (\696(726)  & (\622(733)  & \588B(740) ))),
  \1159(368)  = ~\1158(293)  | ~\1157(355) ,
  \1458(107)  = \529(51) ,
  \513(672)  = ~\512(661)  | ~\511(642) ,
  \1310(375)  = ~\1308(226)  | ~\1305(343) ,
  \1108(307)  = ~\1100(227) ,
  \1350(573)  = ~\1348(521)  | ~\1345(551) ,
  \2(838)  = ~\1513(785)  | ~\1506(90) ,
  \1781(480)  = ~\1777(461) ,
  \414(591)  = ~\1361(568)  | ~\1352(499) ,
  \532(698)  = ~\1472(190)  | ~\1469(690) ,
  \1644(100)  = \934(37)  & \233(57) ,
  \48(850)  = \[6] ,
  \358(389)  = ~\1174(268)  | ~\1171(369) ,
  \669(715)  = ~\537(709) ,
  \388(396)  = ~\1276(288)  | ~\1273(372) ,
  \1238(487)  = ~\1829(463)  | ~\1822(431) ,
  \1187(507)  = ~\1804(466)  | ~\1801(493) ,
  \1638(867)  = ~\1917(842)  | ~\1910(631) ,
  \397(416)  = ~\1321(377)  | ~\1312(166) ,
  \1869(456)  = ~\1865(439) ,
  \979(179)  = \893(111)  & (\949(33)  & \926(42) ),
  \1700(322)  = ~\1694(245) ,
  \23(831)  = ~\1569(792)  | ~\1562(76) ,
  \1569(792)  = ~\1565(765) ,
  \1773(501)  = ~\1769(478) ,
  \1335(114)  = \938(36)  & (\245(56)  & \221(19) ),
  \1203(282)  = ~\1201(263)  | ~\1194(206) ,
  \1134(509)  = \340(484) ,
  \1432(336)  = ~\1426(274) ,
  \544(620)  = ~\1488(188)  | ~\1485(596) ,
  \375(906)  = ~\1220(391)  | ~\1217(897) ,
  \1010(411)  = \269(378) ,
  \1632(121)  = ~\1626(60) ,
  \44(824)  = ~\1625(801)  | ~\1618(62) ,
  \552(667)  = ~\546(656) ,
  \231(58)  = ~\898(28)  | ~\224(20) ,
  \165(81)  = ~\113(4) ,
  \1469(690)  = \441(675) ,
  \1673(502)  = \265(479) ,
  \1368(648)  = ~\1362(627) ,
  \1272(300)  = ~\1853(238)  | ~\1846(220) ,
  \1149(669)  = ~\1148(639)  | ~\1147(658) ,
  \497(721)  = ~\496(714)  | ~\495(708) ,
  \52(92)  = ~\947(34)  | ~\930(41) ,
  \251(175)  = \149(89) ,
  \1082(517)  = ~\1733(488)  | ~\1726(234) ,
  \299(140)  = \184(71) ,
  \1721(119)  = \206(59) ,
  \980(261)  = \251(175) ,
  \1488(188)  = ~\1482(106) ,
  \261(441)  = ~\989(417)  | ~\980(261) ,
  \1749(221)  = ~\1745(130) ,
  \431(877)  = ~\1409(622)  | ~\1402(845) ,
  \893(111)  = ~\237(23)  | ~\248(55) ,
  \1918(632)  = \367(623)  & \856(98) ,
  \565(276)  = ~\482(202) ,
  \453(599)  = ~\918(45)  | ~\401(583) ,
  \393(548)  = ~\392(526)  | ~\391(504) ,
  \1100(227)  = \327(137) ,
  \462(820)  = ~\865(793)  | ~\863(783) ,
  \1256(210)  = \382(120) ,
  \1885(233)  = ~\1881(142) ,
  \1332(132)  = \194(65) ,
  \1473(696)  = ~\1469(690) ,
  \9(863)  = \[2] ,
  \509(662)  = ~\1441(634)  | ~\1434(275) ,
  \1184(370)  = ~\363(344) ,
  \1098(270)  = ~\1090(196) ,
  \1838(219)  = \385(128) ,
  \1853(238)  = ~\1849(147) ,
  \1490(103)  = \553(49) ,
  \1649(882)  = ~\1648(868)  | ~\1647(840) ,
  \1670(472)  = \274(453) ,
  \419(683)  = ~\418(671) ,
  \1071(342)  = ~\1724(290)  | ~\1721(119) ,
  \1405(604)  = \401(583) ,
  \1552(159)  = ~\1546(80) ,
  \156(85)  = ~\107(2) ,
  \958(265)  = ~\978(180)  | ~\956(181) ,
  \1410(279)  = \492(204) ,
  \441(675)  = ~\918(45)  | ~\425(674) ,
  \1320(254)  = ~\1312(166) ,
  \437(688)  = ~\918(45)  | ~\422(680) ,
  \1349(567)  = ~\1345(551) ,
  \318(113)  = \938(36)  & \224(20) ,
  \5(837)  = ~\1521(786)  | ~\1514(88) ,
  \1309(367)  = ~\1305(343) ,
  \1281(318)  = ~\1860(247)  | ~\1857(151) ,
  \382(120)  = \206(59) ,
  \1249(338)  = ~\1248(278)  | ~\1247(291) ,
  \535(697)  = ~\1464(189)  | ~\1461(689) ,
  \1169(356)  = ~\1796(296)  | ~\1793(165) ,
  \1669(256)  = ~\1665(169) ,
  \1247(291)  = ~\1836(203)  | ~\1833(123) ,
  \1243(527)  = ~\1239(505) ,
  \72(909)  = \[23] ,
  \68(904)  = ~\1643(889)  | ~\1634(99) ,
  \40(805)  = ~\1616(129)  | ~\1613(779) ,
  \459(200)  = \954(101)  & \217(18) ,
  \1093(495)  = ~\1740(314)  | ~\1737(469) ,
  \1231(379)  = ~\1227(351) ,
  \1038(325)  = ~\1030(248) ,
  \1271(349)  = ~\1852(301)  | ~\1849(147) ,
  \54(900)  = \[18] ,
  \1594(68)  = \134(11) ,
  \572(737)  = \569(730)  & \565(276) ,
  \588B(740)  = \588(729) ,
  \1210(284)  = ~\1204(207) ,
  \272(414)  = ~\1038(325)  | ~\1035(381) ,
  \326(582)  = ~\325(562)  | ~\324(546) ,
  \191(67)  = ~\134(11) ,
  \1521(786)  = ~\1517(759) ,
  \1045(382)  = ~\1044(320)  | ~\1043(354) ,
  \26(830)  = ~\1577(795)  | ~\1570(74) ,
  \1378(630)  = ~\415(611) ,
  \1600(136)  = ~\1594(68) ,
  \1300(135)  = \191(67) ,
  \1820(250)  = ~\1814(161) ,
  \1294(465)  = ~\1869(456)  | ~\1862(428) ,
  \1924(651)  = ~\1918(632) ,
  \416(660)  = ~\1368(648)  | ~\1365(603) ,
  \1343(532)  = ~\1900(512)  | ~\1897(485) ,
  \1801(493)  = \314(471) ,
  \1153(681)  = ~\1149(669) ,
  \47(823)  = ~\1633(802)  | ~\1626(60) ,
  \365(585)  = ~\1193(566)  | ~\1184(370) ,
  \1769(478)  = \262(458) ,
  \1642(183)  = ~\1634(99) ,
  \1202(359)  = ~\1200(281)  | ~\1197(176) ,
  \1737(469)  = \310(451) ,
  \1237(462)  = ~\1828(450)  | ~\1825(445) ,
  \784(752)  = ~\958(265)  | (~\746(678)  | (~\675(725)  | (~\639A(734)  | ~\588A(739) ))),
  \1132(586)  = ~\1130(530)  | ~\1127(576) ,
  \254(172)  = \153(87) ,
  \820(769)  = ~\969(266)  | (~\746(678)  | (~\696(726)  | (~\639B(735)  | ~\573(738) ))),
  \1877(215)  = ~\1873(124) ,
  \1340(498)  = \407(474) ,
  \376(910)  = ~\1221(907)  | ~\1212(363) ,
  \287(876)  = ~\1029(682)  | ~\1020(844) ,
  \1925(841)  = ~\1921(821) ,
  \420(668)  = ~\1376(664)  | ~\1373(443) ,
  \1073(366)  = ~\1072(286)  | ~\1071(342) ,
  \1660(331)  = ~\1654(258) ,
  \1592(139)  = ~\1586(70) ,
  \1104(302)  = ~\1749(221)  | ~\1742(224) ,
  \1338(223)  = ~\1332(132) ,
  \1753(131)  = \194(65) ,
  \816(768)  = ~\969(266)  | (~\756(677)  | (~\696(726)  | (~\639B(735)  | ~\573(738) ))),
  \547(619)  = ~\1480(187)  | ~\1477(595) ,
  \1509(758)  = \958(265)  & (\731(676)  & (\696(726)  & (\639A(734)  & \588A(739) ))),
  \1621(780)  = \969(266)  & (\770(679)  & (\696(726)  & (\639B(735)  & \588B(740) ))),
  \1004(540)  = ~\1677(524)  | ~\1670(472) ,
  \1365(603)  = ~\326(582) ,
  \389(427)  = ~\1277(401)  | ~\1268(211) ,
  \321(144)  = \179(73) ,
  \1(818)  = ~\1512(178)  | ~\1509(758) ,
  \1273(372)  = ~\1272(300)  | ~\1271(349) ,
  \1742(224)  = \330(134) ,
  \379(575)  = ~\378(557)  | ~\377(542) ,
  \257(422)  = ~\998(334)  | ~\995(385) ,
  \1090(196)  = \318(113) ,
  \29(829)  = ~\1585(796)  | ~\1578(72) ,
  \1710(212)  = \302(122) ,
  \926(42)  = \952(31) ,
  \1633(802)  = ~\1629(781) ,
  \59(898)  = ~\427(880)  | ~\426(888) ,
  \280(569)  = ~\1008(434)  | ~\1005(555) ,
  \1764(536)  = ~\1758(514) ,
  \8(836)  = ~\1529(787)  | ~\1522(86) ,
  \1311(404)  = ~\1309(367)  | ~\1300(135) ,
  \1472(190)  = ~\1466(108) ,
  \1345(551)  = ~\1344(534)  | ~\1343(532) ,
  \1836(203)  = ~\1830(116) ,
  \22(811)  = ~\1568(152)  | ~\1565(765) ,
  \1434(275)  = \505(199) ,
  \875(744)  = ~\979(179)  | (~\731(676)  | (~\696(726)  | (~\622(733)  | ~\573(738) ))),
  \1581(775)  = \969(266)  & (\746(678)  & (\710(728)  & (\639A(734)  & \588B(740) ))),
  \989(417)  = ~\985(384) ,
  \1505(598)  = ~\1501(580) ,
  \168(79)  = ~\116(5) ,
  \423(663)  = ~\1384(649)  | ~\1381(392) ,
  \1849(147)  = \179(73) ,
  \1103(345)  = ~\1748(305)  | ~\1745(130) ,
  \990(262)  = \251(175) ,
  \1900(512)  = ~\1894(490) ,
  \43(804)  = ~\1624(125)  | ~\1621(780) ,
  \1648(868)  = ~\1925(841)  | ~\1918(632) ,
  \265(479)  = ~\259(459) ,
  \1154(193)  = \352(112) ,
  \615(272)  = \487(197) ,
  \1662(259)  = \254(172) ,
  \1053(149)  = \175(75) ,
  \556(601)  = ~\1504(186)  | ~\1501(580) ,
  \983(357)  = ~\1660(331)  | ~\1657(168) ,
  \1921(821)  = \862(38)  & \860(794) ,
  \487(197)  = ~\954(101)  | ~\221(19) ,
  \198(63)  = ~\140(13) ,
  \1283(352)  = ~\1282(324)  | ~\1281(318) ,
  \1465(695)  = ~\1461(689) ,
  \64(96)  = ~\947(34)  | ~\930(41) ,
  \1317(347)  = ~\1316(321)  | ~\1315(312) ,
  \385(128)  = \198(63) ,
  \1860(247)  = ~\1854(158) ,
  \415(611)  = ~\414(591)  | ~\413(574) ,
  \1685(525)  = ~\1681(503) ,
  \859(39)  = ~\953(32) ,
  \1248(278)  = ~\1837(214)  | ~\1830(116) ,
  \1175(398)  = ~\1171(369) ,
  \340(484)  = \336(467) ,
  \430(885)  = ~\1408(870)  | ~\1405(604) ,
  \1821(240)  = ~\1817(150) ,
  \1765(500)  = ~\1761(477) ,
  \947(34)  = \953(32) ,
  \1287(380)  = ~\1283(352) ,
  \860(794)  = ~\836(773)  | (~\832(772)  | (~\828(771)  | (~\824(770)  | (~\820(769)  | (~\816(768)  | (~\812(767)  | ~\808(766) )))))),
  \853(97)  = ~\907(48)  | ~\943(35) ,
  \541(50)  = ~\475(26) ,
  \70(892)  = ~\1652(184)  | ~\1649(882) ,
  \1204(207)  = \369(117) ,
  \672(716)  = \537(709) ,
  \262(458)  = ~\261(441)  | ~\260(421) ,
  \561(635)  = ~\560(617)  | ~\559(600) ,
  \922(43)  = ~\902(30) ,
  \1554(78)  = \119(6) ,
  \1741(489)  = ~\1737(469) ,
  \1152(874)  = ~\1144(849) ,
  \1798(448)  = ~\1111(429)  | ~\1110(405) ,
  \1725(209)  = ~\1721(119) ,
  \622(733)  = \618(722)  & \615(272) ,
  \639B(735)  = \639(724) ,
  \1497(597)  = ~\1493(579) ,
  \401(583)  = ~\400(563)  | ~\399(547) ,
  \4(817)  = ~\1520(174)  | ~\1517(759) ,
  \1713(118)  = \206(59) ,
  \1034(319)  = ~\1701(242)  | ~\1694(245) ,
  \399(547)  = ~\1330(390)  | ~\1327(528) ,
  \1624(125)  = ~\1618(62) ,
  \[10]  = ~\23(831)  | ~\22(811) ,
  \1133(606)  = ~\1131(593)  | ~\1122(508) ,
  \1424(340)  = ~\1418(280) ,
  \511(642)  = ~\1432(336)  | ~\1429(615) ,
  \372(360)  = ~\1210(284)  | ~\1207(177) ,
  \[11]  = ~\26(830)  | ~\25(810) ,
  \1481(613)  = ~\1477(595) ,
  \[12]  = ~\32(828)  | ~\31(808) ,
  \955(102)  = ~\922(43)  | ~\244(53) ,
  \[13]  = ~\35(827)  | ~\34(807) ,
  \30(856)  = \[4] ,
  \1613(779)  = \969(266)  & (\756(677)  & (\688(727)  & (\639B(735)  & \573(738) ))),
  \978(180)  = ~\893(111)  | (~\949(33)  | ~\926(42) ),
  \[14]  = ~\38(826)  | ~\37(806) ,
  \1545(789)  = ~\1541(762) ,
  \1796(296)  = ~\1790(217) ,
  \[15]  = ~\41(825)  | ~\40(805) ,
  \194(65)  = ~\137(12) ,
  \404(273)  = ~\1338(223)  | ~\1335(114) ,
  \396(383)  = ~\1320(254)  | ~\1317(347) ,
  \25(810)  = ~\1576(148)  | ~\1573(774) ,
  \[16]  = ~\74(843)  & ~\73(741) ,
  \938(36)  = ~\953(32) ,
  \495(708)  = ~\1424(340)  | ~\1421(692) ,
  \1774(624)  = ~\1133(606)  | ~\1132(586) ,
  \[17]  = \50(91)  & \49(894) ,
  \1845(237)  = ~\1841(146) ,
  \433(687)  = ~\918(45)  | ~\419(683) ,
  \57(912)  = \[24] ,
  \[18]  = \53(893)  & \52(92) ,
  \1797(253)  = ~\1793(165) ,
  \1716(289)  = ~\1710(212) ,
  \426(888)  = ~\1392(872)  | ~\1389(592) ,
  \1003(519)  = ~\1676(496)  | ~\1673(502) ,
  \[19]  = \59(898)  & \58(94) ,
  \46(803)  = ~\1632(121)  | ~\1629(781) ,
  \943(35)  = \953(32) ,
  \540(717)  = ~\534(710) ,
  \1351(590)  = ~\1349(567)  | ~\1340(498) ,
  \559(600)  = ~\1496(185)  | ~\1493(579) ,
  \1105(373)  = ~\1104(302)  | ~\1103(345) ,
  \1087(553)  = ~\1083(538) ,
  \588A(739)  = \588(729) ,
  \1601(798)  = ~\1597(777) ,
  \1705(154)  = \171(77) ,
  \1886(455)  = ~\398(438) ,
  \1048(326)  = ~\1040(249) ,
  \1520(174)  = ~\1514(88) ,
  \885(749)  = ~\979(179)  | (~\731(676)  | (~\675(725)  | (~\622(733)  | ~\572(737) ))),
  \780(751)  = ~\958(265)  | (~\756(677)  | (~\675(725)  | (~\639A(734)  | ~\588A(739) ))),
  \1162(267)  = ~\1154(193) ,
  \1593(797)  = ~\1589(776) ,
  \1212(363)  = ~\1203(282)  | ~\1202(359) ,
  \719(652)  = ~\561(635) ,
  \1360(522)  = ~\1352(499) ,
  \1652(184)  = ~\1644(100) ,
  \1188(529)  = ~\1805(516)  | ~\1798(448) ,
  \675(725)  = \669(715)  & \663(684) ,
  \776(750)  = ~\958(265)  | (~\731(676)  | (~\696(726)  | (~\639A(734)  | ~\588A(739) ))),
  \360(444)  = ~\359(424)  | ~\358(389) ,
  \[20]  = \62(95)  & \61(896) ,
  \1697(153)  = \171(77) ,
  \1917(842)  = ~\1913(822) ,
  \696(726)  = \672(716)  & \663(684) ,
  \[21]  = \65(895)  & \64(96) ,
  \988(333)  = ~\980(261) ,
  \335(449)  = ~\334(430)  | ~\333(406) ,
  \557(618)  = ~\1505(598)  | ~\1498(104) ,
  \505(199)  = ~\954(101)  | ~\217(18) ,
  \286(884)  = ~\1028(869)  | ~\1025(670) ,
  \1692(647)  = ~\1686(626) ,
  \1916(650)  = ~\1910(631) ,
  \[22]  = ~\68(904)  | ~\67(891) ,
  \618(722)  = ~\525(718) ,
  \1457(702)  = ~\1453(694) ,
  \1905(486)  = \336(467) ,
  \1033(353)  = ~\1700(322)  | ~\1697(153) ,
  \886(782)  = \885(749)  & (\883(748)  & (\881(747)  & (\879(746)  & (\877(745)  & (\875(744)  & (\873(743)  & \871(742) )))))),
  \1014(541)  = ~\1685(525)  | ~\1678(473) ,
  \1259(348)  = ~\1844(299)  | ~\1841(146) ,
  \[23]  = ~\71(905)  | ~\70(892) ,
  \1482(106)  = \541(50) ,
  \33(855)  = \[12] ,
  \[24]  = \56(93)  & \55(911) ,
  \1729(468)  = \310(451) ,
  \28(809)  = ~\1584(143)  | ~\1581(775) ,
  \1693(602)  = ~\1689(581) ,
  \522(719)  = ~\521(712)  | ~\520(706) ,
  \391(504)  = ~\1298(201)  | ~\1295(483) ,
  \1076(310)  = ~\1068(231) ,
  \1316(321)  = ~\1885(233)  | ~\1878(155) ,
  \512(661)  = ~\1433(633)  | ~\1426(274) ,
  \366(605)  = ~\365(585)  | ~\364(565) ,
  \7(816)  = ~\1528(171)  | ~\1525(760) ,
  \268(350)  = ~\298(328)  | ~\297(316) ,
  \1230(260)  = ~\1222(173) ,
  \1252(229)  = ~\1244(138) ,
  \934(37)  = \953(32) ,
  \812(767)  = ~\969(266)  | (~\746(678)  | (~\710(728)  | (~\639A(734)  | ~\588B(740) ))),
  \12(862)  = \[3] ,
  \1745(130)  = \194(65) ,
  \553(49)  = ~\478(27) ,
  \1121(403)  = ~\1117(374) ,
  \1009(571)  = ~\1005(555) ,
  \1078(195)  = \318(113) ,
  \967(182)  = ~\893(111)  | (~\943(35)  | (~\919(44)  | ~\909(47) )),
  \1216(879)  = ~\1813(629)  | ~\1806(848) ,
  \999(418)  = ~\995(385) ,
  \363(344)  = ~\362(315)  | ~\361(297) ,
  \422(680)  = ~\421(657)  | ~\420(668) ,
  \808(766)  = ~\969(266)  | (~\756(677)  | (~\688(727)  | (~\622(733)  | ~\588B(740) ))),
  \1881(142)  = \184(71) ,
  \1625(801)  = ~\1621(780) ,
  \1127(576)  = ~\1126(543)  | ~\1125(558) ,
  \71(905)  = ~\1653(890)  | ~\1644(100) ,
  \1339(198)  = ~\1335(114) ,
  \1897(485)  = \336(467) ,
  \498(707)  = ~\1416(339)  | ~\1413(691) ,
  \1514(88)  = \104(1) ,
  \1541(762)  = \958(265)  & (\756(677)  & (\696(726)  & (\622(733)  & \588A(739) ))),
  \1513(785)  = ~\1509(758) ,
  \1862(428)  = ~\1311(404)  | ~\1310(375) ,
  \1356(535)  = ~\1909(511)  | ~\1902(491) ,
  \1023(659)  = ~\1692(647)  | ~\1689(581) ,
  \496(714)  = ~\1425(700)  | ~\1418(280) ,
  \1544(162)  = ~\1538(82) ,
  \993(358)  = ~\1668(332)  | ~\1665(169) ,
  \160(83)  = ~\110(3) ,
  \1829(463)  = ~\1825(445) ,
  \871(742)  = ~\979(179)  | (~\731(676)  | (~\675(725)  | (~\622(733)  | ~\588B(740) ))),
  \639(724)  = \525(718)  & \615(272) ,
  \1573(774)  = \969(266)  & (\756(677)  & (\688(727)  & (\622(733)  & \588B(740) ))),
  \1913(822)  = \859(39)  & \857(784) ,
  \1286(257)  = ~\1278(170) ,
  \1234(440)  = ~\1233(420)  | ~\1232(387) ,
  \1425(700)  = ~\1421(692) ,
  \1088(545)  = ~\1086(269)  | ~\1083(538) ,
  \1426(274)  = \505(199) ,
  \1067(393)  = ~\1063(365) ,
  \1373(443)  = ~\1165(423)  | ~\1164(388) ,
  \1062(285)  = ~\1717(208)  | ~\1710(212) ,
  \1665(169)  = \156(85) ,
  \1561(791)  = ~\1557(764) ,
  \1806(848)  = \462(820)  & (\911(46)  & \472(25) ),
  \1884(244)  = ~\1878(155) ,
  \1837(214)  = ~\1833(123) ,
  \1376(664)  = ~\1370(646) ,
  \417(641)  = ~\1369(621)  | ~\1362(627) ,
  \1389(592)  = \379(575) ,
  \856(98)  = ~\909(47)  | ~\943(35) ,
  \1634(99)  = \934(37)  & \231(58) ,
  \15(861)  = \[7] ,
  \1654(258)  = \254(172) ,
  \1616(129)  = ~\1610(64) ,
  \336(467)  = ~\335(449) ,
  \867(736)  = ~\487(197)  | (~\503(731)  | (~\528(723)  | (~\482(202)  | (~\540(717)  | (~\552(667)  | (~\564(654)  | ~\516(686) )))))),
  \1276(288)  = ~\1268(211) ,
  \985(384)  = ~\984(329)  | ~\983(357) ,
  \405(304)  = ~\1339(198)  | ~\1332(132) ,
  \58(94)  = ~\947(34)  | ~\930(41) ,
  \1122(508)  = \340(484) ,
  \525(718)  = ~\524(711)  | ~\523(705) ,
  \36(854)  = \[13] ,
  \1137(559)  = ~\1772(537)  | ~\1769(478) ,
  \1142(531)  = ~\1134(509) ,
  \1095(539)  = ~\1094(518)  | ~\1093(495) ,
  \1677(524)  = ~\1673(502) ,
  \1416(339)  = ~\1410(279) ,
  \1809(610)  = ~\1351(590)  | ~\1350(573) ,
  \418(671)  = ~\417(641)  | ~\416(660) ,
  \377(542)  = ~\1242(457)  | ~\1239(505) ,
  \1756(306)  = ~\1750(225) ,
  \367(623)  = ~\366(605) ,
  \1086(269)  = ~\1078(195) ,
  \11(835)  = ~\1537(788)  | ~\1530(84) ,
  \429(878)  = ~\1401(584)  | ~\1394(846) ,
  \1734(235)  = \321(144) ,
  \406(335)  = ~\405(304)  | ~\404(273) ,
  \1873(124)  = \202(61) ,
  \930(41)  = ~\952(31) ,
  \1197(176)  = \149(89) ,
  \278(589)  = ~\1019(572)  | ~\1010(411) ,
  \1005(555)  = ~\1004(540)  | ~\1003(519) ,
  \1239(505)  = ~\1238(487)  | ~\1237(462) ,
  \1480(187)  = ~\1474(105) ,
  \285(628)  = ~\279(609) ,
  \1813(629)  = ~\1809(610) ,
  \1733(488)  = ~\1729(468) ,
  \1717(208)  = ~\1713(118) ,
  \1854(158)  = \168(79) ,
  \407(474)  = ~\296(454) ,
  \32(828)  = ~\1593(797)  | ~\1586(70) ,
  \1584(143)  = ~\1578(72) ,
  \1312(166)  = \160(83) ,
  \1870(141)  = \184(71) ,
  \295(437)  = ~\1049(413)  | ~\1040(249) ,
  \1024(640)  = ~\1693(602)  | ~\1686(626) ,
  \1044(320)  = ~\1709(243)  | ~\1702(246) ,
  \1562(76)  = \122(7) ,
  \1889(464)  = ~\390(446) ,
  \1277(401)  = ~\1273(372) ,
  \1157(355)  = ~\1788(294)  | ~\1785(164) ,
  \260(421)  = ~\988(333)  | ~\985(384) ,
  \520(706)  = ~\1456(192)  | ~\1453(694) ,
  \1709(243)  = ~\1705(154) ,
  \1512(178)  = ~\1506(90) ,
  \327(137)  = \188(69) ,
  \1201(263)  = ~\1197(176) ,
  \1568(152)  = ~\1562(76) ,
  \1409(622)  = ~\1405(604) ,
  \857(784)  = ~\804(757)  | (~\800(756)  | (~\796(755)  | (~\792(754)  | (~\788(753)  | (~\784(752)  | (~\780(751)  | ~\776(750) )))))),
  \60(901)  = \[19] ,
  \1165(423)  = ~\1163(397)  | ~\1154(193) ,
  \1766(515)  = \343(492) ,
  \1910(631)  = \853(97)  & \285(628) ,
  \1192(399)  = ~\1184(370) ,
  \1537(788)  = ~\1533(761) ,
  \499(713)  = ~\1417(699)  | ~\1410(279) ,
  \424(644)  = ~\1385(425)  | ~\1378(630) ,
  \1605(778)  = \969(266)  & (\731(676)  & (\710(728)  & (\639B(735)  & \573(738) ))),
  \1474(105)  = \541(50) ,
  \392(526)  = ~\1299(506)  | ~\1290(115) ,
  \1110(405)  = ~\1108(307)  | ~\1105(373) ,
  \614(271)  = ~\487(197) ,
  \233(57)  = ~\900(29)  | ~\227(21) ,
  \836(773)  = ~\969(266)  | (~\756(677)  | (~\710(728)  | (~\639B(735)  | ~\588B(740) ))),
  \1138(544)  = ~\1773(501)  | ~\1766(515) ,
  \324(546)  = ~\1098(270)  | ~\1095(539) ,
  \1804(466)  = ~\1798(448) ,
  \1597(777)  = \969(266)  & (\746(678)  & (\696(726)  & (\639B(735)  & \573(738) ))),
  \1789(252)  = ~\1785(164) ,
  \1013(520)  = ~\1684(497)  | ~\1681(503) ,
  \1043(354)  = ~\1708(323)  | ~\1705(154) ,
  \1578(72)  = \128(9) ,
  \1143(594)  = ~\1139(577) ,
  \306(433)  = ~\1077(394)  | ~\1068(231) ,
  \998(334)  = ~\990(262) ,
  \528(723)  = ~\522(719) ,
  \1909(511)  = ~\1905(486) ,
  \907(48)  = ~\898(28) ,
  \1322(361)  = ~\406(335) ,
  \425(674)  = ~\424(644)  | ~\423(663) ,
  \956(181)  = ~\893(111)  | (~\943(35)  | (~\919(44)  | ~\907(48) )),
  \188(69)  = ~\131(10) ,
  \346(587)  = ~\1142(531)  | ~\1139(577) ,
  \296(454)  = ~\295(437)  | ~\294(415) ,
  \1397(564)  = \393(548) ,
  \1081(494)  = ~\1732(313)  | ~\1729(468) ,
  \18(860)  = \[8] ,
  \881(747)  = ~\979(179)  | (~\731(676)  | (~\688(727)  | (~\622(733)  | ~\573(738) ))),
  \1602(66)  = \137(12) ,
  \305(409)  = ~\1076(310)  | ~\1073(366) ,
  \1293(476)  = ~\1868(447)  | ~\1865(439) ,
  \1183(218)  = ~\1179(127) ,
  \1585(796)  = ~\1581(775) ,
  \1327(528)  = ~\1326(523)  | ~\1325(481) ,
  \1830(116)  = \938(36)  & (\241(54)  & \214(17) ),
  \1702(246)  = \291(157) ,
  \1788(294)  = ~\1782(216) ,
  \65(895)  = ~\431(877)  | ~\430(885) ,
  \39(853)  = \[14] ,
  \688(727)  = \669(715)  & \666(685) ,
  \325(562)  = ~\1099(554)  | ~\1090(196) ,
  \1865(439)  = ~\1289(419)  | ~\1288(386) ,
  \1761(477)  = \262(458) ,
  \517(52)  = ~\469(24) ,
  \75(866)  = \[16] ,
  \500(720)  = ~\499(713)  | ~\498(707) ,
  \14(834)  = ~\1545(789)  | ~\1538(82) ,
  \639A(734)  = \639(724) ,
  \1408(870)  = ~\1402(845) ,
  \588(729)  = \500(720)  & \566(277) ,
  \1254(376)  = ~\1252(229)  | ~\1249(338) ,
  \1449(701)  = ~\1445(693) ,
  \1661(255)  = ~\1657(168) ,
  \288(160)  = \165(81) ,
  \1226(327)  = ~\1821(240)  | ~\1814(161) ,
  \621(732)  = \618(722)  & \614(271) ,
  \1565(765)  = \958(265)  & (\770(679)  & (\675(725)  & (\622(733)  & \588B(740) ))),
  \364(565)  = ~\1192(399)  | ~\1189(550) ,
  \1381(392)  = ~\374(364) ,
  \1348(521)  = ~\1340(498) ,
  \1058(230)  = \299(140) ,
  \537(709)  = ~\536(703)  | ~\535(697) ,
  \359(424)  = ~\1175(398)  | ~\1166(194) ,
  \1303(292)  = ~\1876(232)  | ~\1873(124) ,
  \1618(62)  = \143(14) ,
  \314(471)  = ~\307(452) ,
  \35(827)  = ~\1601(798)  | ~\1594(68) ,
  \398(438)  = ~\397(416)  | ~\396(383) ,
  \1536(167)  = ~\1530(84) ,
  \1790(217)  = \355(126) ,
  \1147(658)  = ~\1780(645)  | ~\1777(461) ,
  \1315(312)  = ~\1884(244)  | ~\1881(142) ,
  \50(91)  = ~\947(34)  | ~\930(41) ,
  \1369(621)  = ~\1365(603) ,
  \746(678)  = \725(665)  & \722(653) ,
  \1506(90)  = \101(0) ,
  \1233(420)  = ~\1231(379)  | ~\1222(173) ,
  \1019(572)  = ~\1015(556) ,
  \1812(873)  = ~\1806(848) ,
  \51(899)  = \[17] ,
  \1876(232)  = ~\1870(141) ,
  \877(745)  = ~\979(179)  | (~\756(677)  | (~\675(725)  | (~\622(733)  | ~\573(738) ))),
  \1299(506)  = ~\1295(483) ,
  \1077(394)  = ~\1073(366) ,
  \206(59)  = ~\146(15) ,
  \1008(434)  = ~\1000(410) ,
  \503(731)  = ~\497(721) ,
  \149(89)  = ~\101(0) ,
  \1857(151)  = \175(75) ,
  \1109(402)  = ~\1105(373) ,
  \1653(890)  = ~\1649(882) ,
  \984(329)  = ~\1661(255)  | ~\1654(258) ,
  \1305(343)  = ~\1304(311)  | ~\1303(292) ,
  \1637(839)  = ~\1916(650)  | ~\1913(822) ,
  \298(328)  = ~\1057(239)  | ~\1050(163) ,
  \307(452)  = ~\306(433)  | ~\305(409) ,
  \1260(298)  = ~\1845(237)  | ~\1838(219) ,
  \1793(165)  = \160(83) ,
  \954(101)  = ~\922(43)  | ~\248(55) ,
  \1617(800)  = ~\1613(779) ,
  \1684(497)  = ~\1678(473) ,
  \1893(482)  = ~\1889(464) ,
  \1384(649)  = ~\1378(630) ,
  \1020(844)  = \462(820)  & (\911(46)  & \457(205) ),
  \1533(761)  = \958(265)  & (\731(676)  & (\688(727)  & (\639A(734)  & \588A(739) ))),
  \1694(245)  = \291(157) ,
  \309(432)  = ~\1067(393)  | ~\1058(230) ,
  \1442(109)  = \517(52) ,
  \1708(323)  = ~\1702(246) ,
  \352(112)  = \938(36)  & \227(21) ,
  \1261(371)  = ~\1260(298)  | ~\1259(348) ,
  \1841(146)  = \179(73) ,
  \1456(192)  = ~\1450(110) ,
  \1290(115)  = \938(36)  & (\245(56)  & \217(18) ),
  \722(653)  = \561(635) ,
  \63(902)  = \[20] ,
  \1437(616)  = \453(599) ,
  \179(73)  = ~\125(8) ,
  \1522(86)  = \107(2) ,
  \560(617)  = ~\1497(597)  | ~\1490(103) ,
  \1828(450)  = ~\1822(431) ,
  \1094(518)  = ~\1741(489)  | ~\1734(235) ,
  \995(385)  = ~\994(330)  | ~\993(358) ,
  \1072(286)  = ~\1725(209)  | ~\1718(213) ,
  \308(408)  = ~\1066(309)  | ~\1063(365) ,
  \1148(639)  = ~\1781(480)  | ~\1774(624) ,
  \1402(845)  = \462(820)  & (\911(46)  & \459(200) ),
  \545(638)  = ~\1489(614)  | ~\1482(106) ,
  \10(815)  = ~\1536(167)  | ~\1533(761) ,
  \1298(201)  = ~\1290(115) ,
  \1268(211)  = \382(120) ,
  \1289(419)  = ~\1287(380)  | ~\1278(170) ,
  \184(71)  = ~\128(9) ,
  \1370(646)  = ~\348(625) ,
  \1553(790)  = ~\1549(763) ,
  \725(665)  = ~\549(655) ,
  \1657(168)  = \156(85) ,
  \1112(228)  = \327(137) ,
  \31(808)  = ~\1592(139)  | ~\1589(776) ,
  \523(705)  = ~\1448(191)  | ~\1445(693) ,
  \1576(148)  = ~\1570(74) ,
  \804(757)  = ~\958(265)  | (~\770(679)  | (~\675(725)  | (~\622(733)  | ~\588B(740) ))),
  \1453(694)  = \437(688) ,
  \302(122)  = \202(61) ,
  \1163(397)  = ~\1159(368) ,
  \1176(145)  = \179(73) ,
  \374(364)  = ~\373(283)  | ~\372(360) ,
  \1724(290)  = ~\1718(213) ,
  \1308(226)  = ~\1300(135) ,
  \1179(127)  = \198(63) ,
  \1538(82)  = \113(4) ,
  \17(833)  = ~\1553(790)  | ~\1546(80) ,
  \1331(549)  = ~\1327(528) ,
  \1066(309)  = ~\1058(230) ,
  \1498(104)  = \553(49) ,
  \1222(173)  = \153(87) ,
  \350(875)  = ~\1153(681)  | ~\1144(849) ,
  \378(557)  = ~\1243(527)  | ~\1234(440) ,
  \1678(473)  = \274(453) ,
  \1740(314)  = ~\1734(235) ,
  \334(430)  = ~\1121(403)  | ~\1112(228) ,
  \919(44)  = \902(30) ,
  \245(56)  = \234(22) ,
  \1878(155)  = \171(77) ,
  \38(826)  = ~\1609(799)  | ~\1602(66) ,
  \1015(556)  = ~\1014(541)  | ~\1013(520) ,
  \1726(234)  = \321(144) ,
  \1570(74)  = \125(8) ,
  \1805(516)  = ~\1801(493) ,
  \1217(897)  = ~\1216(879)  | ~\1215(887) ,
  \1441(634)  = ~\1437(616) ,
  \333(406)  = ~\1120(308)  | ~\1117(374) ,
  \1211(264)  = ~\1207(177) ,
  \1852(301)  = ~\1846(220) ,
  \279(609)  = ~\278(589)  | ~\277(570) ;
endmodule

