// IWLS benchmark module "CM163" printed on Wed May 29 16:31:28 2002
module cm163a(a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u);
input
  a,
  b,
  c,
  d,
  e,
  f,
  g,
  h,
  i,
  j,
  k,
  l,
  m,
  n,
  o,
  p;
output
  q,
  r,
  s,
  t,
  u;
wire
  o0,
  p0,
  q0,
  r0,
  g0,
  h0,
  \[0] ,
  i0,
  \[1] ,
  j0,
  \[2] ,
  \[3] ,
  l0,
  \[4] ,
  m0,
  n0;
assign
  o0 = (~n & ~r0) | (n & r0),
  p0 = ~p | (~i | (~k | ~o)),
  q0 = ~l & (~j & ~l0),
  r0 = ~l & (~j & (~l0 & ~m)),
  g0 = f & ~e,
  h0 = f & e,
  \[0]  = (~h0 & ~g0) | ((~h0 & ~a) | ((~i0 & ~g0) | (~i0 & ~a))),
  i0 = (~j & l0) | (j & ~l0),
  \[1]  = (~h0 & ~g0) | ((~h0 & ~b) | ((~j0 & ~g0) | (~j0 & ~b))),
  q = \[0] ,
  r = \[1] ,
  s = \[2] ,
  j0 = (~l & ~m0) | (l & m0),
  t = \[3] ,
  \[2]  = (~h0 & ~g0) | ((~h0 & ~g) | ((~n0 & ~g0) | (~n0 & ~g))),
  u = \[4] ,
  \[3]  = (~h0 & ~g0) | ((~h0 & ~h) | ((~o0 & ~g0) | (~o0 & ~h))),
  l0 = ~d | ~c,
  \[4]  = d & ~p0,
  m0 = ~l0 & ~j,
  n0 = (~m & ~q0) | (m & q0);
endmodule

