module in6 (
    x0,
    x1,
    x2,
    x3,
    x4,
    x5,
    x6,
    x7,
    x8,
    x9,
    x10,
    x11,
    x12,
    x13,
    x14,
    x15,
    x16,
    x17,
    x18,
    x19,
    x20,
    x21,
    x22,
    x23,
    x24,
    x25,
    x26,
    x27,
    x28,
    x29,
    x30,
    x31,
    x32,
    y0,
    y1,
    y2,
    y3,
    y4,
    y5,
    y6,
    y7,
    y8,
    y9,
    y10,
    y11,
    y12,
    y13,
    y14,
    y15,
    y16,
    y17,
    y18,
    y19,
    y20,
    y21,
    y22
);
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 ;
  wire n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 ;
  assign n36  = ~x15 & x31;
  assign n37  = ~x16 & n36;
  assign n34  = x28 & ~x31;
  assign n35  = x30 & n34;
  assign n38  = (x1 & n35) | (x1 & n37) | (n35 & n37);
  assign n39  = x22 & ~n38;
  assign n40  = (x22 & n37) | (x22 & ~n39) | (n37 & ~n39);
  assign n41  = ~x0 & n40;
  assign n46  = (~x0 & x4) | (~x0 & x32) | (x4 & x32);
  assign n42  = x28 & ~x32;
  assign n43  = x29 & n42;
  assign n44  = x24 & n43;
  assign n45  = x1 & n44;
  assign n47  = ~x0 & n45;
  assign n48  = (~x4 & n46) | (~x4 & n47) | (n46 & n47);
  assign n49  = x3 & ~x28;
  assign n50  = (x0 & ~x30) | (x0 & n49) | (~x30 & n49);
  assign n51  = ~x0 & n50;
  assign n52  = ~x28 & x29;
  assign n53  = ~x30 & n52;
  assign n54  = x0 | n53;
  assign n55  = (x0 & x3) | (x0 & n54) | (x3 & n54);
  assign n56  = (x11 & ~x12) | (x11 & x29) | (~x12 & x29);
  assign n57  = ~x10 & x29;
  assign n58  = (~x11 & n56) | (~x11 & n57) | (n56 & n57);
  assign n59  = x19 & x21;
  assign n60  = (x20 & ~n58) | (x20 & n59) | (~n58 & n59);
  assign n61  = n58 & n60;
  assign n79  = ~x9 & n61;
  assign n62  = ~x10 & x11;
  assign n63  = (x9 & ~x12) | (x9 & n62) | (~x12 & n62);
  assign n64  = ~x9 & n63;
  assign n65  = x11 | x12;
  assign n70  = (~x12 & x20) | (~x12 & x29) | (x20 & x29);
  assign n71  = (x12 & x21) | (x12 & x29) | (x21 & x29);
  assign n72  = n70 & n71;
  assign n73  = x19 & n72;
  assign n74  = x11 & ~n73;
  assign n75  = n65 & ~n74;
  assign n76  = (~x9 & x10) | (~x9 & n75) | (x10 & n75);
  assign n66  = x21 & ~x29;
  assign n67  = (x12 & ~x21) | (x12 & n66) | (~x21 & n66);
  assign n68  = (x11 & x12) | (x11 & n67) | (x12 & n67);
  assign n69  = (n65 & n67) | (n65 & ~n68) | (n67 & ~n68);
  assign n77  = (x9 & x10) | (x9 & ~n69) | (x10 & ~n69);
  assign n78  = n76 & n77;
  assign n80  = n64 | n78;
  assign n81  = (n61 & ~n79) | (n61 & n80) | (~n79 & n80);
  assign n82  = ~x0 & x30;
  assign n83  = (x28 & n81) | (x28 & ~n82) | (n81 & ~n82);
  assign n84  = n81 & ~n83;
  assign n85  = x10 & ~x11;
  assign n86  = (x9 & ~x12) | (x9 & n85) | (~x12 & n85);
  assign n87  = ~x9 & n86;
  assign n88  = x15 & ~x28;
  assign n89  = (x14 & x17) | (x14 & n88) | (x17 & n88);
  assign n90  = ~x14 & n89;
  assign n101 = (x30 & ~n87) | (x30 & n90) | (~n87 & n90);
  assign n91  = (~x6 & x15) | (~x6 & x17) | (x15 & x17);
  assign n92  = ~x15 & n91;
  assign n93  = (x7 & ~x17) | (x7 & n92) | (~x17 & n92);
  assign n94  = (n91 & n92) | (n91 & n93) | (n92 & n93);
  assign n95  = (~x14 & x15) | (~x14 & n94) | (x15 & n94);
  assign n96  = x17 & ~n95;
  assign n97  = (x17 & n94) | (x17 & ~n96) | (n94 & ~n96);
  assign n98  = x1 & x28;
  assign n99  = (x23 & ~n97) | (x23 & n98) | (~n97 & n98);
  assign n100 = n97 & n99;
  assign n102 = x30 & n100;
  assign n103 = (n87 & n101) | (n87 & n102) | (n101 & n102);
  assign n104 = ~x16 & n103;
  assign n105 = (x0 & ~x18) | (x0 & n104) | (~x18 & n104);
  assign n106 = ~x0 & n105;
  assign n107 = x11 | x28;
  assign n108 = x12 | n107;
  assign n109 = ~x9 & x10;
  assign n110 = ~n108 & n109;
  assign n111 = (x1 & x23) | (x1 & n110) | (x23 & n110);
  assign n112 = x28 & ~n111;
  assign n113 = (x28 & n110) | (x28 & ~n112) | (n110 & ~n112);
  assign n114 = x16 & x18;
  assign n115 = x17 & ~x18;
  assign n116 = x6 | x16;
  assign n117 = x17 & n116;
  assign n118 = (n114 & n115) | (n114 & ~n117) | (n115 & ~n117);
  assign n132 = (x30 & ~n113) | (x30 & n118) | (~n113 & n118);
  assign n119 = ~x17 & x18;
  assign n120 = x18 & ~n119;
  assign n121 = ~x8 & n120;
  assign n122 = (x17 & n119) | (x17 & ~n121) | (n119 & ~n121);
  assign n123 = (~x6 & n119) | (~x6 & n122) | (n119 & n122);
  assign n124 = ~x16 & x23;
  assign n125 = (~x28 & n123) | (~x28 & n124) | (n123 & n124);
  assign n126 = ~n123 & n125;
  assign n127 = x12 & n126;
  assign n128 = (x10 & x11) | (x10 & n127) | (x11 & n127);
  assign n129 = ~x10 & n128;
  assign n130 = ~x9 & n129;
  assign n131 = x1 & n130;
  assign n133 = x30 & n131;
  assign n134 = (n113 & n132) | (n113 & n133) | (n132 & n133);
  assign n135 = ~x0 & n134;
  assign n136 = ~x15 & n135;
  assign n137 = x11 & x12;
  assign n138 = (x9 & x10) | (x9 & ~x28) | (x10 & ~x28);
  assign n139 = n137 & n138;
  assign n140 = (x28 & n137) | (x28 & ~n139) | (n137 & ~n139);
  assign n141 = ~x18 & x22;
  assign n142 = (x15 & ~n140) | (x15 & n141) | (~n140 & n141);
  assign n143 = n140 & n142;
  assign n150 = (x1 & x30) | (x1 & ~n143) | (x30 & ~n143);
  assign n144 = (x1 & x22) | (x1 & n110) | (x22 & n110);
  assign n145 = x28 & ~n144;
  assign n146 = (x28 & n110) | (x28 & ~n145) | (n110 & ~n145);
  assign n147 = ~x0 & x18;
  assign n148 = (x15 & n146) | (x15 & ~n147) | (n146 & ~n147);
  assign n149 = n146 & ~n148;
  assign n151 = x30 & n149;
  assign n152 = (n143 & n150) | (n143 & n151) | (n150 & n151);
  assign n153 = (x0 & x16) | (x0 & ~x17) | (x16 & ~x17);
  assign n154 = n152 & ~n153;
  assign n155 = (x0 & n152) | (x0 & ~n154) | (n152 & ~n154);
  assign n156 = x16 & ~x17;
  assign n157 = x22 & x28;
  assign n158 = (~x16 & n156) | (~x16 & n157) | (n156 & n157);
  assign n181 = (x1 & x30) | (x1 & ~n158) | (x30 & ~n158);
  assign n165 = x16 & x22;
  assign n166 = (x17 & n137) | (x17 & n165) | (n137 & n165);
  assign n167 = ~x17 & n166;
  assign n168 = x1 & ~x10;
  assign n169 = (x6 & x8) | (x6 & n168) | (x8 & n168);
  assign n170 = ~x6 & n169;
  assign n175 = (x0 & n167) | (x0 & ~n170) | (n167 & ~n170);
  assign n171 = ~x12 & n85;
  assign n172 = ~x16 & x17;
  assign n173 = (x14 & n171) | (x14 & n172) | (n171 & n172);
  assign n174 = ~x14 & n173;
  assign n176 = ~x0 & n174;
  assign n177 = (n167 & ~n175) | (n167 & n176) | (~n175 & n176);
  assign n159 = x12 | x17;
  assign n160 = (~x11 & x16) | (~x11 & n159) | (x16 & n159);
  assign n161 = x11 | n160;
  assign n162 = x10 & ~n161;
  assign n163 = (x6 & x7) | (x6 & n162) | (x7 & n162);
  assign n164 = ~x6 & n163;
  assign n178 = n164 & ~n177;
  assign n179 = x9 | x28;
  assign n180 = (n177 & n178) | (n177 & ~n179) | (n178 & ~n179);
  assign n182 = x30 & n180;
  assign n183 = (n158 & n181) | (n158 & n182) | (n181 & n182);
  assign n184 = (x0 & x15) | (x0 & ~x18) | (x15 & ~x18);
  assign n185 = n183 & ~n184;
  assign n186 = (x0 & n183) | (x0 & ~n185) | (n183 & ~n185);
  assign n187 = x17 & n88;
  assign n188 = ~x12 & n187;
  assign n189 = ~x14 & n188;
  assign n190 = (x0 & ~x11) | (x0 & n109) | (~x11 & n109);
  assign n191 = ~x0 & n190;
  assign n201 = (x30 & ~n189) | (x30 & n191) | (~n189 & n191);
  assign n192 = (x14 & x15) | (x14 & ~x17) | (x15 & ~x17);
  assign n193 = n91 & ~n192;
  assign n194 = ~x6 & x7;
  assign n195 = ~x17 & n194;
  assign n196 = x15 & n195;
  assign n197 = x0 & ~n196;
  assign n198 = (n193 & n196) | (n193 & ~n197) | (n196 & ~n197);
  assign n199 = (x22 & n98) | (x22 & ~n198) | (n98 & ~n198);
  assign n200 = n198 & n199;
  assign n202 = x30 & n200;
  assign n203 = (n189 & n201) | (n189 & n202) | (n201 & n202);
  assign n204 = x0 & x7;
  assign n205 = (x16 & x18) | (x16 & ~n204) | (x18 & ~n204);
  assign n206 = n203 & n205;
  assign n207 = (n203 & n204) | (n203 & ~n206) | (n204 & ~n206);
  assign n220 = x6 & ~x16;
  assign n221 = (x6 & x8) | (x6 & x16) | (x8 & x16);
  assign n222 = ~x15 & x16;
  assign n223 = (n220 & n221) | (n220 & ~n222) | (n221 & ~n222);
  assign n226 = (x0 & x28) | (x0 & n223) | (x28 & n223);
  assign n224 = x7 & ~x15;
  assign n225 = ~x16 & n224;
  assign n227 = ~x28 & n225;
  assign n228 = (n223 & ~n226) | (n223 & n227) | (~n226 & n227);
  assign n229 = x12 & n228;
  assign n230 = (x10 & x11) | (x10 & n229) | (x11 & n229);
  assign n231 = ~x10 & n230;
  assign n235 = (x9 & ~x18) | (x9 & n231) | (~x18 & n231);
  assign n232 = x15 & x28;
  assign n233 = (x16 & n194) | (x16 & n232) | (n194 & n232);
  assign n234 = ~x16 & n233;
  assign n236 = ~x18 & n234;
  assign n237 = (~x9 & n235) | (~x9 & n236) | (n235 & n236);
  assign n208 = x0 | x15;
  assign n217 = x16 & x28;
  assign n218 = (x18 & n208) | (x18 & n217) | (n208 & n217);
  assign n219 = ~n208 & n218;
  assign n238 = n219 & ~n237;
  assign n239 = x1 & x22;
  assign n240 = (n237 & n238) | (n237 & n239) | (n238 & n239);
  assign n209 = x15 & ~x18;
  assign n210 = (x16 & n194) | (x16 & n209) | (n194 & n209);
  assign n211 = ~x16 & n210;
  assign n212 = (x16 & ~n208) | (x16 & n211) | (~n208 & n211);
  assign n213 = x18 & ~n212;
  assign n214 = (x18 & n211) | (x18 & ~n213) | (n211 & ~n213);
  assign n215 = (x12 & n107) | (x12 & n214) | (n107 & n214);
  assign n216 = n214 & ~n215;
  assign n241 = (~x9 & n216) | (~x9 & n240) | (n216 & n240);
  assign n242 = x10 & ~n241;
  assign n243 = (x10 & n240) | (x10 & ~n242) | (n240 & ~n242);
  assign n244 = (~x17 & n204) | (~x17 & n243) | (n204 & n243);
  assign n245 = x30 & ~n244;
  assign n246 = (x30 & n204) | (x30 & ~n245) | (n204 & ~n245);
  assign n247 = (x16 & x17) | (x16 & x23) | (x17 & x23);
  assign n248 = (x16 & x17) | (x16 & ~x28) | (x17 & ~x28);
  assign n249 = n247 & ~n248;
  assign n250 = ~x28 & n156;
  assign n257 = (x9 & n171) | (x9 & ~n250) | (n171 & ~n250);
  assign n251 = x12 & x23;
  assign n252 = (x16 & x17) | (x16 & n251) | (x17 & n251);
  assign n253 = ~x16 & n252;
  assign n254 = x1 & x11;
  assign n255 = (x10 & n253) | (x10 & n254) | (n253 & n254);
  assign n256 = ~x10 & n255;
  assign n258 = ~x9 & n256;
  assign n259 = (n171 & ~n257) | (n171 & n258) | (~n257 & n258);
  assign n260 = x1 | n259;
  assign n261 = (n249 & n259) | (n249 & n260) | (n259 & n260);
  assign n262 = ~x15 & x30;
  assign n263 = (x18 & ~n261) | (x18 & n262) | (~n261 & n262);
  assign n264 = n261 & n263;
  assign n265 = ~x0 & n264;
  assign n266 = (x0 & ~n204) | (x0 & n265) | (~n204 & n265);
  assign n267 = x23 & x28;
  assign n268 = (~x15 & n209) | (~x15 & n267) | (n209 & n267);
  assign n285 = (x1 & x30) | (x1 & ~n268) | (x30 & ~n268);
  assign n275 = x1 & ~x8;
  assign n276 = ~x10 & n275;
  assign n277 = x23 & n276;
  assign n278 = (x18 & ~n137) | (x18 & n277) | (~n137 & n277);
  assign n279 = n137 & n278;
  assign n272 = x10 & ~x12;
  assign n273 = (x11 & ~x18) | (x11 & n272) | (~x18 & n272);
  assign n274 = ~x11 & n273;
  assign n280 = n274 & ~n279;
  assign n281 = x6 | x15;
  assign n282 = (n279 & n280) | (n279 & ~n281) | (n280 & ~n281);
  assign n269 = ~x18 & n171;
  assign n270 = (x14 & x15) | (x14 & n269) | (x15 & n269);
  assign n271 = ~x14 & n270;
  assign n283 = n271 & ~n282;
  assign n284 = (~n179 & n282) | (~n179 & n283) | (n282 & n283);
  assign n286 = x30 & n284;
  assign n287 = (n268 & n285) | (n268 & n286) | (n285 & n286);
  assign n288 = n172 & n287;
  assign n289 = ~x0 & n288;
  assign n290 = (x0 & ~n204) | (x0 & n289) | (~n204 & n289);
  assign n291 = (x0 & x24) | (x0 & x29) | (x24 & x29);
  assign n292 = x25 & x29;
  assign n293 = (~x0 & n291) | (~x0 & n292) | (n291 & n292);
  assign n294 = (x0 & x1) | (x0 & n293) | (x1 & n293);
  assign n295 = x28 & ~n294;
  assign n296 = (x0 & x28) | (x0 & ~n295) | (x28 & ~n295);
  assign n297 = x1 & ~x22;
  assign n298 = (x0 & x13) | (x0 & n297) | (x13 & n297);
  assign n299 = ~x0 & n298;
  assign n300 = x24 & x29;
  assign n301 = (x28 & ~n299) | (x28 & n300) | (~n299 & n300);
  assign n302 = n299 & n301;
  assign n303 = (x0 & x24) | (x0 & n98) | (x24 & n98);
  assign n304 = ~x0 & n303;
  assign n305 = x29 & n304;
  assign n306 = (x5 & x22) | (x5 & x28) | (x22 & x28);
  assign n307 = x30 & ~n306;
  assign n308 = (x5 & x30) | (x5 & ~n307) | (x30 & ~n307);
  assign n309 = ~x0 & n308;
  assign n310 = ~x12 & x30;
  assign n311 = (x11 & ~x28) | (x11 & n310) | (~x28 & n310);
  assign n312 = ~x11 & n311;
  assign n313 = (x0 & n109) | (x0 & n312) | (n109 & n312);
  assign n314 = ~x0 & n313;
  assign n315 = (x3 & x27) | (x3 & ~n314) | (x27 & ~n314);
  assign n316 = x26 | n314;
  assign n317 = (x27 & ~n315) | (x27 & n316) | (~n315 & n316);
  assign n318 = x0 | n317;
  assign n319 = (~x3 & x27) | (~x3 & n314) | (x27 & n314);
  assign n320 = (x3 & x26) | (x3 & n314) | (x26 & n314);
  assign n321 = n319 | n320;
  assign n322 = (~x27 & n319) | (~x27 & n321) | (n319 & n321);
  assign n323 = x0 | n322;
  assign n324 = (x10 & ~x11) | (x10 & n61) | (~x11 & n61);
  assign n325 = x12 & ~n324;
  assign n326 = (x12 & n61) | (x12 & ~n325) | (n61 & ~n325);
  assign n327 = (~x12 & x19) | (~x12 & x20) | (x19 & x20);
  assign n328 = (x12 & x19) | (x12 & x21) | (x19 & x21);
  assign n329 = n327 & n328;
  assign n330 = x9 & ~n329;
  assign n331 = x12 & x21;
  assign n332 = x9 | n331;
  assign n333 = ~n330 & n332;
  assign n334 = x29 & n333;
  assign n335 = x10 & ~n334;
  assign n336 = x9 | x12;
  assign n337 = ~x10 & n336;
  assign n338 = n335 | n337;
  assign n339 = x11 & ~n338;
  assign n340 = x9 | n339;
  assign n341 = (n326 & n339) | (n326 & n340) | (n339 & n340);
  assign n342 = (x28 & ~n82) | (x28 & n341) | (~n82 & n341);
  assign n343 = n341 & ~n342;
  assign n344 = (x2 & x29) | (x2 & ~x30) | (x29 & ~x30);
  assign n345 = (x3 & x29) | (x3 & x30) | (x29 & x30);
  assign n346 = n344 & ~n345;
  assign n347 = x21 & x29;
  assign n348 = (x11 & ~n65) | (x11 & n347) | (~n65 & n347);
  assign n349 = x20 & n348;
  assign n350 = (x10 & x19) | (x10 & n349) | (x19 & n349);
  assign n351 = ~x10 & n350;
  assign n354 = (~x10 & x11) | (~x10 & x12) | (x11 & x12);
  assign n355 = x12 & ~n354;
  assign n352 = x19 & x29;
  assign n353 = x21 & n352;
  assign n356 = (x11 & n353) | (x11 & n355) | (n353 & n355);
  assign n357 = (~n354 & n355) | (~n354 & n356) | (n355 & n356);
  assign n358 = x12 & x29;
  assign n359 = x21 & n358;
  assign n360 = x11 & n359;
  assign n361 = (x9 & x10) | (x9 & n360) | (x10 & n360);
  assign n362 = ~x9 & n361;
  assign n363 = (~n351 & n357) | (~n351 & n362) | (n357 & n362);
  assign n364 = x9 | n362;
  assign n365 = (n351 & n363) | (n351 & n364) | (n363 & n364);
  assign n366 = x30 & ~n365;
  assign n367 = x3 & ~x29;
  assign n368 = x30 | n367;
  assign n369 = ~n366 & n368;
  assign n370 = (x0 & ~n346) | (x0 & n369) | (~n346 & n369);
  assign n371 = ~x0 & x28;
  assign n372 = (n346 & n370) | (n346 & ~n371) | (n370 & ~n371);
  assign n391 = (x3 & ~x28) | (x3 & x30) | (~x28 & x30);
  assign n380 = x20 & x29;
  assign n381 = x21 & n380;
  assign n382 = x9 & x19;
  assign n383 = (x12 & ~n381) | (x12 & n382) | (~n381 & n382);
  assign n384 = n381 & n383;
  assign n385 = (x9 & x12) | (x9 & ~n384) | (x12 & ~n384);
  assign n386 = x11 & n385;
  assign n387 = (x11 & n384) | (x11 & ~n386) | (n384 & ~n386);
  assign n388 = ~x10 & n387;
  assign n373 = ~x11 & x12;
  assign n374 = x12 & ~n373;
  assign n375 = x10 & n374;
  assign n376 = (x21 & ~n373) | (x21 & n374) | (~n373 & n374);
  assign n377 = (~x11 & n375) | (~x11 & n376) | (n375 & n376);
  assign n378 = (x20 & n352) | (x20 & ~n377) | (n352 & ~n377);
  assign n379 = n377 & n378;
  assign n389 = n379 | n388;
  assign n390 = (x9 & n388) | (x9 & n389) | (n388 & n389);
  assign n392 = (x28 & x30) | (x28 & ~n390) | (x30 & ~n390);
  assign n393 = n391 & ~n392;
  assign n394 = ~x0 & n393;
  assign n395 = x9 & x11;
  assign n396 = (x0 & x10) | (x0 & n395) | (x10 & n395);
  assign n397 = ~x0 & n396;
  assign n398 = x12 & x20;
  assign n399 = (x19 & ~n397) | (x19 & n398) | (~n397 & n398);
  assign n400 = n397 & n399;
  assign n401 = x30 & n400;
  assign n402 = (x28 & x29) | (x28 & n401) | (x29 & n401);
  assign n403 = ~x28 & n402;
  assign y0   = n41;
  assign y1   = n48;
  assign y2   = n51;
  assign y3   = n55;
  assign y4   = n84;
  assign y5   = n106;
  assign y6   = n136;
  assign y7   = n155;
  assign y8   = n186;
  assign y9   = n207;
  assign y10  = n246;
  assign y11  = n266;
  assign y12  = n290;
  assign y13  = n296;
  assign y14  = n302;
  assign y15  = n305;
  assign y16  = n309;
  assign y17  = n318;
  assign y18  = n323;
  assign y19  = n343;
  assign y20  = n372;
  assign y21  = n394;
  assign y22  = n403;
endmodule
