// IWLS benchmark module "x4" printed on Wed May 29 17:30:39 2002
module x4(a, b, g, h, i, k, l, m, n, o, p, q, r, s, t, u, v, w, \xx , y, z, a0, b0, c0, d0, e0, f0, g0, h0, i0, k0, l0, m0, n0, o0, p0, q0, r0, s0, t0, u0, v0, w0, x0, y0, z0, a1, b1, c1, d1, e1, f1, g1, h1, i1, j1, k1, l1, m1, n1, o1, p1, q1, r1, s1, t1, u1, v1, w1, x1, y1, z1, a2, b2, c2, d2, e2, f2, g2, h2, i2, j2, k2, l2, m2, n2, o2, p2, q2, r2, s2, t2, u2, v2, w2, x2, y2, z2, a3, b3, c3, d3, e3, f3, g3, h3, i3, j3, k3, l3, m3, n3, o3, p3, q3, r3, s3, t3, u3, v3, w3, x3, y3, z3, a4, b4, c4, d4, e4, f4, g4, h4, i4, j4, k4, l4, m4, n4, o4, p4, q4, r4, s4, t4, u4, v4, w4, x4, y4, z4, a5, b5, c5, d5, e5, f5, g5, h5, i5, j5, k5, l5, m5, n5, o5);
input
  z0,
  z1,
  a,
  b,
  g,
  h,
  i,
  k,
  l,
  m,
  n,
  o,
  p,
  q,
  r,
  s,
  t,
  u,
  v,
  w,
  \xx ,
  y,
  z,
  a0,
  a1,
  a2,
  b0,
  b1,
  b2,
  c0,
  c1,
  c2,
  d0,
  d1,
  d2,
  e0,
  e1,
  e2,
  f0,
  f1,
  f2,
  g0,
  g1,
  g2,
  h0,
  h1,
  h2,
  i0,
  i1,
  i2,
  j1,
  j2,
  k0,
  k1,
  k2,
  l0,
  l1,
  l2,
  m0,
  m1,
  m2,
  n0,
  n1,
  n2,
  o0,
  o1,
  o2,
  p0,
  p1,
  p2,
  q0,
  q1,
  q2,
  r0,
  r1,
  r2,
  s0,
  s1,
  s2,
  t0,
  t1,
  t2,
  u0,
  u1,
  u2,
  v0,
  v1,
  v2,
  w0,
  w1,
  x0,
  x1,
  y0,
  y1;
output
  z2,
  z3,
  z4,
  a3,
  a4,
  a5,
  b3,
  b4,
  b5,
  c3,
  c4,
  c5,
  d3,
  d4,
  d5,
  e3,
  e4,
  e5,
  f3,
  f4,
  f5,
  g3,
  g4,
  g5,
  h3,
  h4,
  h5,
  i3,
  i4,
  i5,
  j3,
  j4,
  j5,
  k3,
  k4,
  k5,
  l3,
  l4,
  l5,
  m3,
  m4,
  m5,
  n3,
  n4,
  n5,
  o3,
  o4,
  o5,
  p3,
  p4,
  q3,
  q4,
  r3,
  r4,
  s3,
  s4,
  t3,
  t4,
  u3,
  u4,
  v3,
  v4,
  w2,
  w3,
  w4,
  x2,
  x3,
  x4,
  y2,
  y3,
  y4;
wire
  \[60] ,
  j11,
  j13,
  j14,
  \[61] ,
  \[62] ,
  \[63] ,
  r12,
  \[64] ,
  \[65] ,
  \[66] ,
  z10,
  z11,
  z13,
  \[67] ,
  \[68] ,
  \[69] ,
  \[0] ,
  \[1] ,
  c11,
  c12,
  c14,
  \[2] ,
  \[3] ,
  \[4] ,
  \[70] ,
  k11,
  k14,
  \[5] ,
  \[6] ,
  \[7] ,
  \[8] ,
  \[9] ,
  d10,
  d13,
  d14,
  l10,
  l11,
  l12,
  l14,
  t11,
  \[10] ,
  e10,
  e11,
  e14,
  \[11] ,
  \[12] ,
  \[13] ,
  m13,
  \[14] ,
  \[15] ,
  \[16] ,
  u10,
  u12,
  u13,
  \[17] ,
  \[18] ,
  \[19] ,
  \[20] ,
  f10,
  f11,
  f12,
  f14,
  \[21] ,
  \[22] ,
  \[23] ,
  n10,
  n11,
  \[24] ,
  \[25] ,
  \[26] ,
  v10,
  v13,
  \[27] ,
  \[28] ,
  \[29] ,
  \[30] ,
  g10,
  g13,
  g14,
  \[31] ,
  \[32] ,
  \[33] ,
  o12,
  \[34] ,
  \[35] ,
  \[36] ,
  w11,
  w13,
  \[37] ,
  \[38] ,
  \[39] ,
  \[40] ,
  h14,
  \[41] ,
  \[42] ,
  \[43] ,
  p13,
  \[44] ,
  \[45] ,
  \[46] ,
  x10,
  x12,
  x13,
  \[47] ,
  \[48] ,
  \[49] ,
  f9,
  a11,
  a13,
  a14,
  i9,
  \[50] ,
  j8,
  i11,
  i12,
  \[51] ,
  k8,
  k9,
  \[52] ,
  l9,
  \[53] ,
  m8,
  q11,
  \[54] ,
  \[55] ,
  o8,
  \[56] ,
  y10,
  y13,
  \[57] ,
  \[58] ,
  \[59] ,
  w8,
  b14,
  x8;
assign
  \[60]  = (~x13 & (~w13 & ~u13)) | ((~x13 & (~w13 & u2)) | ((~x13 & (~w13 & l2)) | ((~x13 & (~u13 & ~l2)) | ((~x13 & (~u13 & ~k2)) | ((~x13 & (u2 & ~l2)) | ((~x13 & (u2 & ~k2)) | (~x13 & (l2 & ~k2)))))))),
  z2 = \[3] ,
  z3 = \[29] ,
  z4 = \[55] ,
  j11 = ~e1 | ~q1,
  j13 = ~e1 | ~h2,
  j14 = (u0 & ~u2) | ((~u2 & ~b) | i0),
  \[61]  = (~y13 & (~w13 & ~u13)) | ((~y13 & (~w13 & u2)) | ((~y13 & (~w13 & m2)) | ((~y13 & (~u13 & ~m2)) | ((~y13 & (~u13 & ~l2)) | ((~y13 & (u2 & ~m2)) | ((~y13 & (u2 & ~l2)) | (~y13 & (m2 & ~l2)))))))),
  \[62]  = (~a14 & ~z13) | ((~a14 & d1) | ((~a14 & e1) | (~a14 & n2))),
  \[63]  = (~c14 & (~b14 & ~z13)) | ((~c14 & (~b14 & d1)) | ((~c14 & (~b14 & e1)) | ((~c14 & (~b14 & o2)) | ((~c14 & (~z13 & ~o2)) | ((~c14 & (~z13 & ~n2)) | ((~c14 & (d1 & ~o2)) | ((~c14 & (d1 & ~n2)) | ((~c14 & (e1 & ~o2)) | ((~c14 & (e1 & ~n2)) | (~c14 & (o2 & ~n2))))))))))),
  r12 = ~e1 | ~b2,
  \[64]  = (~d14 & (~b14 & ~z13)) | ((~d14 & (~b14 & d1)) | ((~d14 & (~b14 & e1)) | ((~d14 & (~b14 & p2)) | ((~d14 & (~z13 & ~p2)) | ((~d14 & (~z13 & ~o2)) | ((~d14 & (~z13 & ~n2)) | ((~d14 & (d1 & ~p2)) | ((~d14 & (d1 & ~o2)) | ((~d14 & (d1 & ~n2)) | ((~d14 & (e1 & ~p2)) | ((~d14 & (e1 & ~o2)) | ((~d14 & (e1 & ~n2)) | ((~d14 & (p2 & ~o2)) | (~d14 & (p2 & ~n2))))))))))))))),
  \[65]  = (~f14 & (~z13 & ~b14)) | ((~f14 & (~z13 & ~e14)) | ((~f14 & (~z13 & ~n2)) | ((~f14 & (~z13 & ~o2)) | ((~f14 & (d1 & ~b14)) | ((~f14 & (d1 & ~e14)) | ((~f14 & (d1 & ~n2)) | ((~f14 & (d1 & ~o2)) | ((~f14 & (e1 & ~b14)) | ((~f14 & (e1 & ~e14)) | ((~f14 & (e1 & ~n2)) | ((~f14 & (e1 & ~o2)) | ((~f14 & (q2 & ~b14)) | ((~f14 & (q2 & ~e14)) | ((~f14 & (q2 & ~n2)) | (~f14 & (q2 & ~o2)))))))))))))))),
  \[66]  = (~c1 & (~h14 & (~g14 & ~z13))) | ((~c1 & (~h14 & (~g14 & d1))) | ((~c1 & (~h14 & (~g14 & e1))) | ((~c1 & (~h14 & (~b14 & ~z13))) | ((~c1 & (~h14 & (~b14 & d1))) | ((~c1 & (~h14 & (~b14 & e1))) | ((~c1 & (~h14 & (~z13 & ~o2))) | ((~c1 & (~h14 & (~z13 & ~n2))) | ((~c1 & (~h14 & (d1 & ~o2))) | ((~c1 & (~h14 & (d1 & ~n2))) | ((~c1 & (~h14 & (e1 & ~o2))) | ((~c1 & (~h14 & (e1 & ~n2))) | ((~c1 & (~g14 & r2)) | ((~c1 & (~b14 & r2)) | ((~c1 & (r2 & ~o2)) | (~c1 & (r2 & ~n2)))))))))))))))),
  z10 = (m1 & (v2 & (g0 & ~h0))) | ((m1 & (v2 & (g0 & h))) | (m1 & (v2 & (g0 & g)))),
  z11 = ~e1 | ~v1,
  z13 = k2 | (~l2 | ~m2),
  \[67]  = (n1 & (e1 & (~m0 & ~i0))) | ((n1 & (b1 & ~i0)) | ((b1 & (~e1 & ~i0)) | (b1 & (m0 & ~i0)))),
  \[68]  = (~t2 & (s2 & (l1 & ~c1))) | ((t2 & (~s2 & ~c1)) | (t2 & (~l1 & ~c1))),
  \[69]  = (~j14 & ~u13) | ((~j14 & k2) | ((~j14 & ~l2) | (~j14 & ~m2))),
  \[0]  = ~f1,
  \[1]  = ~g1,
  c11 = (m1 & (h & (g0 & v2))) | ((m1 & (g & (g0 & v2))) | ((m1 & (g0 & (v2 & ~h0))) | (e1 & ~m0))),
  c12 = ~e1 | ~w1,
  c14 = (~o2 & ~n2) | c1,
  \[2]  = ~h1,
  \[3]  = ~i1,
  \[4]  = ~j1,
  \[70]  = (~v10 & (v2 & ~f0)) | (~k14 & ~v10),
  k11 = (m1 & (v2 & (g0 & ~h0))) | ((m1 & (v2 & (g0 & i))) | ((m1 & (v2 & (g0 & h))) | (m1 & (v2 & (g0 & g))))),
  k14 = ~l14 | (~n2 | ~e1),
  \[5]  = ~k1,
  \[6]  = (~k8 & (~j8 & (e1 & ~i0))) | (~m8 & (s2 & ~i0)),
  \[7]  = (~w8 & (g0 & (~c1 & v2))) | ~x8,
  \[8]  = (~f9 & (n2 & (e1 & ~c1))) | (l0 & ~c1),
  \[9]  = (~w8 & (g0 & v2)) | ~i9,
  d10 = o2 | (p2 | ~r2),
  d13 = ~e1 | ~f2,
  d14 = (~p2 & ~o2) | ((~p2 & ~n2) | c1),
  l10 = o2 & (~p2 & (~q2 & ~r2)),
  l11 = (~e11 & (g0 & (m1 & v2))) | (~m0 & e1),
  l12 = ~e1 | ~z1,
  l14 = (r2 & (~o2 & (~p2 & q2))) | (r2 & (~o2 & (~p2 & i))),
  t11 = ~e1 | ~t1,
  \[10]  = ~k9 & (~i0 & ~c1),
  e10 = ~i & ~q2,
  e11 = ~g & (~h & (~i & h0)),
  e14 = p2 & q2,
  \[11]  = ~i0 & (o0 & ~c1),
  \[12]  = ~i0 & (p0 & ~c1),
  \[13]  = ~i0 & (q0 & ~c1),
  m13 = ~e1 | ~i2,
  \[14]  = ~i0 & (r0 & ~c1),
  \[15]  = ~i0 & (s0 & ~c1),
  \[16]  = ~i0 & (t0 & ~c1),
  u10 = ~x10 | (g | (h | k2)),
  u12 = ~e1 | ~c2,
  u13 = ~b | u0,
  \[17]  = b & ~i0,
  \[18]  = a & ~i0,
  \[19]  = ~i0 & v0,
  \[20]  = ~i0 & w0,
  f10 = (~v2 & ~i0) | (~i0 & ~f0),
  f11 = (p1 & (e1 & (~m0 & ~i0))) | ((p1 & (~o1 & ~i0)) | ((~o1 & (~e1 & ~i0)) | (~o1 & (m0 & ~i0)))),
  f12 = ~e1 | ~x1,
  f14 = (~q2 & ~p2) | ((~q2 & ~o2) | ((~q2 & ~n2) | c1)),
  \[21]  = ~i0 & x0,
  \[22]  = ~i0 & y0,
  \[23]  = ~i0 & z0,
  n10 = ~l9 | (~e1 | (n2 | ~o2)),
  n11 = ~e1 | ~r1,
  \[24]  = ~i0 & a1,
  \[25]  = (~e10 & (~d10 & (e1 & n2))) | ((~w8 & (g0 & v2)) | ~f10),
  \[26]  = ~g10 & v2,
  v10 = (g0 & v2) | i0,
  v13 = (k2 & (b & ~u0)) | ((u2 & k2) | c1),
  \[27]  = (m2 & (l2 & (~k2 & ~c1))) | ((d1 & ~c1) | (e1 & ~c1)),
  \[28]  = (~c1 & (~n10 & ~l10)) | ((~c1 & (~n10 & o0)) | ((~c1 & (~n10 & ~e1)) | ((~c1 & (~n10 & n2)) | ((~c1 & (f1 & ~l10)) | ((~c1 & (f1 & o0)) | ((~c1 & (f1 & ~e1)) | (~c1 & (f1 & n2)))))))),
  \[29]  = (~c1 & (~n10 & ~l10)) | ((~c1 & (~n10 & p0)) | ((~c1 & (~n10 & ~e1)) | ((~c1 & (~n10 & n2)) | ((~c1 & (g1 & ~l10)) | ((~c1 & (g1 & p0)) | ((~c1 & (g1 & ~e1)) | (~c1 & (g1 & n2)))))))),
  \[30]  = (~c1 & (~n10 & ~l10)) | ((~c1 & (~n10 & q0)) | ((~c1 & (~n10 & ~e1)) | ((~c1 & (~n10 & n2)) | ((~c1 & (h1 & ~l10)) | ((~c1 & (h1 & q0)) | ((~c1 & (h1 & ~e1)) | (~c1 & (h1 & n2)))))))),
  g10 = (h0 & (~i & (~h & ~g))) | (m1 | (g0 | ~i0)),
  g13 = ~e1 | ~g2,
  g14 = p2 & (q2 & r2),
  \[31]  = (~c1 & (~n10 & ~l10)) | ((~c1 & (~n10 & r0)) | ((~c1 & (~n10 & ~e1)) | ((~c1 & (~n10 & n2)) | ((~c1 & (i1 & ~l10)) | ((~c1 & (i1 & r0)) | ((~c1 & (i1 & ~e1)) | (~c1 & (i1 & n2)))))))),
  \[32]  = (~c1 & (~n10 & ~l10)) | ((~c1 & (~n10 & s0)) | ((~c1 & (~n10 & ~e1)) | ((~c1 & (~n10 & n2)) | ((~c1 & (j1 & ~l10)) | ((~c1 & (j1 & s0)) | ((~c1 & (j1 & ~e1)) | (~c1 & (j1 & n2)))))))),
  \[33]  = (~c1 & (~n10 & ~l10)) | ((~c1 & (~n10 & t0)) | ((~c1 & (~n10 & ~e1)) | ((~c1 & (~n10 & n2)) | ((~c1 & (k1 & ~l10)) | ((~c1 & (k1 & t0)) | ((~c1 & (k1 & ~e1)) | (~c1 & (k1 & n2)))))))),
  o12 = ~e1 | ~a2,
  \[34]  = (~f9 & (n2 & (e1 & ~c1))) | (l1 & ~c1),
  \[35]  = (~v10 & ~u10) | (~v10 & m1),
  \[36]  = (~a11 & (i & (g0 & ~i0))) | ((~z10 & (~y10 & (~m0 & ~i0))) | (~c11 & (n1 & ~i0))),
  w11 = ~e1 | ~u1,
  w13 = (b & ~u0) | u2,
  \[37]  = (~e11 & (g0 & (m1 & v2))) | ~f11,
  \[38]  = (~k11 & (~j11 & (~m0 & ~i0))) | ((~i11 & (k & (~e11 & g0))) | (~l11 & (p1 & ~i0))),
  \[39]  = (~n11 & (~k11 & (~m0 & ~i0))) | ((l & (~i11 & (~e11 & g0))) | (q1 & (~l11 & ~i0))),
  \[40]  = (~q11 & (~k11 & (~m0 & ~i0))) | ((m & (~i11 & (~e11 & g0))) | (r1 & (~l11 & ~i0))),
  h14 = ~n2 | (~o2 | (~p2 | ~q2)),
  \[41]  = (~t11 & (~k11 & (~m0 & ~i0))) | ((n & (~i11 & (~e11 & g0))) | (s1 & (~l11 & ~i0))),
  \[42]  = (~w11 & (~k11 & (~m0 & ~i0))) | ((o & (~i11 & (~e11 & g0))) | (t1 & (~l11 & ~i0))),
  \[43]  = (~z11 & (~k11 & (~m0 & ~i0))) | ((p & (~i11 & (~e11 & g0))) | (u1 & (~l11 & ~i0))),
  p13 = ~e1 | ~j2,
  \[44]  = (~c12 & (~k11 & (~m0 & ~i0))) | ((q & (~i11 & (~e11 & g0))) | (v1 & (~l11 & ~i0))),
  \[45]  = (~f12 & (~k11 & (~m0 & ~i0))) | ((r & (~i11 & (~e11 & g0))) | (w1 & (~l11 & ~i0))),
  \[46]  = (~i12 & (~k11 & (~m0 & ~i0))) | ((s & (~i11 & (~e11 & g0))) | (x1 & (~l11 & ~i0))),
  x10 = l2 & m2,
  x12 = ~e1 | ~d2,
  x13 = (m2 & ~k2) | ((~l2 & ~k2) | c1),
  \[47]  = (~l12 & (~k11 & (~m0 & ~i0))) | ((t & (~i11 & (~e11 & g0))) | (y1 & (~l11 & ~i0))),
  a3 = \[4] ,
  a4 = \[30] ,
  a5 = \[56] ,
  \[48]  = (~o12 & (~k11 & (~m0 & ~i0))) | ((u & (~i11 & (~e11 & g0))) | (z1 & (~l11 & ~i0))),
  b3 = \[5] ,
  b4 = \[31] ,
  b5 = \[57] ,
  \[49]  = (~r12 & (~k11 & (~m0 & ~i0))) | ((v & (~i11 & (~e11 & g0))) | (a2 & (~l11 & ~i0))),
  c3 = \[6] ,
  c4 = \[32] ,
  c5 = \[58] ,
  d3 = \[7] ,
  d4 = \[33] ,
  d5 = \[59] ,
  e3 = \[8] ,
  e4 = \[34] ,
  e5 = \[60] ,
  f3 = \[9] ,
  f4 = \[35] ,
  f5 = \[61] ,
  f9 = o2 | (p2 | (q2 | r2)),
  g3 = \[10] ,
  g4 = \[36] ,
  g5 = \[62] ,
  a11 = ~m1 | ~v2,
  a13 = ~e1 | ~e2,
  a14 = (m2 & (l2 & (n2 & ~k2))) | ((d1 & n2) | ((n2 & e1) | c1)),
  h3 = \[11] ,
  h4 = \[37] ,
  h5 = \[63] ,
  i3 = \[12] ,
  i4 = \[38] ,
  i5 = \[64] ,
  i9 = (g0 & (v2 & ~i0)) | (~m0 & ~i0),
  \[50]  = (~u12 & (~k11 & (~m0 & ~i0))) | ((w & (~i11 & (~e11 & g0))) | (b2 & (~l11 & ~i0))),
  j3 = \[13] ,
  j4 = \[39] ,
  j5 = \[65] ,
  j8 = ~n2 | (o2 | (p2 | ~r2)),
  i11 = i0 | (~m1 | ~v2),
  i12 = ~e1 | ~y1,
  \[51]  = (~x12 & (~k11 & (~m0 & ~i0))) | ((\xx  & (~i11 & (~e11 & g0))) | (c2 & (~l11 & ~i0))),
  k3 = \[14] ,
  k4 = \[40] ,
  k5 = \[66] ,
  k8 = (~t2 & h0) | ((t2 & ~h0) | (~q2 & ~i)),
  k9 = (~n0 & ~l9) | ((~n0 & ~e1) | ((~n0 & ~n2) | (~n0 & o2))),
  \[52]  = (~a13 & (~k11 & (~m0 & ~i0))) | ((y & (~i11 & (~e11 & g0))) | (d2 & (~l11 & ~i0))),
  l3 = \[15] ,
  l4 = \[41] ,
  l5 = \[67] ,
  l9 = ~p2 & (~q2 & ~r2),
  \[53]  = (~d13 & (~k11 & (~m0 & ~i0))) | ((z & (~i11 & (~e11 & g0))) | (e2 & (~l11 & ~i0))),
  m3 = \[16] ,
  m4 = \[42] ,
  m5 = \[68] ,
  m8 = ~o8 & (r2 & ~p2),
  q11 = ~e1 | ~s1,
  \[54]  = (~g13 & (~k11 & (~m0 & ~i0))) | ((a0 & (~i11 & (~e11 & g0))) | (f2 & (~l11 & ~i0))),
  n3 = \[17] ,
  n4 = \[43] ,
  n5 = \[69] ,
  \[55]  = (~j13 & (~k11 & (~m0 & ~i0))) | ((b0 & (~i11 & (~e11 & g0))) | (g2 & (~l11 & ~i0))),
  o3 = \[18] ,
  o4 = \[44] ,
  o5 = \[70] ,
  o8 = (~q2 & ~i) | (o2 | (~e1 | ~n2)),
  \[56]  = (~m13 & (~k11 & (~m0 & ~i0))) | ((c0 & (~i11 & (~e11 & g0))) | (h2 & (~l11 & ~i0))),
  p3 = \[19] ,
  p4 = \[45] ,
  y10 = ~e1 | o1,
  y13 = (~m2 & ~l2) | ((~m2 & ~k2) | ((l2 & ~k2) | c1)),
  \[57]  = (~p13 & (~k11 & (~m0 & ~i0))) | ((d0 & (~i11 & (~e11 & g0))) | (i2 & (~l11 & ~i0))),
  q3 = \[20] ,
  q4 = \[46] ,
  \[58]  = (~e11 & (~i11 & (e0 & g0))) | (~l11 & (~i0 & j2)),
  r3 = \[21] ,
  r4 = \[47] ,
  \[59]  = (~v13 & ~u13) | ((~v13 & k2) | (~v13 & u2)),
  s3 = \[22] ,
  s4 = \[48] ,
  t3 = \[23] ,
  t4 = \[49] ,
  u3 = \[24] ,
  u4 = \[50] ,
  v3 = \[25] ,
  v4 = \[51] ,
  w2 = \[0] ,
  w3 = \[26] ,
  w4 = \[52] ,
  w8 = (m1 & ~h0) | ((m1 & i) | ((m1 & h) | (m1 & g))),
  b14 = (m2 & (l2 & ~k2)) | (d1 | e1),
  x2 = \[1] ,
  x3 = \[27] ,
  x4 = \[53] ,
  x8 = (~v2 & ~k0) | ((~k0 & ~f0) | c1),
  y2 = \[2] ,
  y3 = \[28] ,
  y4 = \[54] ;
endmodule

